module handshake_synchronizer (dst_clk,
    dst_ready,
    dst_rst_n,
    dst_valid,
    src_clk,
    src_ready,
    src_rst_n,
    src_valid,
    dst_data,
    src_data);
 input dst_clk;
 input dst_ready;
 input dst_rst_n;
 output dst_valid;
 input src_clk;
 output src_ready;
 input src_rst_n;
 input src_valid;
 output [31:0] dst_data;
 input [31:0] src_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire \ack_sync[0] ;
 wire \ack_sync[1] ;
 wire \data_reg[0] ;
 wire \data_reg[10] ;
 wire \data_reg[11] ;
 wire \data_reg[12] ;
 wire \data_reg[13] ;
 wire \data_reg[14] ;
 wire \data_reg[15] ;
 wire \data_reg[16] ;
 wire \data_reg[17] ;
 wire \data_reg[18] ;
 wire \data_reg[19] ;
 wire \data_reg[1] ;
 wire \data_reg[20] ;
 wire \data_reg[21] ;
 wire \data_reg[22] ;
 wire \data_reg[23] ;
 wire \data_reg[24] ;
 wire \data_reg[25] ;
 wire \data_reg[26] ;
 wire \data_reg[27] ;
 wire \data_reg[28] ;
 wire \data_reg[29] ;
 wire \data_reg[2] ;
 wire \data_reg[30] ;
 wire \data_reg[31] ;
 wire \data_reg[3] ;
 wire \data_reg[4] ;
 wire \data_reg[5] ;
 wire \data_reg[6] ;
 wire \data_reg[7] ;
 wire \data_reg[8] ;
 wire \data_reg[9] ;
 wire dst_ack;
 wire dst_req;
 wire \req_sync[0] ;
 wire src_req;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire clknet_0_src_clk;
 wire clknet_2_0__leaf_src_clk;
 wire clknet_2_1__leaf_src_clk;
 wire clknet_2_2__leaf_src_clk;
 wire clknet_2_3__leaf_src_clk;
 wire net72;
 wire net73;
 wire net74;

 XNOR2_X2 _154_ (.A(src_req),
    .B(\ack_sync[1] ),
    .ZN(net71));
 NAND2_X4 _155_ (.A1(net37),
    .A2(net71),
    .ZN(_068_));
 BUF_X4 _156_ (.A(_068_),
    .Z(_069_));
 MUX2_X1 _157_ (.A(net4),
    .B(\data_reg[0] ),
    .S(_069_),
    .Z(_001_));
 MUX2_X1 _158_ (.A(net5),
    .B(\data_reg[10] ),
    .S(_069_),
    .Z(_002_));
 MUX2_X1 _159_ (.A(net6),
    .B(\data_reg[11] ),
    .S(_069_),
    .Z(_003_));
 MUX2_X1 _160_ (.A(net7),
    .B(\data_reg[12] ),
    .S(_069_),
    .Z(_004_));
 MUX2_X1 _161_ (.A(net8),
    .B(\data_reg[13] ),
    .S(_069_),
    .Z(_005_));
 MUX2_X1 _162_ (.A(net9),
    .B(\data_reg[14] ),
    .S(_069_),
    .Z(_006_));
 MUX2_X1 _163_ (.A(net10),
    .B(\data_reg[15] ),
    .S(_069_),
    .Z(_007_));
 MUX2_X1 _164_ (.A(net11),
    .B(\data_reg[16] ),
    .S(_069_),
    .Z(_008_));
 MUX2_X1 _165_ (.A(net12),
    .B(\data_reg[17] ),
    .S(_069_),
    .Z(_009_));
 MUX2_X1 _166_ (.A(net13),
    .B(\data_reg[18] ),
    .S(_069_),
    .Z(_010_));
 BUF_X8 _167_ (.A(_068_),
    .Z(_070_));
 MUX2_X1 _168_ (.A(net14),
    .B(\data_reg[19] ),
    .S(_070_),
    .Z(_011_));
 MUX2_X1 _169_ (.A(net15),
    .B(\data_reg[1] ),
    .S(_070_),
    .Z(_012_));
 MUX2_X1 _170_ (.A(net16),
    .B(\data_reg[20] ),
    .S(_070_),
    .Z(_013_));
 MUX2_X1 _171_ (.A(net17),
    .B(\data_reg[21] ),
    .S(_070_),
    .Z(_014_));
 MUX2_X1 _172_ (.A(net18),
    .B(\data_reg[22] ),
    .S(_070_),
    .Z(_015_));
 MUX2_X1 _173_ (.A(net19),
    .B(\data_reg[23] ),
    .S(_070_),
    .Z(_016_));
 MUX2_X1 _174_ (.A(net20),
    .B(\data_reg[24] ),
    .S(_070_),
    .Z(_017_));
 MUX2_X1 _175_ (.A(net21),
    .B(\data_reg[25] ),
    .S(_070_),
    .Z(_018_));
 MUX2_X1 _176_ (.A(net22),
    .B(\data_reg[26] ),
    .S(_070_),
    .Z(_019_));
 MUX2_X1 _177_ (.A(net23),
    .B(\data_reg[27] ),
    .S(_070_),
    .Z(_020_));
 BUF_X8 _178_ (.A(_068_),
    .Z(_071_));
 MUX2_X1 _179_ (.A(net24),
    .B(\data_reg[28] ),
    .S(_071_),
    .Z(_021_));
 MUX2_X1 _180_ (.A(net25),
    .B(\data_reg[29] ),
    .S(_071_),
    .Z(_022_));
 MUX2_X1 _181_ (.A(net26),
    .B(\data_reg[2] ),
    .S(_071_),
    .Z(_023_));
 MUX2_X1 _182_ (.A(net27),
    .B(\data_reg[30] ),
    .S(_071_),
    .Z(_024_));
 MUX2_X1 _183_ (.A(net28),
    .B(\data_reg[31] ),
    .S(_071_),
    .Z(_025_));
 MUX2_X1 _184_ (.A(net29),
    .B(\data_reg[3] ),
    .S(_071_),
    .Z(_026_));
 MUX2_X1 _185_ (.A(net30),
    .B(\data_reg[4] ),
    .S(_071_),
    .Z(_027_));
 MUX2_X1 _186_ (.A(net31),
    .B(\data_reg[5] ),
    .S(_071_),
    .Z(_028_));
 MUX2_X1 _187_ (.A(net32),
    .B(\data_reg[6] ),
    .S(_071_),
    .Z(_029_));
 MUX2_X1 _188_ (.A(net33),
    .B(\data_reg[7] ),
    .S(_071_),
    .Z(_030_));
 MUX2_X1 _189_ (.A(net34),
    .B(\data_reg[8] ),
    .S(_068_),
    .Z(_031_));
 MUX2_X1 _190_ (.A(net35),
    .B(\data_reg[9] ),
    .S(_068_),
    .Z(_032_));
 NAND2_X1 _191_ (.A1(net2),
    .A2(net70),
    .ZN(_072_));
 MUX2_X1 _192_ (.A(dst_req),
    .B(dst_ack),
    .S(_072_),
    .Z(_033_));
 XNOR2_X2 _193_ (.A(dst_ack),
    .B(dst_req),
    .ZN(_073_));
 NOR2_X4 _194_ (.A1(net70),
    .A2(_073_),
    .ZN(_074_));
 BUF_X8 _195_ (.A(_074_),
    .Z(_075_));
 MUX2_X1 _196_ (.A(net38),
    .B(\data_reg[0] ),
    .S(_075_),
    .Z(_034_));
 MUX2_X1 _197_ (.A(net39),
    .B(\data_reg[10] ),
    .S(_075_),
    .Z(_035_));
 MUX2_X1 _198_ (.A(net40),
    .B(\data_reg[11] ),
    .S(_075_),
    .Z(_036_));
 MUX2_X1 _199_ (.A(net41),
    .B(\data_reg[12] ),
    .S(_075_),
    .Z(_037_));
 MUX2_X1 _200_ (.A(net42),
    .B(\data_reg[13] ),
    .S(_075_),
    .Z(_038_));
 MUX2_X1 _201_ (.A(net43),
    .B(\data_reg[14] ),
    .S(_075_),
    .Z(_039_));
 MUX2_X1 _202_ (.A(net44),
    .B(\data_reg[15] ),
    .S(_075_),
    .Z(_040_));
 MUX2_X1 _203_ (.A(net45),
    .B(\data_reg[16] ),
    .S(_075_),
    .Z(_041_));
 MUX2_X1 _204_ (.A(net46),
    .B(\data_reg[17] ),
    .S(_075_),
    .Z(_042_));
 MUX2_X1 _205_ (.A(net47),
    .B(\data_reg[18] ),
    .S(_075_),
    .Z(_043_));
 BUF_X8 _206_ (.A(_074_),
    .Z(_076_));
 MUX2_X1 _207_ (.A(net48),
    .B(\data_reg[19] ),
    .S(_076_),
    .Z(_044_));
 MUX2_X1 _208_ (.A(net49),
    .B(\data_reg[1] ),
    .S(_076_),
    .Z(_045_));
 MUX2_X1 _209_ (.A(net50),
    .B(\data_reg[20] ),
    .S(_076_),
    .Z(_046_));
 MUX2_X1 _210_ (.A(net51),
    .B(\data_reg[21] ),
    .S(_076_),
    .Z(_047_));
 MUX2_X1 _211_ (.A(net52),
    .B(\data_reg[22] ),
    .S(_076_),
    .Z(_048_));
 MUX2_X1 _212_ (.A(net53),
    .B(\data_reg[23] ),
    .S(_076_),
    .Z(_049_));
 MUX2_X1 _213_ (.A(net54),
    .B(\data_reg[24] ),
    .S(_076_),
    .Z(_050_));
 MUX2_X1 _214_ (.A(net55),
    .B(\data_reg[25] ),
    .S(_076_),
    .Z(_051_));
 MUX2_X1 _215_ (.A(net56),
    .B(\data_reg[26] ),
    .S(_076_),
    .Z(_052_));
 MUX2_X1 _216_ (.A(net57),
    .B(\data_reg[27] ),
    .S(_076_),
    .Z(_053_));
 BUF_X8 _217_ (.A(_074_),
    .Z(_077_));
 MUX2_X1 _218_ (.A(net58),
    .B(\data_reg[28] ),
    .S(_077_),
    .Z(_054_));
 MUX2_X1 _219_ (.A(net59),
    .B(\data_reg[29] ),
    .S(_077_),
    .Z(_055_));
 MUX2_X1 _220_ (.A(net60),
    .B(\data_reg[2] ),
    .S(_077_),
    .Z(_056_));
 MUX2_X1 _221_ (.A(net61),
    .B(\data_reg[30] ),
    .S(_077_),
    .Z(_057_));
 MUX2_X1 _222_ (.A(net62),
    .B(\data_reg[31] ),
    .S(_077_),
    .Z(_058_));
 MUX2_X1 _223_ (.A(net63),
    .B(\data_reg[3] ),
    .S(_077_),
    .Z(_059_));
 MUX2_X1 _224_ (.A(net64),
    .B(\data_reg[4] ),
    .S(_077_),
    .Z(_060_));
 MUX2_X1 _225_ (.A(net65),
    .B(\data_reg[5] ),
    .S(_077_),
    .Z(_061_));
 MUX2_X1 _226_ (.A(net66),
    .B(\data_reg[6] ),
    .S(_077_),
    .Z(_062_));
 MUX2_X1 _227_ (.A(net67),
    .B(\data_reg[7] ),
    .S(_077_),
    .Z(_063_));
 MUX2_X1 _228_ (.A(net68),
    .B(\data_reg[8] ),
    .S(_074_),
    .Z(_064_));
 MUX2_X1 _229_ (.A(net69),
    .B(\data_reg[9] ),
    .S(_074_),
    .Z(_065_));
 INV_X1 _230_ (.A(net70),
    .ZN(_078_));
 NAND2_X1 _231_ (.A1(_078_),
    .A2(_073_),
    .ZN(_079_));
 AND2_X1 _232_ (.A1(_072_),
    .A2(_079_),
    .ZN(_066_));
 INV_X1 _233_ (.A(\ack_sync[1] ),
    .ZN(_080_));
 AOI21_X1 _234_ (.A(src_req),
    .B1(_080_),
    .B2(net37),
    .ZN(_081_));
 NAND2_X1 _235_ (.A1(net37),
    .A2(\ack_sync[1] ),
    .ZN(_082_));
 AOI21_X1 _236_ (.A(_000_),
    .B1(_082_),
    .B2(src_req),
    .ZN(_083_));
 NOR2_X1 _237_ (.A1(_081_),
    .A2(_083_),
    .ZN(_067_));
 DFFR_X1 \ack_sync[0]$_DFF_PN0_  (.D(dst_ack),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\ack_sync[0] ),
    .QN(_151_));
 DFFR_X1 \ack_sync[1]$_DFF_PN0_  (.D(\ack_sync[0] ),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\ack_sync[1] ),
    .QN(_150_));
 DFFR_X1 \data_reg[0]$_DFFE_PN0P_  (.D(_001_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[0] ),
    .QN(_149_));
 DFFR_X1 \data_reg[10]$_DFFE_PN0P_  (.D(_002_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[10] ),
    .QN(_148_));
 DFFR_X1 \data_reg[11]$_DFFE_PN0P_  (.D(_003_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[11] ),
    .QN(_147_));
 DFFR_X1 \data_reg[12]$_DFFE_PN0P_  (.D(_004_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[12] ),
    .QN(_146_));
 DFFR_X1 \data_reg[13]$_DFFE_PN0P_  (.D(_005_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[13] ),
    .QN(_145_));
 DFFR_X1 \data_reg[14]$_DFFE_PN0P_  (.D(_006_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[14] ),
    .QN(_144_));
 DFFR_X1 \data_reg[15]$_DFFE_PN0P_  (.D(_007_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[15] ),
    .QN(_143_));
 DFFR_X1 \data_reg[16]$_DFFE_PN0P_  (.D(_008_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[16] ),
    .QN(_142_));
 DFFR_X1 \data_reg[17]$_DFFE_PN0P_  (.D(_009_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[17] ),
    .QN(_141_));
 DFFR_X1 \data_reg[18]$_DFFE_PN0P_  (.D(_010_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[18] ),
    .QN(_140_));
 DFFR_X1 \data_reg[19]$_DFFE_PN0P_  (.D(_011_),
    .RN(net36),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[19] ),
    .QN(_139_));
 DFFR_X1 \data_reg[1]$_DFFE_PN0P_  (.D(_012_),
    .RN(net36),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[1] ),
    .QN(_138_));
 DFFR_X1 \data_reg[20]$_DFFE_PN0P_  (.D(_013_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[20] ),
    .QN(_137_));
 DFFR_X1 \data_reg[21]$_DFFE_PN0P_  (.D(_014_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[21] ),
    .QN(_136_));
 DFFR_X1 \data_reg[22]$_DFFE_PN0P_  (.D(_015_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[22] ),
    .QN(_135_));
 DFFR_X1 \data_reg[23]$_DFFE_PN0P_  (.D(_016_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[23] ),
    .QN(_134_));
 DFFR_X1 \data_reg[24]$_DFFE_PN0P_  (.D(_017_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[24] ),
    .QN(_133_));
 DFFR_X1 \data_reg[25]$_DFFE_PN0P_  (.D(_018_),
    .RN(net73),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[25] ),
    .QN(_132_));
 DFFR_X1 \data_reg[26]$_DFFE_PN0P_  (.D(_019_),
    .RN(net73),
    .CK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[26] ),
    .QN(_131_));
 DFFR_X1 \data_reg[27]$_DFFE_PN0P_  (.D(_020_),
    .RN(net36),
    .CK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[27] ),
    .QN(_130_));
 DFFR_X1 \data_reg[28]$_DFFE_PN0P_  (.D(_021_),
    .RN(net36),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[28] ),
    .QN(_129_));
 DFFR_X1 \data_reg[29]$_DFFE_PN0P_  (.D(_022_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[29] ),
    .QN(_128_));
 DFFR_X1 \data_reg[2]$_DFFE_PN0P_  (.D(_023_),
    .RN(net36),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[2] ),
    .QN(_127_));
 DFFR_X1 \data_reg[30]$_DFFE_PN0P_  (.D(_024_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[30] ),
    .QN(_126_));
 DFFR_X1 \data_reg[31]$_DFFE_PN0P_  (.D(_025_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[31] ),
    .QN(_125_));
 DFFR_X1 \data_reg[3]$_DFFE_PN0P_  (.D(_026_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[3] ),
    .QN(_124_));
 DFFR_X1 \data_reg[4]$_DFFE_PN0P_  (.D(_027_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[4] ),
    .QN(_123_));
 DFFR_X1 \data_reg[5]$_DFFE_PN0P_  (.D(_028_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[5] ),
    .QN(_122_));
 DFFR_X1 \data_reg[6]$_DFFE_PN0P_  (.D(_029_),
    .RN(net36),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[6] ),
    .QN(_121_));
 DFFR_X1 \data_reg[7]$_DFFE_PN0P_  (.D(_030_),
    .RN(net73),
    .CK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[7] ),
    .QN(_120_));
 DFFR_X1 \data_reg[8]$_DFFE_PN0P_  (.D(_031_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[8] ),
    .QN(_119_));
 DFFR_X1 \data_reg[9]$_DFFE_PN0P_  (.D(_032_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[9] ),
    .QN(_118_));
 DFFR_X1 \dst_ack$_DFFE_PN0P_  (.D(_033_),
    .RN(net3),
    .CK(net1),
    .Q(dst_ack),
    .QN(_117_));
 DFFR_X1 \dst_data_reg[0]$_DFFE_PN0P_  (.D(_034_),
    .RN(net3),
    .CK(net1),
    .Q(net38),
    .QN(_116_));
 DFFR_X1 \dst_data_reg[10]$_DFFE_PN0P_  (.D(_035_),
    .RN(net3),
    .CK(net1),
    .Q(net39),
    .QN(_115_));
 DFFR_X1 \dst_data_reg[11]$_DFFE_PN0P_  (.D(_036_),
    .RN(net3),
    .CK(net1),
    .Q(net40),
    .QN(_114_));
 DFFR_X1 \dst_data_reg[12]$_DFFE_PN0P_  (.D(_037_),
    .RN(net3),
    .CK(net1),
    .Q(net41),
    .QN(_113_));
 DFFR_X1 \dst_data_reg[13]$_DFFE_PN0P_  (.D(_038_),
    .RN(net3),
    .CK(net1),
    .Q(net42),
    .QN(_112_));
 DFFR_X1 \dst_data_reg[14]$_DFFE_PN0P_  (.D(_039_),
    .RN(net3),
    .CK(net1),
    .Q(net43),
    .QN(_111_));
 DFFR_X1 \dst_data_reg[15]$_DFFE_PN0P_  (.D(_040_),
    .RN(net3),
    .CK(net1),
    .Q(net44),
    .QN(_110_));
 DFFR_X1 \dst_data_reg[16]$_DFFE_PN0P_  (.D(_041_),
    .RN(net3),
    .CK(net1),
    .Q(net45),
    .QN(_109_));
 DFFR_X1 \dst_data_reg[17]$_DFFE_PN0P_  (.D(_042_),
    .RN(net3),
    .CK(net1),
    .Q(net46),
    .QN(_108_));
 DFFR_X1 \dst_data_reg[18]$_DFFE_PN0P_  (.D(_043_),
    .RN(net3),
    .CK(net1),
    .Q(net47),
    .QN(_107_));
 DFFR_X1 \dst_data_reg[19]$_DFFE_PN0P_  (.D(_044_),
    .RN(net3),
    .CK(net1),
    .Q(net48),
    .QN(_106_));
 DFFR_X1 \dst_data_reg[1]$_DFFE_PN0P_  (.D(_045_),
    .RN(net3),
    .CK(net1),
    .Q(net49),
    .QN(_105_));
 DFFR_X1 \dst_data_reg[20]$_DFFE_PN0P_  (.D(_046_),
    .RN(net3),
    .CK(net1),
    .Q(net50),
    .QN(_104_));
 DFFR_X1 \dst_data_reg[21]$_DFFE_PN0P_  (.D(_047_),
    .RN(net3),
    .CK(net1),
    .Q(net51),
    .QN(_103_));
 DFFR_X1 \dst_data_reg[22]$_DFFE_PN0P_  (.D(_048_),
    .RN(net3),
    .CK(net1),
    .Q(net52),
    .QN(_102_));
 DFFR_X1 \dst_data_reg[23]$_DFFE_PN0P_  (.D(_049_),
    .RN(net3),
    .CK(net1),
    .Q(net53),
    .QN(_101_));
 DFFR_X1 \dst_data_reg[24]$_DFFE_PN0P_  (.D(_050_),
    .RN(net3),
    .CK(net1),
    .Q(net54),
    .QN(_100_));
 DFFR_X1 \dst_data_reg[25]$_DFFE_PN0P_  (.D(_051_),
    .RN(net3),
    .CK(net1),
    .Q(net55),
    .QN(_099_));
 DFFR_X1 \dst_data_reg[26]$_DFFE_PN0P_  (.D(_052_),
    .RN(net3),
    .CK(net1),
    .Q(net56),
    .QN(_098_));
 DFFR_X1 \dst_data_reg[27]$_DFFE_PN0P_  (.D(_053_),
    .RN(net3),
    .CK(net1),
    .Q(net57),
    .QN(_097_));
 DFFR_X1 \dst_data_reg[28]$_DFFE_PN0P_  (.D(_054_),
    .RN(net3),
    .CK(net1),
    .Q(net58),
    .QN(_096_));
 DFFR_X1 \dst_data_reg[29]$_DFFE_PN0P_  (.D(_055_),
    .RN(net3),
    .CK(net1),
    .Q(net59),
    .QN(_095_));
 DFFR_X1 \dst_data_reg[2]$_DFFE_PN0P_  (.D(_056_),
    .RN(net3),
    .CK(net1),
    .Q(net60),
    .QN(_094_));
 DFFR_X1 \dst_data_reg[30]$_DFFE_PN0P_  (.D(_057_),
    .RN(net3),
    .CK(net1),
    .Q(net61),
    .QN(_093_));
 DFFR_X1 \dst_data_reg[31]$_DFFE_PN0P_  (.D(_058_),
    .RN(net3),
    .CK(net1),
    .Q(net62),
    .QN(_092_));
 DFFR_X1 \dst_data_reg[3]$_DFFE_PN0P_  (.D(_059_),
    .RN(net3),
    .CK(net1),
    .Q(net63),
    .QN(_091_));
 DFFR_X1 \dst_data_reg[4]$_DFFE_PN0P_  (.D(_060_),
    .RN(net3),
    .CK(net1),
    .Q(net64),
    .QN(_090_));
 DFFR_X1 \dst_data_reg[5]$_DFFE_PN0P_  (.D(_061_),
    .RN(net3),
    .CK(net1),
    .Q(net65),
    .QN(_089_));
 DFFR_X1 \dst_data_reg[6]$_DFFE_PN0P_  (.D(_062_),
    .RN(net3),
    .CK(net1),
    .Q(net66),
    .QN(_088_));
 DFFR_X1 \dst_data_reg[7]$_DFFE_PN0P_  (.D(_063_),
    .RN(net3),
    .CK(net1),
    .Q(net67),
    .QN(_087_));
 DFFR_X1 \dst_data_reg[8]$_DFFE_PN0P_  (.D(_064_),
    .RN(net3),
    .CK(net1),
    .Q(net68),
    .QN(_086_));
 DFFR_X1 \dst_data_reg[9]$_DFFE_PN0P_  (.D(_065_),
    .RN(net3),
    .CK(net1),
    .Q(net69),
    .QN(_085_));
 DFFR_X2 \dst_valid_reg$_DFFE_PN0P_  (.D(_066_),
    .RN(net3),
    .CK(net1),
    .Q(net70),
    .QN(_152_));
 DFFR_X1 \req_sync[0]$_DFF_PN0_  (.D(src_req),
    .RN(net3),
    .CK(net1),
    .Q(\req_sync[0] ),
    .QN(_153_));
 DFFR_X1 \req_sync[1]$_DFF_PN0_  (.D(\req_sync[0] ),
    .RN(net3),
    .CK(net1),
    .Q(dst_req),
    .QN(_084_));
 DFFR_X1 \src_req$_DFFE_PN0P_  (.D(_067_),
    .RN(net73),
    .CK(clknet_2_0__leaf_src_clk),
    .Q(src_req),
    .QN(_000_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_45 ();
 BUF_X4 input1 (.A(dst_clk),
    .Z(net1));
 BUF_X1 input2 (.A(dst_ready),
    .Z(net2));
 BUF_X8 input3 (.A(dst_rst_n),
    .Z(net3));
 BUF_X1 input4 (.A(src_data[0]),
    .Z(net4));
 BUF_X1 input5 (.A(src_data[10]),
    .Z(net5));
 BUF_X1 input6 (.A(src_data[11]),
    .Z(net6));
 BUF_X1 input7 (.A(src_data[12]),
    .Z(net7));
 BUF_X1 input8 (.A(src_data[13]),
    .Z(net8));
 BUF_X1 input9 (.A(src_data[14]),
    .Z(net9));
 BUF_X1 input10 (.A(src_data[15]),
    .Z(net10));
 BUF_X1 input11 (.A(src_data[16]),
    .Z(net11));
 BUF_X1 input12 (.A(src_data[17]),
    .Z(net12));
 BUF_X1 input13 (.A(src_data[18]),
    .Z(net13));
 BUF_X1 input14 (.A(src_data[19]),
    .Z(net14));
 BUF_X1 input15 (.A(src_data[1]),
    .Z(net15));
 BUF_X1 input16 (.A(src_data[20]),
    .Z(net16));
 BUF_X1 input17 (.A(src_data[21]),
    .Z(net17));
 BUF_X1 input18 (.A(src_data[22]),
    .Z(net18));
 BUF_X1 input19 (.A(src_data[23]),
    .Z(net19));
 BUF_X1 input20 (.A(src_data[24]),
    .Z(net20));
 BUF_X1 input21 (.A(src_data[25]),
    .Z(net21));
 BUF_X1 input22 (.A(src_data[26]),
    .Z(net22));
 BUF_X1 input23 (.A(src_data[27]),
    .Z(net23));
 BUF_X1 input24 (.A(src_data[28]),
    .Z(net24));
 BUF_X1 input25 (.A(src_data[29]),
    .Z(net25));
 BUF_X1 input26 (.A(src_data[2]),
    .Z(net26));
 BUF_X1 input27 (.A(src_data[30]),
    .Z(net27));
 BUF_X1 input28 (.A(src_data[31]),
    .Z(net28));
 BUF_X1 input29 (.A(src_data[3]),
    .Z(net29));
 BUF_X1 input30 (.A(src_data[4]),
    .Z(net30));
 BUF_X1 input31 (.A(src_data[5]),
    .Z(net31));
 BUF_X1 input32 (.A(src_data[6]),
    .Z(net32));
 BUF_X1 input33 (.A(src_data[7]),
    .Z(net33));
 BUF_X1 input34 (.A(src_data[8]),
    .Z(net34));
 BUF_X1 input35 (.A(src_data[9]),
    .Z(net35));
 BUF_X8 input36 (.A(net72),
    .Z(net36));
 BUF_X1 input37 (.A(src_valid),
    .Z(net37));
 BUF_X1 output38 (.A(net38),
    .Z(dst_data[0]));
 BUF_X1 output39 (.A(net39),
    .Z(dst_data[10]));
 BUF_X1 output40 (.A(net40),
    .Z(dst_data[11]));
 BUF_X1 output41 (.A(net41),
    .Z(dst_data[12]));
 BUF_X1 output42 (.A(net42),
    .Z(dst_data[13]));
 BUF_X1 output43 (.A(net43),
    .Z(dst_data[14]));
 BUF_X1 output44 (.A(net44),
    .Z(dst_data[15]));
 BUF_X1 output45 (.A(net45),
    .Z(dst_data[16]));
 BUF_X1 output46 (.A(net46),
    .Z(dst_data[17]));
 BUF_X1 output47 (.A(net47),
    .Z(dst_data[18]));
 BUF_X1 output48 (.A(net48),
    .Z(dst_data[19]));
 BUF_X1 output49 (.A(net49),
    .Z(dst_data[1]));
 BUF_X1 output50 (.A(net50),
    .Z(dst_data[20]));
 BUF_X1 output51 (.A(net51),
    .Z(dst_data[21]));
 BUF_X1 output52 (.A(net52),
    .Z(dst_data[22]));
 BUF_X1 output53 (.A(net53),
    .Z(dst_data[23]));
 BUF_X1 output54 (.A(net54),
    .Z(dst_data[24]));
 BUF_X1 output55 (.A(net55),
    .Z(dst_data[25]));
 BUF_X1 output56 (.A(net56),
    .Z(dst_data[26]));
 BUF_X1 output57 (.A(net57),
    .Z(dst_data[27]));
 BUF_X1 output58 (.A(net58),
    .Z(dst_data[28]));
 BUF_X1 output59 (.A(net59),
    .Z(dst_data[29]));
 BUF_X1 output60 (.A(net60),
    .Z(dst_data[2]));
 BUF_X1 output61 (.A(net61),
    .Z(dst_data[30]));
 BUF_X1 output62 (.A(net62),
    .Z(dst_data[31]));
 BUF_X1 output63 (.A(net63),
    .Z(dst_data[3]));
 BUF_X1 output64 (.A(net64),
    .Z(dst_data[4]));
 BUF_X1 output65 (.A(net65),
    .Z(dst_data[5]));
 BUF_X1 output66 (.A(net66),
    .Z(dst_data[6]));
 BUF_X1 output67 (.A(net67),
    .Z(dst_data[7]));
 BUF_X1 output68 (.A(net68),
    .Z(dst_data[8]));
 BUF_X1 output69 (.A(net69),
    .Z(dst_data[9]));
 BUF_X1 output70 (.A(net70),
    .Z(dst_valid));
 BUF_X1 output71 (.A(net71),
    .Z(src_ready));
 CLKBUF_X3 clkbuf_0_src_clk (.A(src_clk),
    .Z(clknet_0_src_clk));
 CLKBUF_X3 clkbuf_2_0__f_src_clk (.A(clknet_0_src_clk),
    .Z(clknet_2_0__leaf_src_clk));
 CLKBUF_X3 clkbuf_2_1__f_src_clk (.A(clknet_0_src_clk),
    .Z(clknet_2_1__leaf_src_clk));
 CLKBUF_X3 clkbuf_2_2__f_src_clk (.A(clknet_0_src_clk),
    .Z(clknet_2_2__leaf_src_clk));
 CLKBUF_X3 clkbuf_2_3__f_src_clk (.A(clknet_0_src_clk),
    .Z(clknet_2_3__leaf_src_clk));
 INV_X1 clkload0 (.A(clknet_2_0__leaf_src_clk));
 CLKBUF_X1 clkload1 (.A(clknet_2_1__leaf_src_clk));
 INV_X1 clkload2 (.A(clknet_2_3__leaf_src_clk));
 CLKBUF_X1 hold1 (.A(net74),
    .Z(net72));
 BUF_X8 hold2 (.A(net36),
    .Z(net73));
 CLKBUF_X1 hold3 (.A(src_rst_n),
    .Z(net74));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_33 ();
 FILLCELL_X2 FILLER_0_56 ();
 FILLCELL_X2 FILLER_0_96 ();
 FILLCELL_X2 FILLER_0_101 ();
 FILLCELL_X1 FILLER_0_103 ();
 FILLCELL_X4 FILLER_0_110 ();
 FILLCELL_X1 FILLER_0_114 ();
 FILLCELL_X8 FILLER_0_118 ();
 FILLCELL_X1 FILLER_0_126 ();
 FILLCELL_X8 FILLER_0_136 ();
 FILLCELL_X4 FILLER_0_144 ();
 FILLCELL_X2 FILLER_0_148 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X8 FILLER_1_17 ();
 FILLCELL_X2 FILLER_1_25 ();
 FILLCELL_X8 FILLER_1_52 ();
 FILLCELL_X1 FILLER_1_83 ();
 FILLCELL_X1 FILLER_1_91 ();
 FILLCELL_X2 FILLER_1_112 ();
 FILLCELL_X2 FILLER_1_134 ();
 FILLCELL_X8 FILLER_1_143 ();
 FILLCELL_X2 FILLER_1_151 ();
 FILLCELL_X2 FILLER_1_160 ();
 FILLCELL_X1 FILLER_1_162 ();
 FILLCELL_X4 FILLER_2_1 ();
 FILLCELL_X8 FILLER_2_52 ();
 FILLCELL_X2 FILLER_2_67 ();
 FILLCELL_X1 FILLER_2_69 ();
 FILLCELL_X2 FILLER_2_110 ();
 FILLCELL_X8 FILLER_2_159 ();
 FILLCELL_X2 FILLER_2_167 ();
 FILLCELL_X1 FILLER_2_169 ();
 FILLCELL_X2 FILLER_3_1 ();
 FILLCELL_X1 FILLER_3_3 ();
 FILLCELL_X4 FILLER_3_54 ();
 FILLCELL_X1 FILLER_3_92 ();
 FILLCELL_X8 FILLER_3_107 ();
 FILLCELL_X1 FILLER_3_115 ();
 FILLCELL_X1 FILLER_3_130 ();
 FILLCELL_X2 FILLER_3_151 ();
 FILLCELL_X1 FILLER_3_153 ();
 FILLCELL_X8 FILLER_4_1 ();
 FILLCELL_X2 FILLER_4_9 ();
 FILLCELL_X1 FILLER_4_11 ();
 FILLCELL_X8 FILLER_4_34 ();
 FILLCELL_X1 FILLER_4_42 ();
 FILLCELL_X32 FILLER_4_52 ();
 FILLCELL_X32 FILLER_4_84 ();
 FILLCELL_X16 FILLER_4_116 ();
 FILLCELL_X8 FILLER_4_132 ();
 FILLCELL_X4 FILLER_4_140 ();
 FILLCELL_X2 FILLER_4_164 ();
 FILLCELL_X1 FILLER_4_166 ();
 FILLCELL_X4 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_36 ();
 FILLCELL_X32 FILLER_5_68 ();
 FILLCELL_X32 FILLER_5_112 ();
 FILLCELL_X2 FILLER_5_144 ();
 FILLCELL_X4 FILLER_5_166 ();
 FILLCELL_X4 FILLER_6_1 ();
 FILLCELL_X1 FILLER_6_5 ();
 FILLCELL_X2 FILLER_6_9 ();
 FILLCELL_X1 FILLER_6_11 ();
 FILLCELL_X1 FILLER_6_28 ();
 FILLCELL_X4 FILLER_6_38 ();
 FILLCELL_X4 FILLER_6_69 ();
 FILLCELL_X2 FILLER_6_73 ();
 FILLCELL_X1 FILLER_6_75 ();
 FILLCELL_X2 FILLER_6_89 ();
 FILLCELL_X1 FILLER_6_91 ();
 FILLCELL_X16 FILLER_6_122 ();
 FILLCELL_X2 FILLER_6_138 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X8 FILLER_7_17 ();
 FILLCELL_X4 FILLER_7_25 ();
 FILLCELL_X2 FILLER_7_29 ();
 FILLCELL_X1 FILLER_7_31 ();
 FILLCELL_X16 FILLER_7_81 ();
 FILLCELL_X2 FILLER_7_97 ();
 FILLCELL_X1 FILLER_7_149 ();
 FILLCELL_X2 FILLER_8_1 ();
 FILLCELL_X4 FILLER_8_6 ();
 FILLCELL_X1 FILLER_8_30 ();
 FILLCELL_X2 FILLER_8_38 ();
 FILLCELL_X1 FILLER_8_40 ();
 FILLCELL_X8 FILLER_8_46 ();
 FILLCELL_X4 FILLER_8_54 ();
 FILLCELL_X1 FILLER_8_58 ();
 FILLCELL_X32 FILLER_8_72 ();
 FILLCELL_X8 FILLER_8_104 ();
 FILLCELL_X2 FILLER_8_112 ();
 FILLCELL_X1 FILLER_8_114 ();
 FILLCELL_X8 FILLER_8_129 ();
 FILLCELL_X2 FILLER_8_137 ();
 FILLCELL_X1 FILLER_8_139 ();
 FILLCELL_X1 FILLER_9_1 ();
 FILLCELL_X1 FILLER_9_5 ();
 FILLCELL_X1 FILLER_9_26 ();
 FILLCELL_X2 FILLER_9_30 ();
 FILLCELL_X32 FILLER_9_59 ();
 FILLCELL_X16 FILLER_9_91 ();
 FILLCELL_X8 FILLER_9_107 ();
 FILLCELL_X2 FILLER_9_115 ();
 FILLCELL_X1 FILLER_9_117 ();
 FILLCELL_X8 FILLER_9_138 ();
 FILLCELL_X4 FILLER_9_146 ();
 FILLCELL_X4 FILLER_9_157 ();
 FILLCELL_X2 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_37 ();
 FILLCELL_X16 FILLER_10_45 ();
 FILLCELL_X8 FILLER_10_61 ();
 FILLCELL_X4 FILLER_10_69 ();
 FILLCELL_X32 FILLER_10_86 ();
 FILLCELL_X32 FILLER_10_118 ();
 FILLCELL_X16 FILLER_10_150 ();
 FILLCELL_X4 FILLER_10_166 ();
 FILLCELL_X8 FILLER_11_41 ();
 FILLCELL_X2 FILLER_11_49 ();
 FILLCELL_X1 FILLER_11_51 ();
 FILLCELL_X8 FILLER_11_65 ();
 FILLCELL_X4 FILLER_11_73 ();
 FILLCELL_X1 FILLER_11_77 ();
 FILLCELL_X32 FILLER_11_91 ();
 FILLCELL_X16 FILLER_11_123 ();
 FILLCELL_X4 FILLER_11_139 ();
 FILLCELL_X2 FILLER_11_143 ();
 FILLCELL_X1 FILLER_11_145 ();
 FILLCELL_X1 FILLER_11_166 ();
 FILLCELL_X2 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_3 ();
 FILLCELL_X32 FILLER_12_7 ();
 FILLCELL_X32 FILLER_12_39 ();
 FILLCELL_X4 FILLER_12_71 ();
 FILLCELL_X2 FILLER_12_75 ();
 FILLCELL_X32 FILLER_12_82 ();
 FILLCELL_X1 FILLER_12_114 ();
 FILLCELL_X1 FILLER_12_135 ();
 FILLCELL_X2 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_30 ();
 FILLCELL_X2 FILLER_13_34 ();
 FILLCELL_X32 FILLER_13_56 ();
 FILLCELL_X8 FILLER_13_88 ();
 FILLCELL_X4 FILLER_13_96 ();
 FILLCELL_X2 FILLER_13_100 ();
 FILLCELL_X2 FILLER_13_109 ();
 FILLCELL_X1 FILLER_13_111 ();
 FILLCELL_X16 FILLER_13_119 ();
 FILLCELL_X1 FILLER_13_135 ();
 FILLCELL_X1 FILLER_13_169 ();
 FILLCELL_X2 FILLER_14_4 ();
 FILLCELL_X8 FILLER_14_43 ();
 FILLCELL_X4 FILLER_14_51 ();
 FILLCELL_X1 FILLER_14_55 ();
 FILLCELL_X16 FILLER_14_83 ();
 FILLCELL_X1 FILLER_14_99 ();
 FILLCELL_X16 FILLER_14_120 ();
 FILLCELL_X2 FILLER_14_136 ();
 FILLCELL_X1 FILLER_14_138 ();
 FILLCELL_X1 FILLER_14_166 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X16 FILLER_15_8 ();
 FILLCELL_X8 FILLER_15_24 ();
 FILLCELL_X4 FILLER_15_32 ();
 FILLCELL_X1 FILLER_15_39 ();
 FILLCELL_X32 FILLER_15_74 ();
 FILLCELL_X16 FILLER_15_106 ();
 FILLCELL_X8 FILLER_15_122 ();
 FILLCELL_X4 FILLER_15_130 ();
 FILLCELL_X2 FILLER_15_134 ();
 FILLCELL_X1 FILLER_15_136 ();
 FILLCELL_X1 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_35 ();
 FILLCELL_X2 FILLER_16_39 ();
 FILLCELL_X1 FILLER_16_41 ();
 FILLCELL_X32 FILLER_16_62 ();
 FILLCELL_X32 FILLER_16_94 ();
 FILLCELL_X8 FILLER_16_126 ();
 FILLCELL_X4 FILLER_16_134 ();
 FILLCELL_X1 FILLER_16_138 ();
 FILLCELL_X1 FILLER_16_166 ();
 FILLCELL_X2 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_3 ();
 FILLCELL_X4 FILLER_17_11 ();
 FILLCELL_X16 FILLER_17_35 ();
 FILLCELL_X32 FILLER_17_56 ();
 FILLCELL_X16 FILLER_17_88 ();
 FILLCELL_X8 FILLER_17_104 ();
 FILLCELL_X1 FILLER_17_112 ();
 FILLCELL_X16 FILLER_17_120 ();
 FILLCELL_X8 FILLER_17_136 ();
 FILLCELL_X2 FILLER_17_144 ();
 FILLCELL_X4 FILLER_17_166 ();
 FILLCELL_X16 FILLER_18_14 ();
 FILLCELL_X8 FILLER_18_30 ();
 FILLCELL_X4 FILLER_18_38 ();
 FILLCELL_X1 FILLER_18_42 ();
 FILLCELL_X2 FILLER_18_70 ();
 FILLCELL_X4 FILLER_18_112 ();
 FILLCELL_X1 FILLER_18_116 ();
 FILLCELL_X8 FILLER_18_124 ();
 FILLCELL_X4 FILLER_18_132 ();
 FILLCELL_X2 FILLER_18_136 ();
 FILLCELL_X1 FILLER_18_138 ();
 FILLCELL_X1 FILLER_18_146 ();
 FILLCELL_X2 FILLER_19_31 ();
 FILLCELL_X1 FILLER_19_33 ();
 FILLCELL_X2 FILLER_19_68 ();
 FILLCELL_X1 FILLER_19_70 ();
 FILLCELL_X2 FILLER_19_165 ();
 FILLCELL_X4 FILLER_20_54 ();
 FILLCELL_X1 FILLER_20_58 ();
 FILLCELL_X1 FILLER_20_79 ();
 FILLCELL_X1 FILLER_20_94 ();
 FILLCELL_X1 FILLER_20_115 ();
 FILLCELL_X2 FILLER_20_136 ();
 FILLCELL_X1 FILLER_20_138 ();
 FILLCELL_X16 FILLER_20_146 ();
 FILLCELL_X8 FILLER_20_162 ();
 FILLCELL_X2 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_10 ();
 FILLCELL_X4 FILLER_21_27 ();
 FILLCELL_X1 FILLER_21_31 ();
 FILLCELL_X8 FILLER_21_75 ();
 FILLCELL_X4 FILLER_21_83 ();
 FILLCELL_X2 FILLER_21_87 ();
 FILLCELL_X1 FILLER_21_110 ();
 FILLCELL_X2 FILLER_21_118 ();
 FILLCELL_X2 FILLER_21_167 ();
 FILLCELL_X1 FILLER_21_169 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_17 ();
 FILLCELL_X2 FILLER_22_28 ();
 FILLCELL_X4 FILLER_22_33 ();
 FILLCELL_X4 FILLER_22_40 ();
 FILLCELL_X1 FILLER_22_54 ();
 FILLCELL_X1 FILLER_22_58 ();
 FILLCELL_X2 FILLER_22_78 ();
 FILLCELL_X8 FILLER_22_83 ();
 FILLCELL_X4 FILLER_22_94 ();
 FILLCELL_X16 FILLER_22_116 ();
 FILLCELL_X1 FILLER_22_135 ();
 FILLCELL_X16 FILLER_22_142 ();
 FILLCELL_X8 FILLER_22_158 ();
 FILLCELL_X4 FILLER_22_166 ();
endmodule
