module configurable_prng (clk,
    enable,
    reseed,
    rst_n,
    valid,
    random,
    seed_in);
 input clk;
 input enable;
 input reseed;
 input rst_n;
 output valid;
 output [15:0] random;
 input [15:0] seed_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net36;

 sky130_fd_sc_hd__buf_2 _057_ (.A(reseed),
    .X(_023_));
 sky130_fd_sc_hd__nor4_1 _058_ (.A(net18),
    .B(net17),
    .C(net5),
    .D(net8),
    .Y(_024_));
 sky130_fd_sc_hd__nor4_1 _059_ (.A(net4),
    .B(net7),
    .C(net6),
    .D(net9),
    .Y(_025_));
 sky130_fd_sc_hd__nor4_1 _060_ (.A(net10),
    .B(net3),
    .C(net12),
    .D(net15),
    .Y(_026_));
 sky130_fd_sc_hd__nor4_1 _061_ (.A(net11),
    .B(net14),
    .C(net13),
    .D(net16),
    .Y(_027_));
 sky130_fd_sc_hd__nand4_1 _062_ (.A(_024_),
    .B(_025_),
    .C(_026_),
    .D(_027_),
    .Y(_028_));
 sky130_fd_sc_hd__nand2_4 _063_ (.A(_023_),
    .B(_028_),
    .Y(_029_));
 sky130_fd_sc_hd__buf_4 _064_ (.A(enable),
    .X(_030_));
 sky130_fd_sc_hd__buf_6 _065_ (.A(_030_),
    .X(_031_));
 sky130_fd_sc_hd__xnor2_1 _066_ (.A(net25),
    .B(net20),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_1 _067_ (.A(net23),
    .B(net22),
    .Y(_033_));
 sky130_fd_sc_hd__xnor2_1 _068_ (.A(_032_),
    .B(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__nor2_1 _069_ (.A(_030_),
    .B(net19),
    .Y(_035_));
 sky130_fd_sc_hd__a21oi_1 _070_ (.A1(_031_),
    .A2(_034_),
    .B1(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__buf_2 _071_ (.A(_023_),
    .X(_037_));
 sky130_fd_sc_hd__o22a_1 _072_ (.A1(net3),
    .A2(_029_),
    .B1(_036_),
    .B2(_037_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _073_ (.A0(net20),
    .A1(net34),
    .S(_030_),
    .X(_038_));
 sky130_fd_sc_hd__buf_2 _074_ (.A(_023_),
    .X(_039_));
 sky130_fd_sc_hd__o22a_1 _075_ (.A1(net4),
    .A2(_029_),
    .B1(_038_),
    .B2(_039_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _076_ (.A0(net21),
    .A1(net20),
    .S(_030_),
    .X(_040_));
 sky130_fd_sc_hd__o22a_1 _077_ (.A1(net5),
    .A2(_029_),
    .B1(_040_),
    .B2(_039_),
    .X(_002_));
 sky130_fd_sc_hd__mux2i_1 _078_ (.A0(net22),
    .A1(net21),
    .S(_031_),
    .Y(_041_));
 sky130_fd_sc_hd__nand2_1 _079_ (.A(_037_),
    .B(net6),
    .Y(_042_));
 sky130_fd_sc_hd__o21ai_0 _080_ (.A1(_039_),
    .A2(_041_),
    .B1(_042_),
    .Y(_003_));
 sky130_fd_sc_hd__mux2_1 _081_ (.A0(net23),
    .A1(net22),
    .S(_030_),
    .X(_043_));
 sky130_fd_sc_hd__o22a_1 _082_ (.A1(net7),
    .A2(_029_),
    .B1(_043_),
    .B2(_039_),
    .X(_004_));
 sky130_fd_sc_hd__mux2i_1 _083_ (.A0(net24),
    .A1(net23),
    .S(_031_),
    .Y(_044_));
 sky130_fd_sc_hd__nand2_1 _084_ (.A(_037_),
    .B(net8),
    .Y(_045_));
 sky130_fd_sc_hd__o21ai_0 _085_ (.A1(_039_),
    .A2(_044_),
    .B1(_045_),
    .Y(_005_));
 sky130_fd_sc_hd__mux2_1 _086_ (.A0(net25),
    .A1(net24),
    .S(_030_),
    .X(_046_));
 sky130_fd_sc_hd__o22a_1 _087_ (.A1(net9),
    .A2(_029_),
    .B1(_046_),
    .B2(_039_),
    .X(_006_));
 sky130_fd_sc_hd__mux2i_1 _088_ (.A0(net26),
    .A1(net19),
    .S(_031_),
    .Y(_047_));
 sky130_fd_sc_hd__nand2_1 _089_ (.A(_037_),
    .B(net10),
    .Y(_048_));
 sky130_fd_sc_hd__o21ai_0 _090_ (.A1(_039_),
    .A2(_047_),
    .B1(_048_),
    .Y(_007_));
 sky130_fd_sc_hd__mux2i_1 _091_ (.A0(net27),
    .A1(net26),
    .S(_031_),
    .Y(_049_));
 sky130_fd_sc_hd__nand2_1 _092_ (.A(_037_),
    .B(net11),
    .Y(_050_));
 sky130_fd_sc_hd__o21ai_0 _093_ (.A1(_023_),
    .A2(_049_),
    .B1(_050_),
    .Y(_008_));
 sky130_fd_sc_hd__mux2i_1 _094_ (.A0(net28),
    .A1(net27),
    .S(_031_),
    .Y(_051_));
 sky130_fd_sc_hd__nand2_1 _095_ (.A(_037_),
    .B(net12),
    .Y(_052_));
 sky130_fd_sc_hd__o21ai_0 _096_ (.A1(_023_),
    .A2(_051_),
    .B1(_052_),
    .Y(_009_));
 sky130_fd_sc_hd__mux2i_1 _097_ (.A0(net29),
    .A1(net28),
    .S(_031_),
    .Y(_053_));
 sky130_fd_sc_hd__nand2_1 _098_ (.A(_037_),
    .B(net13),
    .Y(_054_));
 sky130_fd_sc_hd__o21ai_0 _099_ (.A1(_023_),
    .A2(_053_),
    .B1(_054_),
    .Y(_010_));
 sky130_fd_sc_hd__mux2_1 _100_ (.A0(net30),
    .A1(net29),
    .S(_030_),
    .X(_055_));
 sky130_fd_sc_hd__o22a_1 _101_ (.A1(net14),
    .A2(_029_),
    .B1(_055_),
    .B2(_039_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _102_ (.A0(net31),
    .A1(net30),
    .S(_030_),
    .X(_056_));
 sky130_fd_sc_hd__o22a_1 _103_ (.A1(net15),
    .A2(_029_),
    .B1(_056_),
    .B2(_039_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _104_ (.A0(net32),
    .A1(net31),
    .S(_030_),
    .X(_017_));
 sky130_fd_sc_hd__o22a_1 _105_ (.A1(net16),
    .A2(_029_),
    .B1(_017_),
    .B2(_039_),
    .X(_013_));
 sky130_fd_sc_hd__mux2i_1 _106_ (.A0(net33),
    .A1(net32),
    .S(_031_),
    .Y(_018_));
 sky130_fd_sc_hd__nand2_1 _107_ (.A(_037_),
    .B(net17),
    .Y(_019_));
 sky130_fd_sc_hd__o21ai_0 _108_ (.A1(_023_),
    .A2(_018_),
    .B1(_019_),
    .Y(_014_));
 sky130_fd_sc_hd__mux2i_1 _109_ (.A0(net34),
    .A1(net33),
    .S(_031_),
    .Y(_020_));
 sky130_fd_sc_hd__nand2_1 _110_ (.A(_037_),
    .B(net18),
    .Y(_021_));
 sky130_fd_sc_hd__o21ai_0 _111_ (.A1(_023_),
    .A2(_020_),
    .B1(_021_),
    .Y(_015_));
 sky130_fd_sc_hd__nor2_1 _112_ (.A(_031_),
    .B(net35),
    .Y(_022_));
 sky130_fd_sc_hd__nor2_1 _113_ (.A(_037_),
    .B(_022_),
    .Y(_016_));
 sky130_fd_sc_hd__dfstp_1 \lfsr_reg[0]$_DFFE_PN1P_  (.D(_000_),
    .Q(net19),
    .SET_B(net2),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \lfsr_reg[10]$_DFFE_PN1P_  (.D(_001_),
    .Q(net20),
    .SET_B(net2),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \lfsr_reg[11]$_DFFE_PN1P_  (.D(_002_),
    .Q(net21),
    .SET_B(net2),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[12]$_DFFE_PN0P_  (.D(_003_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \lfsr_reg[13]$_DFFE_PN1P_  (.D(_004_),
    .Q(net23),
    .SET_B(net2),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[14]$_DFFE_PN0P_  (.D(_005_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \lfsr_reg[15]$_DFFE_PN1P_  (.D(_006_),
    .Q(net25),
    .SET_B(net2),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[1]$_DFFE_PN0P_  (.D(_007_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[2]$_DFFE_PN0P_  (.D(_008_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[3]$_DFFE_PN0P_  (.D(_009_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[4]$_DFFE_PN0P_  (.D(_010_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \lfsr_reg[5]$_DFFE_PN1P_  (.D(_011_),
    .Q(net30),
    .SET_B(net2),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \lfsr_reg[6]$_DFFE_PN1P_  (.D(_012_),
    .Q(net31),
    .SET_B(net2),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \lfsr_reg[7]$_DFFE_PN1P_  (.D(_013_),
    .Q(net32),
    .SET_B(net2),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[8]$_DFFE_PN0P_  (.D(_014_),
    .Q(net33),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[9]$_DFFE_PN0P_  (.D(_015_),
    .Q(net34),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_reg$_DFFE_PN0P_  (.D(_016_),
    .Q(net35),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 hold1 (.A(net2),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_71 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(net36),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(seed_in[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(seed_in[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(seed_in[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(seed_in[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(seed_in[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(seed_in[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(seed_in[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(seed_in[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(seed_in[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(seed_in[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(seed_in[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(seed_in[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(seed_in[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(seed_in[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(seed_in[8]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(seed_in[9]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(random[0]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(random[10]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(random[11]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(random[12]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(random[13]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(random[14]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(random[15]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(random[1]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(random[2]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(random[3]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(random[4]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(random[5]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(random[6]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(random[7]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(random[8]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(random[9]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(valid));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net36));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_159 ();
endmodule
