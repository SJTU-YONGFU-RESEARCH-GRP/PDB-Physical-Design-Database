module parameterized_decade_counter (clk,
    enable,
    rst_n,
    tc,
    count);
 input clk;
 input enable;
 input rst_n;
 output tc;
 output [3:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net8;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22_ (.I(net5),
    .ZN(_04_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23_ (.A1(net6),
    .A2(_18_),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24_ (.A1(_04_),
    .A2(_05_),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25_ (.I(net4),
    .ZN(_17_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26_ (.I(net2),
    .ZN(_06_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _27_ (.A1(_04_),
    .A2(_05_),
    .B(net3),
    .C(_06_),
    .ZN(_07_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28_ (.A1(_06_),
    .A2(net3),
    .Z(_08_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29_ (.A1(_07_),
    .A2(_08_),
    .Z(_00_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30_ (.A1(_04_),
    .A2(_05_),
    .B(_19_),
    .ZN(_09_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31_ (.I0(net4),
    .I1(_09_),
    .S(net2),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _32_ (.A1(net2),
    .A2(_20_),
    .ZN(_10_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _33_ (.A1(_05_),
    .A2(_10_),
    .ZN(_11_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _34_ (.I0(_10_),
    .I1(_11_),
    .S(_04_),
    .Z(_02_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _35_ (.A1(net2),
    .A2(net4),
    .A3(net3),
    .ZN(_12_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _36_ (.A1(net4),
    .A2(net3),
    .Z(_13_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _37_ (.I0(_12_),
    .I1(_13_),
    .S(net6),
    .Z(_14_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _38_ (.A1(net5),
    .A2(_18_),
    .B(net2),
    .ZN(_15_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _39_ (.A1(net6),
    .A2(_15_),
    .ZN(_16_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _40_ (.A1(_04_),
    .A2(_14_),
    .B(_16_),
    .ZN(_03_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _41_ (.A(net3),
    .B(_17_),
    .CO(_18_),
    .S(_19_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _42_ (.A(net3),
    .B(net4),
    .CO(_20_),
    .S(_21_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[0]$_DFFE_PN0P_  (.D(_00_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net3));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[1]$_DFFE_PN0P_  (.D(_01_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[2]$_DFFE_PN0P_  (.D(_02_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[3]$_DFFE_PN0P_  (.D(_03_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 hold1 (.I(net8),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_40 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_41 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_42 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_43 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_44 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_50 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input1 (.I(enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output2 (.I(net3),
    .Z(count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output3 (.I(net4),
    .Z(count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output4 (.I(net5),
    .Z(count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output5 (.I(net6),
    .Z(count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output6 (.I(net7),
    .Z(tc));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_184 ();
endmodule
