module arbiter_rr (active,
    clk,
    rst_n,
    grant,
    request);
 output active;
 input clk;
 input rst_n;
 output [3:0] grant;
 input [3:0] request;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire \priority_ptr[0] ;
 wire \priority_ptr[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net12;

 sky130_fd_sc_hd__buf_2 _056_ (.A(_049_),
    .X(_006_));
 sky130_fd_sc_hd__mux4_4 _057_ (.A0(net5),
    .A1(net4),
    .A2(net3),
    .A3(net2),
    .S0(\priority_ptr[0] ),
    .S1(_006_),
    .X(_007_));
 sky130_fd_sc_hd__buf_6 _058_ (.A(\priority_ptr[0] ),
    .X(_008_));
 sky130_fd_sc_hd__mux4_1 _059_ (.A0(net4),
    .A1(net5),
    .A2(net2),
    .A3(net3),
    .S0(_008_),
    .S1(\priority_ptr[1] ),
    .X(_009_));
 sky130_fd_sc_hd__nor2b_1 _060_ (.A(_007_),
    .B_N(_009_),
    .Y(_010_));
 sky130_fd_sc_hd__mux4_1 _061_ (.A0(net2),
    .A1(net3),
    .A2(net4),
    .A3(net5),
    .S0(_008_),
    .S1(\priority_ptr[1] ),
    .X(_011_));
 sky130_fd_sc_hd__buf_6 _062_ (.A(_011_),
    .X(_012_));
 sky130_fd_sc_hd__a221oi_1 _063_ (.A1(_052_),
    .A2(_007_),
    .B1(_010_),
    .B2(_050_),
    .C1(_012_),
    .Y(_013_));
 sky130_fd_sc_hd__nor2b_1 _064_ (.A(_048_),
    .B_N(_012_),
    .Y(_014_));
 sky130_fd_sc_hd__mux4_1 _065_ (.A0(net3),
    .A1(net5),
    .A2(net2),
    .A3(net4),
    .S0(_006_),
    .S1(_008_),
    .X(_015_));
 sky130_fd_sc_hd__nor4b_2 _066_ (.A(_012_),
    .B(_007_),
    .C(_009_),
    .D_N(_015_),
    .Y(_016_));
 sky130_fd_sc_hd__nand2_1 _067_ (.A(_054_),
    .B(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__o21ai_0 _068_ (.A1(_013_),
    .A2(_014_),
    .B1(_017_),
    .Y(_000_));
 sky130_fd_sc_hd__a221oi_1 _069_ (.A1(_050_),
    .A2(_007_),
    .B1(_010_),
    .B2(_054_),
    .C1(_012_),
    .Y(_018_));
 sky130_fd_sc_hd__nor2b_1 _070_ (.A(_052_),
    .B_N(_012_),
    .Y(_019_));
 sky130_fd_sc_hd__nand2_1 _071_ (.A(_048_),
    .B(_016_),
    .Y(_020_));
 sky130_fd_sc_hd__o21ai_0 _072_ (.A1(_018_),
    .A2(_019_),
    .B1(_020_),
    .Y(_001_));
 sky130_fd_sc_hd__a221oi_1 _073_ (.A1(_054_),
    .A2(_007_),
    .B1(_010_),
    .B2(_048_),
    .C1(_012_),
    .Y(_021_));
 sky130_fd_sc_hd__nor2b_1 _074_ (.A(_050_),
    .B_N(_012_),
    .Y(_022_));
 sky130_fd_sc_hd__nand2_1 _075_ (.A(_052_),
    .B(_016_),
    .Y(_023_));
 sky130_fd_sc_hd__o21ai_0 _076_ (.A1(_021_),
    .A2(_022_),
    .B1(_023_),
    .Y(_002_));
 sky130_fd_sc_hd__a221oi_1 _077_ (.A1(_048_),
    .A2(_007_),
    .B1(_010_),
    .B2(_052_),
    .C1(_012_),
    .Y(_024_));
 sky130_fd_sc_hd__nor2b_1 _078_ (.A(_054_),
    .B_N(_012_),
    .Y(_025_));
 sky130_fd_sc_hd__nand2_1 _079_ (.A(_050_),
    .B(_016_),
    .Y(_026_));
 sky130_fd_sc_hd__o21ai_0 _080_ (.A1(_024_),
    .A2(_025_),
    .B1(_026_),
    .Y(_003_));
 sky130_fd_sc_hd__inv_1 _081_ (.A(_008_),
    .Y(_046_));
 sky130_fd_sc_hd__inv_1 _082_ (.A(\priority_ptr[1] ),
    .Y(_047_));
 sky130_fd_sc_hd__nor2_1 _083_ (.A(_012_),
    .B(_010_),
    .Y(_027_));
 sky130_fd_sc_hd__xnor2_1 _084_ (.A(_008_),
    .B(_027_),
    .Y(_004_));
 sky130_fd_sc_hd__mux2_1 _085_ (.A0(net5),
    .A1(net3),
    .S(_006_),
    .X(_028_));
 sky130_fd_sc_hd__mux2i_1 _086_ (.A0(net4),
    .A1(net2),
    .S(_006_),
    .Y(_029_));
 sky130_fd_sc_hd__nor3b_1 _087_ (.A(net5),
    .B(\priority_ptr[1] ),
    .C_N(_008_),
    .Y(_030_));
 sky130_fd_sc_hd__a221oi_2 _088_ (.A1(_046_),
    .A2(_028_),
    .B1(_029_),
    .B2(_030_),
    .C1(_011_),
    .Y(_031_));
 sky130_fd_sc_hd__or4_1 _089_ (.A(net2),
    .B(net3),
    .C(net4),
    .D(net5),
    .X(_032_));
 sky130_fd_sc_hd__nand2_1 _090_ (.A(_006_),
    .B(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__nor2_1 _091_ (.A(_031_),
    .B(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__inv_1 _092_ (.A(_006_),
    .Y(_035_));
 sky130_fd_sc_hd__nor2_1 _093_ (.A(\priority_ptr[1] ),
    .B(_032_),
    .Y(_036_));
 sky130_fd_sc_hd__a31o_1 _094_ (.A1(net3),
    .A2(_035_),
    .A3(_031_),
    .B1(_036_),
    .X(_037_));
 sky130_fd_sc_hd__and2b_1 _095_ (.A_N(_008_),
    .B(net5),
    .X(_038_));
 sky130_fd_sc_hd__a2111o_1 _096_ (.A1(_008_),
    .A2(_035_),
    .B1(_038_),
    .C1(_047_),
    .D1(net2),
    .X(_039_));
 sky130_fd_sc_hd__nor2_1 _097_ (.A(net4),
    .B(_006_),
    .Y(_040_));
 sky130_fd_sc_hd__nor4_1 _098_ (.A(_008_),
    .B(net4),
    .C(net5),
    .D(\priority_ptr[1] ),
    .Y(_041_));
 sky130_fd_sc_hd__a31oi_1 _099_ (.A1(_008_),
    .A2(\priority_ptr[1] ),
    .A3(_040_),
    .B1(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__nand3b_1 _100_ (.A_N(net3),
    .B(_006_),
    .C(_032_),
    .Y(_043_));
 sky130_fd_sc_hd__a21oi_1 _101_ (.A1(_039_),
    .A2(_042_),
    .B1(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__nand4_1 _102_ (.A(_035_),
    .B(_031_),
    .C(_039_),
    .D(_042_),
    .Y(_045_));
 sky130_fd_sc_hd__nor4b_1 _103_ (.A(_034_),
    .B(_037_),
    .C(_044_),
    .D_N(_045_),
    .Y(_005_));
 sky130_fd_sc_hd__or4_1 _104_ (.A(net9),
    .B(net8),
    .C(net11),
    .D(net10),
    .X(net7));
 sky130_fd_sc_hd__ha_1 _105_ (.A(_046_),
    .B(_047_),
    .COUT(_048_),
    .SUM(_049_));
 sky130_fd_sc_hd__ha_1 _106_ (.A(_046_),
    .B(\priority_ptr[1] ),
    .COUT(_050_),
    .SUM(_051_));
 sky130_fd_sc_hd__ha_1 _107_ (.A(\priority_ptr[0] ),
    .B(_047_),
    .COUT(_052_),
    .SUM(_053_));
 sky130_fd_sc_hd__ha_1 _108_ (.A(\priority_ptr[0] ),
    .B(\priority_ptr[1] ),
    .COUT(_054_),
    .SUM(_055_));
 sky130_fd_sc_hd__dfrtp_1 \grant[0]$_DFF_PN0_  (.D(_000_),
    .Q(net8),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \grant[1]$_DFF_PN0_  (.D(_001_),
    .Q(net9),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \grant[2]$_DFF_PN0_  (.D(_002_),
    .Q(net10),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \grant[3]$_DFF_PN0_  (.D(_003_),
    .Q(net11),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfstp_1 \priority_ptr[0]$_DFFE_PN1P_  (.D(_004_),
    .Q(\priority_ptr[0] ),
    .SET_B(net6),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfstp_2 \priority_ptr[1]$_DFFE_PN1P_  (.D(_005_),
    .Q(\priority_ptr[1] ),
    .SET_B(net6),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1 (.A(net6),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_49 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(request[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(request[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(request[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(request[3]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(net12),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 output6 (.A(net7),
    .X(active));
 sky130_fd_sc_hd__clkbuf_1 output7 (.A(net8),
    .X(grant[0]));
 sky130_fd_sc_hd__clkbuf_1 output8 (.A(net9),
    .X(grant[1]));
 sky130_fd_sc_hd__clkbuf_1 output9 (.A(net10),
    .X(grant[2]));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net11),
    .X(grant[3]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net12));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_137 ();
endmodule
