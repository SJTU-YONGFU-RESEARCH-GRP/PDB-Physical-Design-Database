module parameterized_decade_counter (clk,
    enable,
    rst_n,
    tc,
    count);
 input clk;
 input enable;
 input rst_n;
 output tc;
 output [3:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X2 _26_ (.A(net4),
    .Z(_05_));
 NAND2_X1 _27_ (.A1(net5),
    .A2(_22_),
    .ZN(_06_));
 NOR2_X1 _28_ (.A1(_05_),
    .A2(_06_),
    .ZN(net6));
 INV_X1 _29_ (.A(net1),
    .ZN(_07_));
 BUF_X4 _30_ (.A(enable),
    .Z(_08_));
 NAND2_X1 _31_ (.A1(_08_),
    .A2(_00_),
    .ZN(_09_));
 INV_X1 _32_ (.A(_08_),
    .ZN(_10_));
 NAND2_X1 _33_ (.A1(_10_),
    .A2(net2),
    .ZN(_11_));
 AOI221_X1 _34_ (.A(_07_),
    .B1(_09_),
    .B2(_11_),
    .C1(net6),
    .C2(_08_),
    .ZN(_01_));
 NOR3_X2 _35_ (.A1(_05_),
    .A2(_10_),
    .A3(_06_),
    .ZN(_12_));
 NAND2_X1 _36_ (.A1(_08_),
    .A2(_23_),
    .ZN(_13_));
 OAI21_X1 _37_ (.A(_13_),
    .B1(net3),
    .B2(_08_),
    .ZN(_14_));
 NOR3_X1 _38_ (.A1(_07_),
    .A2(_12_),
    .A3(_14_),
    .ZN(_02_));
 NAND2_X1 _39_ (.A1(_08_),
    .A2(_24_),
    .ZN(_15_));
 XOR2_X1 _40_ (.A(_05_),
    .B(_15_),
    .Z(_16_));
 NOR3_X1 _41_ (.A1(_07_),
    .A2(_12_),
    .A3(_16_),
    .ZN(_03_));
 NAND4_X1 _42_ (.A1(_05_),
    .A2(_08_),
    .A3(net3),
    .A4(net2),
    .ZN(_17_));
 XOR2_X1 _43_ (.A(net5),
    .B(_17_),
    .Z(_18_));
 NOR3_X1 _44_ (.A1(_07_),
    .A2(_12_),
    .A3(_18_),
    .ZN(_04_));
 HA_X1 _45_ (.A(net2),
    .B(_21_),
    .CO(_22_),
    .S(_23_));
 HA_X1 _46_ (.A(net2),
    .B(net3),
    .CO(_24_),
    .S(_25_));
 DFF_X2 \count[0]$_SDFFE_PP0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net2),
    .QN(_00_));
 DFF_X2 \count[1]$_SDFFE_PP0P_  (.D(_02_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net3),
    .QN(_21_));
 DFF_X1 \count[2]$_SDFFE_PP0P_  (.D(_03_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net4),
    .QN(_20_));
 DFF_X1 \count[3]$_SDFFE_PP0P_  (.D(_04_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net5),
    .QN(_19_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_41 ();
 BUF_X1 input1 (.A(rst_n),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(count[0]));
 BUF_X1 output3 (.A(net3),
    .Z(count[1]));
 BUF_X1 output4 (.A(net4),
    .Z(count[2]));
 BUF_X1 output5 (.A(net5),
    .Z(count[3]));
 BUF_X1 output6 (.A(net6),
    .Z(tc));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X4 FILLER_0_71 ();
 FILLCELL_X1 FILLER_0_75 ();
 FILLCELL_X8 FILLER_0_81 ();
 FILLCELL_X8 FILLER_0_92 ();
 FILLCELL_X4 FILLER_0_100 ();
 FILLCELL_X1 FILLER_0_104 ();
 FILLCELL_X32 FILLER_0_112 ();
 FILLCELL_X16 FILLER_0_144 ();
 FILLCELL_X2 FILLER_0_160 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X4 FILLER_1_65 ();
 FILLCELL_X8 FILLER_1_71 ();
 FILLCELL_X4 FILLER_1_79 ();
 FILLCELL_X1 FILLER_1_83 ();
 FILLCELL_X32 FILLER_1_96 ();
 FILLCELL_X32 FILLER_1_128 ();
 FILLCELL_X2 FILLER_1_160 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X4 FILLER_2_49 ();
 FILLCELL_X2 FILLER_2_53 ();
 FILLCELL_X1 FILLER_2_55 ();
 FILLCELL_X2 FILLER_2_77 ();
 FILLCELL_X32 FILLER_2_100 ();
 FILLCELL_X16 FILLER_2_132 ();
 FILLCELL_X8 FILLER_2_148 ();
 FILLCELL_X4 FILLER_2_156 ();
 FILLCELL_X2 FILLER_2_160 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_65 ();
 FILLCELL_X4 FILLER_3_73 ();
 FILLCELL_X1 FILLER_3_77 ();
 FILLCELL_X32 FILLER_3_111 ();
 FILLCELL_X16 FILLER_3_143 ();
 FILLCELL_X2 FILLER_3_159 ();
 FILLCELL_X1 FILLER_3_161 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X16 FILLER_4_65 ();
 FILLCELL_X8 FILLER_4_81 ();
 FILLCELL_X2 FILLER_4_89 ();
 FILLCELL_X32 FILLER_4_96 ();
 FILLCELL_X32 FILLER_4_128 ();
 FILLCELL_X2 FILLER_4_160 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X8 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_84 ();
 FILLCELL_X1 FILLER_5_88 ();
 FILLCELL_X16 FILLER_5_99 ();
 FILLCELL_X8 FILLER_5_115 ();
 FILLCELL_X32 FILLER_5_126 ();
 FILLCELL_X4 FILLER_5_158 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X16 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_49 ();
 FILLCELL_X2 FILLER_6_57 ();
 FILLCELL_X4 FILLER_6_84 ();
 FILLCELL_X2 FILLER_6_88 ();
 FILLCELL_X1 FILLER_6_90 ();
 FILLCELL_X32 FILLER_6_98 ();
 FILLCELL_X32 FILLER_6_130 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_65 ();
 FILLCELL_X4 FILLER_7_73 ();
 FILLCELL_X32 FILLER_7_96 ();
 FILLCELL_X32 FILLER_7_128 ();
 FILLCELL_X2 FILLER_7_160 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X16 FILLER_8_97 ();
 FILLCELL_X8 FILLER_8_113 ();
 FILLCELL_X2 FILLER_8_121 ();
 FILLCELL_X32 FILLER_8_126 ();
 FILLCELL_X4 FILLER_8_158 ();
 FILLCELL_X4 FILLER_9_1 ();
 FILLCELL_X1 FILLER_9_5 ();
 FILLCELL_X32 FILLER_9_9 ();
 FILLCELL_X32 FILLER_9_41 ();
 FILLCELL_X32 FILLER_9_73 ();
 FILLCELL_X32 FILLER_9_105 ();
 FILLCELL_X16 FILLER_9_137 ();
 FILLCELL_X8 FILLER_9_153 ();
 FILLCELL_X1 FILLER_9_161 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X8 FILLER_10_65 ();
 FILLCELL_X4 FILLER_10_73 ();
 FILLCELL_X32 FILLER_10_82 ();
 FILLCELL_X32 FILLER_10_114 ();
 FILLCELL_X16 FILLER_10_146 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X1 FILLER_11_161 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X1 FILLER_12_161 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X1 FILLER_13_161 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X1 FILLER_14_161 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X1 FILLER_15_161 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X1 FILLER_16_161 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X1 FILLER_17_161 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X1 FILLER_18_161 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X1 FILLER_19_161 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X1 FILLER_20_161 ();
endmodule
