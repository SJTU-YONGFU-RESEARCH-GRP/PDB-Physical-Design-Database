module configurable_carry_lookahead_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 sky130_fd_sc_hd__inv_1 _070_ (.A(net65),
    .Y(_000_));
 sky130_fd_sc_hd__inv_1 _071_ (.A(net25),
    .Y(_052_));
 sky130_fd_sc_hd__inv_1 _072_ (.A(net1),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _073_ (.A(net57),
    .Y(_053_));
 sky130_fd_sc_hd__inv_1 _074_ (.A(net33),
    .Y(_002_));
 sky130_fd_sc_hd__inv_1 _075_ (.A(_006_),
    .Y(net68));
 sky130_fd_sc_hd__inv_1 _076_ (.A(_008_),
    .Y(net69));
 sky130_fd_sc_hd__inv_1 _077_ (.A(_010_),
    .Y(net70));
 sky130_fd_sc_hd__inv_1 _078_ (.A(_012_),
    .Y(net71));
 sky130_fd_sc_hd__inv_1 _079_ (.A(_014_),
    .Y(net72));
 sky130_fd_sc_hd__inv_1 _080_ (.A(_016_),
    .Y(net73));
 sky130_fd_sc_hd__inv_4 _081_ (.A(_018_),
    .Y(net74));
 sky130_fd_sc_hd__inv_1 _082_ (.A(_020_),
    .Y(net75));
 sky130_fd_sc_hd__inv_1 _083_ (.A(_022_),
    .Y(net76));
 sky130_fd_sc_hd__inv_1 _084_ (.A(_024_),
    .Y(net77));
 sky130_fd_sc_hd__inv_1 _085_ (.A(_027_),
    .Y(net78));
 sky130_fd_sc_hd__inv_1 _086_ (.A(_029_),
    .Y(net79));
 sky130_fd_sc_hd__inv_1 _087_ (.A(_031_),
    .Y(net80));
 sky130_fd_sc_hd__inv_1 _088_ (.A(_033_),
    .Y(net81));
 sky130_fd_sc_hd__inv_1 _089_ (.A(_035_),
    .Y(net82));
 sky130_fd_sc_hd__inv_1 _090_ (.A(_037_),
    .Y(net83));
 sky130_fd_sc_hd__inv_1 _091_ (.A(_039_),
    .Y(net84));
 sky130_fd_sc_hd__inv_1 _092_ (.A(_041_),
    .Y(net85));
 sky130_fd_sc_hd__inv_1 _093_ (.A(_043_),
    .Y(net86));
 sky130_fd_sc_hd__inv_1 _094_ (.A(_045_),
    .Y(net87));
 sky130_fd_sc_hd__inv_1 _095_ (.A(_047_),
    .Y(net88));
 sky130_fd_sc_hd__inv_1 _096_ (.A(_049_),
    .Y(net89));
 sky130_fd_sc_hd__inv_1 _097_ (.A(_051_),
    .Y(net90));
 sky130_fd_sc_hd__inv_1 _098_ (.A(_056_),
    .Y(net91));
 sky130_fd_sc_hd__inv_1 _099_ (.A(_058_),
    .Y(net92));
 sky130_fd_sc_hd__inv_1 _100_ (.A(_060_),
    .Y(net93));
 sky130_fd_sc_hd__inv_1 _101_ (.A(_062_),
    .Y(net94));
 sky130_fd_sc_hd__inv_1 _102_ (.A(_064_),
    .Y(net95));
 sky130_fd_sc_hd__inv_1 _103_ (.A(_066_),
    .Y(net96));
 sky130_fd_sc_hd__inv_1 _104_ (.A(_068_),
    .Y(net97));
 sky130_fd_sc_hd__inv_1 _105_ (.A(_069_),
    .Y(net98));
 sky130_fd_sc_hd__inv_1 _106_ (.A(_050_),
    .Y(_054_));
 sky130_fd_sc_hd__inv_1 _107_ (.A(_055_),
    .Y(net66));
 sky130_fd_sc_hd__inv_1 _108_ (.A(_003_),
    .Y(_025_));
 sky130_fd_sc_hd__fa_1 _109_ (.A(_000_),
    .B(_001_),
    .CIN(_002_),
    .COUT(_003_),
    .SUM(net67));
 sky130_fd_sc_hd__fa_1 _110_ (.A(net2),
    .B(net34),
    .CIN(_004_),
    .COUT(_005_),
    .SUM(_006_));
 sky130_fd_sc_hd__fa_1 _111_ (.A(net3),
    .B(net35),
    .CIN(_005_),
    .COUT(_007_),
    .SUM(_008_));
 sky130_fd_sc_hd__fa_1 _112_ (.A(net4),
    .B(net36),
    .CIN(_007_),
    .COUT(_009_),
    .SUM(_010_));
 sky130_fd_sc_hd__fa_1 _113_ (.A(net5),
    .B(net37),
    .CIN(_009_),
    .COUT(_011_),
    .SUM(_012_));
 sky130_fd_sc_hd__fa_1 _114_ (.A(net6),
    .B(net38),
    .CIN(_011_),
    .COUT(_013_),
    .SUM(_014_));
 sky130_fd_sc_hd__fa_4 _115_ (.A(net7),
    .B(net39),
    .CIN(_013_),
    .COUT(_015_),
    .SUM(_016_));
 sky130_fd_sc_hd__fa_1 _116_ (.A(net8),
    .B(net40),
    .CIN(_015_),
    .COUT(_017_),
    .SUM(_018_));
 sky130_fd_sc_hd__fa_1 _117_ (.A(net9),
    .B(net41),
    .CIN(_017_),
    .COUT(_019_),
    .SUM(_020_));
 sky130_fd_sc_hd__fa_1 _118_ (.A(net10),
    .B(net42),
    .CIN(_019_),
    .COUT(_021_),
    .SUM(_022_));
 sky130_fd_sc_hd__fa_1 _119_ (.A(net11),
    .B(net43),
    .CIN(_021_),
    .COUT(_023_),
    .SUM(_024_));
 sky130_fd_sc_hd__fa_1 _120_ (.A(net12),
    .B(net44),
    .CIN(_025_),
    .COUT(_026_),
    .SUM(_027_));
 sky130_fd_sc_hd__fa_1 _121_ (.A(net13),
    .B(net45),
    .CIN(_023_),
    .COUT(_028_),
    .SUM(_029_));
 sky130_fd_sc_hd__fa_1 _122_ (.A(net14),
    .B(net46),
    .CIN(_028_),
    .COUT(_030_),
    .SUM(_031_));
 sky130_fd_sc_hd__fa_1 _123_ (.A(net15),
    .B(net47),
    .CIN(_030_),
    .COUT(_032_),
    .SUM(_033_));
 sky130_fd_sc_hd__fa_1 _124_ (.A(net16),
    .B(net48),
    .CIN(_032_),
    .COUT(_034_),
    .SUM(_035_));
 sky130_fd_sc_hd__fa_1 _125_ (.A(net17),
    .B(net49),
    .CIN(_034_),
    .COUT(_036_),
    .SUM(_037_));
 sky130_fd_sc_hd__fa_1 _126_ (.A(net18),
    .B(net50),
    .CIN(_036_),
    .COUT(_038_),
    .SUM(_039_));
 sky130_fd_sc_hd__fa_1 _127_ (.A(net19),
    .B(net51),
    .CIN(_038_),
    .COUT(_040_),
    .SUM(_041_));
 sky130_fd_sc_hd__fa_1 _128_ (.A(net20),
    .B(net52),
    .CIN(_040_),
    .COUT(_042_),
    .SUM(_043_));
 sky130_fd_sc_hd__fa_1 _129_ (.A(net21),
    .B(net53),
    .CIN(_042_),
    .COUT(_044_),
    .SUM(_045_));
 sky130_fd_sc_hd__fa_1 _130_ (.A(net22),
    .B(net54),
    .CIN(_044_),
    .COUT(_046_),
    .SUM(_047_));
 sky130_fd_sc_hd__fa_1 _131_ (.A(net23),
    .B(net55),
    .CIN(_026_),
    .COUT(_048_),
    .SUM(_049_));
 sky130_fd_sc_hd__fa_1 _132_ (.A(net24),
    .B(net56),
    .CIN(_046_),
    .COUT(_050_),
    .SUM(_051_));
 sky130_fd_sc_hd__fa_1 _133_ (.A(_052_),
    .B(_053_),
    .CIN(_054_),
    .COUT(_055_),
    .SUM(_056_));
 sky130_fd_sc_hd__fa_1 _134_ (.A(net26),
    .B(net58),
    .CIN(_048_),
    .COUT(_057_),
    .SUM(_058_));
 sky130_fd_sc_hd__fa_1 _135_ (.A(net27),
    .B(net59),
    .CIN(_057_),
    .COUT(_059_),
    .SUM(_060_));
 sky130_fd_sc_hd__fa_1 _136_ (.A(net28),
    .B(net60),
    .CIN(_059_),
    .COUT(_061_),
    .SUM(_062_));
 sky130_fd_sc_hd__fa_1 _137_ (.A(net29),
    .B(net61),
    .CIN(_061_),
    .COUT(_063_),
    .SUM(_064_));
 sky130_fd_sc_hd__fa_1 _138_ (.A(net30),
    .B(net62),
    .CIN(_063_),
    .COUT(_065_),
    .SUM(_066_));
 sky130_fd_sc_hd__fa_1 _139_ (.A(net31),
    .B(net63),
    .CIN(_065_),
    .COUT(_067_),
    .SUM(_068_));
 sky130_fd_sc_hd__fa_1 _140_ (.A(net32),
    .B(net64),
    .CIN(_067_),
    .COUT(_004_),
    .SUM(_069_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1889 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(cin),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(cout));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(sum[0]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(sum[10]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(sum[11]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(sum[12]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(sum[13]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(sum[14]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(sum[15]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(sum[16]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(sum[17]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(sum[18]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(sum[19]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(sum[1]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(sum[20]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(sum[21]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(sum[22]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(sum[23]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(sum[24]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(sum[25]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .X(sum[26]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .X(sum[27]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(sum[28]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(sum[29]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(sum[2]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .X(sum[30]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .X(sum[31]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(sum[3]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .X(sum[4]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .X(sum[5]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(sum[6]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .X(sum[7]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .X(sum[8]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .X(sum[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_015_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_819 ();
endmodule
