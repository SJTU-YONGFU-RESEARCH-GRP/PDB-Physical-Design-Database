module pipelined_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    rd_en,
    rst_n,
    wr_en,
    data_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input rd_en;
 input rst_n;
 input wr_en;
 output [4:0] data_count;
 output [31:0] rd_data;
 input [31:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire clknet_0_clk;
 wire \pipeline_count[0] ;
 wire \pipeline_count[1] ;
 wire \pipeline_count[2] ;
 wire \pipeline_count[3] ;
 wire \pipeline_count[4] ;
 wire rd_en_pipe;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_en_pipe[0] ;
 wire \wr_en_pipe[1] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net45;

 sky130_fd_sc_hd__inv_1 _115_ (.A(_077_),
    .Y(_079_));
 sky130_fd_sc_hd__nand3_1 _116_ (.A(_109_),
    .B(_112_),
    .C(_076_),
    .Y(_062_));
 sky130_fd_sc_hd__a21oi_1 _117_ (.A1(_112_),
    .A2(_108_),
    .B1(_111_),
    .Y(_063_));
 sky130_fd_sc_hd__xnor2_1 _118_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .Y(_064_));
 sky130_fd_sc_hd__a21oi_1 _119_ (.A1(_062_),
    .A2(_063_),
    .B1(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__and3_1 _120_ (.A(_062_),
    .B(_063_),
    .C(_064_),
    .X(_066_));
 sky130_fd_sc_hd__or2_0 _121_ (.A(_065_),
    .B(_066_),
    .X(_067_));
 sky130_fd_sc_hd__buf_2 _122_ (.A(_067_),
    .X(_068_));
 sky130_fd_sc_hd__or4_1 _123_ (.A(\pipeline_count[1] ),
    .B(\pipeline_count[3] ),
    .C(\pipeline_count[2] ),
    .D(\pipeline_count[4] ),
    .X(_069_));
 sky130_fd_sc_hd__nand3b_1 _124_ (.A_N(_103_),
    .B(_106_),
    .C(_109_),
    .Y(_070_));
 sky130_fd_sc_hd__a21oi_1 _125_ (.A1(_109_),
    .A2(_105_),
    .B1(_108_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_1 _126_ (.A(_112_),
    .Y(_021_));
 sky130_fd_sc_hd__a21oi_1 _127_ (.A1(_070_),
    .A2(_020_),
    .B1(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__and3b_1 _128_ (.A_N(_103_),
    .B(_106_),
    .C(_109_),
    .X(_023_));
 sky130_fd_sc_hd__a21o_1 _129_ (.A1(_109_),
    .A2(_105_),
    .B1(_108_),
    .X(_024_));
 sky130_fd_sc_hd__nor3_1 _130_ (.A(_112_),
    .B(_023_),
    .C(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__nor2_1 _131_ (.A(_022_),
    .B(_025_),
    .Y(_092_));
 sky130_fd_sc_hd__xor2_2 _132_ (.A(_109_),
    .B(_076_),
    .X(_089_));
 sky130_fd_sc_hd__nand2_1 _133_ (.A(_104_),
    .B(_079_),
    .Y(_026_));
 sky130_fd_sc_hd__nor3_2 _134_ (.A(\pipeline_count[0] ),
    .B(_089_),
    .C(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__nor4b_1 _135_ (.A(_068_),
    .B(_069_),
    .C(_092_),
    .D_N(_027_),
    .Y(net11));
 sky130_fd_sc_hd__a211o_1 _136_ (.A1(_070_),
    .A2(_020_),
    .B1(_021_),
    .C1(_069_),
    .X(_028_));
 sky130_fd_sc_hd__or4_1 _137_ (.A(_112_),
    .B(_069_),
    .C(_023_),
    .D(_024_),
    .X(_029_));
 sky130_fd_sc_hd__a211oi_2 _138_ (.A1(_028_),
    .A2(_029_),
    .B1(_065_),
    .C1(_066_),
    .Y(_030_));
 sky130_fd_sc_hd__inv_1 _139_ (.A(net2),
    .Y(_031_));
 sky130_fd_sc_hd__a21o_1 _140_ (.A1(_027_),
    .A2(_030_),
    .B1(_031_),
    .X(_032_));
 sky130_fd_sc_hd__inv_1 _141_ (.A(_032_),
    .Y(_000_));
 sky130_fd_sc_hd__nor4b_4 _142_ (.A(_079_),
    .B(_022_),
    .C(_025_),
    .D_N(_089_),
    .Y(_033_));
 sky130_fd_sc_hd__or2_0 _143_ (.A(_068_),
    .B(_033_),
    .X(net12));
 sky130_fd_sc_hd__nor3b_2 _144_ (.A(_033_),
    .B(_068_),
    .C_N(net3),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _145_ (.A(\pipeline_count[1] ),
    .Y(_078_));
 sky130_fd_sc_hd__inv_1 _146_ (.A(_083_),
    .Y(_080_));
 sky130_fd_sc_hd__inv_1 _147_ (.A(_082_),
    .Y(net7));
 sky130_fd_sc_hd__inv_1 _148_ (.A(rd_en_pipe),
    .Y(_084_));
 sky130_fd_sc_hd__inv_1 _149_ (.A(\rd_ptr[1] ),
    .Y(_074_));
 sky130_fd_sc_hd__inv_1 _150_ (.A(_103_),
    .Y(_075_));
 sky130_fd_sc_hd__inv_1 _151_ (.A(\rd_ptr[2] ),
    .Y(_107_));
 sky130_fd_sc_hd__inv_1 _152_ (.A(\rd_ptr[3] ),
    .Y(_110_));
 sky130_fd_sc_hd__inv_1 _153_ (.A(_085_),
    .Y(_071_));
 sky130_fd_sc_hd__inv_1 _154_ (.A(\wr_ptr[0] ),
    .Y(_003_));
 sky130_fd_sc_hd__inv_1 _155_ (.A(_104_),
    .Y(_113_));
 sky130_fd_sc_hd__xnor2_1 _156_ (.A(\rd_ptr[0] ),
    .B(_032_),
    .Y(_010_));
 sky130_fd_sc_hd__mux2_1 _157_ (.A0(_002_),
    .A1(\rd_ptr[1] ),
    .S(_032_),
    .X(_011_));
 sky130_fd_sc_hd__nand2_1 _158_ (.A(net2),
    .B(_096_),
    .Y(_034_));
 sky130_fd_sc_hd__a21oi_1 _159_ (.A1(_027_),
    .A2(_030_),
    .B1(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__xnor2_1 _160_ (.A(_107_),
    .B(_035_),
    .Y(_012_));
 sky130_fd_sc_hd__nand3_1 _161_ (.A(\rd_ptr[2] ),
    .B(\rd_ptr[1] ),
    .C(\rd_ptr[0] ),
    .Y(_036_));
 sky130_fd_sc_hd__a211oi_1 _162_ (.A1(_027_),
    .A2(_030_),
    .B1(_036_),
    .C1(_031_),
    .Y(_037_));
 sky130_fd_sc_hd__xnor2_1 _163_ (.A(_110_),
    .B(_037_),
    .Y(_013_));
 sky130_fd_sc_hd__a2111oi_1 _164_ (.A1(_027_),
    .A2(_030_),
    .B1(_034_),
    .C1(_110_),
    .D1(_107_),
    .Y(_038_));
 sky130_fd_sc_hd__xor2_1 _165_ (.A(\rd_ptr[4] ),
    .B(_038_),
    .X(_014_));
 sky130_fd_sc_hd__xnor2_1 _166_ (.A(_003_),
    .B(_001_),
    .Y(_015_));
 sky130_fd_sc_hd__mux2_1 _167_ (.A0(\wr_ptr[1] ),
    .A1(_004_),
    .S(_001_),
    .X(_016_));
 sky130_fd_sc_hd__nand2_1 _168_ (.A(net3),
    .B(_095_),
    .Y(_039_));
 sky130_fd_sc_hd__nor3_1 _169_ (.A(_068_),
    .B(_033_),
    .C(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__xor2_1 _170_ (.A(\wr_ptr[2] ),
    .B(_040_),
    .X(_017_));
 sky130_fd_sc_hd__nand4_1 _171_ (.A(net3),
    .B(\wr_ptr[2] ),
    .C(\wr_ptr[1] ),
    .D(\wr_ptr[0] ),
    .Y(_041_));
 sky130_fd_sc_hd__nor3_1 _172_ (.A(_068_),
    .B(_033_),
    .C(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__xor2_1 _173_ (.A(\wr_ptr[3] ),
    .B(_042_),
    .X(_018_));
 sky130_fd_sc_hd__nand2_1 _174_ (.A(\wr_ptr[2] ),
    .B(\wr_ptr[3] ),
    .Y(_043_));
 sky130_fd_sc_hd__nor4_1 _175_ (.A(_068_),
    .B(_033_),
    .C(_039_),
    .D(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__xor2_1 _176_ (.A(\wr_ptr[4] ),
    .B(_044_),
    .X(_019_));
 sky130_fd_sc_hd__clkbuf_2 _177_ (.A(_086_),
    .X(_045_));
 sky130_fd_sc_hd__xnor2_1 _178_ (.A(\pipeline_count[0] ),
    .B(_045_),
    .Y(_005_));
 sky130_fd_sc_hd__mux2i_1 _179_ (.A0(_073_),
    .A1(_078_),
    .S(_045_),
    .Y(_006_));
 sky130_fd_sc_hd__xnor2_1 _180_ (.A(_072_),
    .B(_100_),
    .Y(_046_));
 sky130_fd_sc_hd__nand2_1 _181_ (.A(\pipeline_count[2] ),
    .B(_045_),
    .Y(_047_));
 sky130_fd_sc_hd__o21ai_0 _182_ (.A1(_045_),
    .A2(_046_),
    .B1(_047_),
    .Y(_007_));
 sky130_fd_sc_hd__a21o_1 _183_ (.A1(\pipeline_count[0] ),
    .A2(_098_),
    .B1(_097_),
    .X(_048_));
 sky130_fd_sc_hd__a21oi_1 _184_ (.A1(_100_),
    .A2(_048_),
    .B1(_099_),
    .Y(_049_));
 sky130_fd_sc_hd__xor2_1 _185_ (.A(_102_),
    .B(_049_),
    .X(_050_));
 sky130_fd_sc_hd__nand2_1 _186_ (.A(\pipeline_count[3] ),
    .B(_045_),
    .Y(_051_));
 sky130_fd_sc_hd__o21ai_0 _187_ (.A1(_045_),
    .A2(_050_),
    .B1(_051_),
    .Y(_008_));
 sky130_fd_sc_hd__a21o_1 _188_ (.A1(_072_),
    .A2(_100_),
    .B1(_099_),
    .X(_052_));
 sky130_fd_sc_hd__a21oi_1 _189_ (.A1(_102_),
    .A2(_052_),
    .B1(_101_),
    .Y(_053_));
 sky130_fd_sc_hd__xnor2_1 _190_ (.A(_085_),
    .B(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _191_ (.A(_045_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__xor2_1 _192_ (.A(\pipeline_count[4] ),
    .B(_055_),
    .X(_009_));
 sky130_fd_sc_hd__a21boi_0 _193_ (.A1(_089_),
    .A2(_026_),
    .B1_N(_030_),
    .Y(net4));
 sky130_fd_sc_hd__a21o_1 _194_ (.A1(_092_),
    .A2(_089_),
    .B1(_068_),
    .X(net5));
 sky130_fd_sc_hd__xnor2_1 _195_ (.A(_091_),
    .B(_081_),
    .Y(net8));
 sky130_fd_sc_hd__a21o_1 _196_ (.A1(_088_),
    .A2(_083_),
    .B1(_087_),
    .X(_056_));
 sky130_fd_sc_hd__a21oi_1 _197_ (.A1(_091_),
    .A2(_056_),
    .B1(_090_),
    .Y(_057_));
 sky130_fd_sc_hd__xnor2_1 _198_ (.A(_094_),
    .B(_057_),
    .Y(net9));
 sky130_fd_sc_hd__inv_1 _199_ (.A(_081_),
    .Y(_058_));
 sky130_fd_sc_hd__a21o_1 _200_ (.A1(_091_),
    .A2(_058_),
    .B1(_090_),
    .X(_059_));
 sky130_fd_sc_hd__a21oi_1 _201_ (.A1(_094_),
    .A2(_059_),
    .B1(_093_),
    .Y(_060_));
 sky130_fd_sc_hd__xor2_1 _202_ (.A(\pipeline_count[4] ),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hd__xnor2_1 _203_ (.A(_068_),
    .B(_061_),
    .Y(net10));
 sky130_fd_sc_hd__fa_1 _204_ (.A(\pipeline_count[0] ),
    .B(\pipeline_count[1] ),
    .CIN(_071_),
    .COUT(_072_),
    .SUM(_073_));
 sky130_fd_sc_hd__fa_1 _205_ (.A(_074_),
    .B(\wr_ptr[1] ),
    .CIN(_075_),
    .COUT(_076_),
    .SUM(_077_));
 sky130_fd_sc_hd__fa_1 _206_ (.A(_078_),
    .B(_079_),
    .CIN(_080_),
    .COUT(_081_),
    .SUM(_082_));
 sky130_fd_sc_hd__ha_1 _207_ (.A(_084_),
    .B(\wr_en_pipe[1] ),
    .COUT(_085_),
    .SUM(_086_));
 sky130_fd_sc_hd__ha_1 _208_ (.A(\pipeline_count[1] ),
    .B(_077_),
    .COUT(_087_),
    .SUM(_088_));
 sky130_fd_sc_hd__ha_1 _209_ (.A(\pipeline_count[2] ),
    .B(_089_),
    .COUT(_090_),
    .SUM(_091_));
 sky130_fd_sc_hd__ha_1 _210_ (.A(\pipeline_count[3] ),
    .B(_092_),
    .COUT(_093_),
    .SUM(_094_));
 sky130_fd_sc_hd__ha_1 _211_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .COUT(_095_),
    .SUM(_004_));
 sky130_fd_sc_hd__ha_1 _212_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .COUT(_096_),
    .SUM(_002_));
 sky130_fd_sc_hd__ha_1 _213_ (.A(\pipeline_count[1] ),
    .B(_071_),
    .COUT(_097_),
    .SUM(_098_));
 sky130_fd_sc_hd__ha_1 _214_ (.A(\pipeline_count[2] ),
    .B(_071_),
    .COUT(_099_),
    .SUM(_100_));
 sky130_fd_sc_hd__ha_1 _215_ (.A(\pipeline_count[3] ),
    .B(_071_),
    .COUT(_101_),
    .SUM(_102_));
 sky130_fd_sc_hd__ha_1 _216_ (.A(\rd_ptr[0] ),
    .B(_003_),
    .COUT(_103_),
    .SUM(_104_));
 sky130_fd_sc_hd__ha_1 _217_ (.A(_074_),
    .B(\wr_ptr[1] ),
    .COUT(_105_),
    .SUM(_106_));
 sky130_fd_sc_hd__ha_2 _218_ (.A(_107_),
    .B(\wr_ptr[2] ),
    .COUT(_108_),
    .SUM(_109_));
 sky130_fd_sc_hd__ha_1 _219_ (.A(_110_),
    .B(\wr_ptr[3] ),
    .COUT(_111_),
    .SUM(_112_));
 sky130_fd_sc_hd__ha_1 _220_ (.A(\pipeline_count[0] ),
    .B(_113_),
    .COUT(_083_),
    .SUM(net6));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_4 _222_ (.A(net13),
    .X(rd_data[0]));
 sky130_fd_sc_hd__buf_4 _223_ (.A(net14),
    .X(rd_data[1]));
 sky130_fd_sc_hd__buf_4 _224_ (.A(net15),
    .X(rd_data[2]));
 sky130_fd_sc_hd__buf_4 _225_ (.A(net16),
    .X(rd_data[3]));
 sky130_fd_sc_hd__buf_4 _226_ (.A(net17),
    .X(rd_data[4]));
 sky130_fd_sc_hd__buf_4 _227_ (.A(net18),
    .X(rd_data[5]));
 sky130_fd_sc_hd__buf_4 _228_ (.A(net19),
    .X(rd_data[6]));
 sky130_fd_sc_hd__buf_4 _229_ (.A(net20),
    .X(rd_data[7]));
 sky130_fd_sc_hd__buf_4 _230_ (.A(net21),
    .X(rd_data[8]));
 sky130_fd_sc_hd__buf_4 _231_ (.A(net22),
    .X(rd_data[9]));
 sky130_fd_sc_hd__buf_4 _232_ (.A(net23),
    .X(rd_data[10]));
 sky130_fd_sc_hd__buf_4 _233_ (.A(net24),
    .X(rd_data[11]));
 sky130_fd_sc_hd__buf_4 _234_ (.A(net25),
    .X(rd_data[12]));
 sky130_fd_sc_hd__buf_4 _235_ (.A(net26),
    .X(rd_data[13]));
 sky130_fd_sc_hd__buf_4 _236_ (.A(net27),
    .X(rd_data[14]));
 sky130_fd_sc_hd__buf_4 _237_ (.A(net28),
    .X(rd_data[15]));
 sky130_fd_sc_hd__buf_4 _238_ (.A(net29),
    .X(rd_data[16]));
 sky130_fd_sc_hd__buf_4 _239_ (.A(net30),
    .X(rd_data[17]));
 sky130_fd_sc_hd__buf_4 _240_ (.A(net31),
    .X(rd_data[18]));
 sky130_fd_sc_hd__buf_4 _241_ (.A(net32),
    .X(rd_data[19]));
 sky130_fd_sc_hd__buf_4 _242_ (.A(net33),
    .X(rd_data[20]));
 sky130_fd_sc_hd__buf_4 _243_ (.A(net34),
    .X(rd_data[21]));
 sky130_fd_sc_hd__buf_4 _244_ (.A(net35),
    .X(rd_data[22]));
 sky130_fd_sc_hd__buf_4 _245_ (.A(net36),
    .X(rd_data[23]));
 sky130_fd_sc_hd__buf_4 _246_ (.A(net37),
    .X(rd_data[24]));
 sky130_fd_sc_hd__buf_4 _247_ (.A(net38),
    .X(rd_data[25]));
 sky130_fd_sc_hd__buf_4 _248_ (.A(net39),
    .X(rd_data[26]));
 sky130_fd_sc_hd__buf_4 _249_ (.A(net40),
    .X(rd_data[27]));
 sky130_fd_sc_hd__buf_4 _250_ (.A(net41),
    .X(rd_data[28]));
 sky130_fd_sc_hd__buf_4 _251_ (.A(net42),
    .X(rd_data[29]));
 sky130_fd_sc_hd__buf_4 _252_ (.A(net43),
    .X(rd_data[30]));
 sky130_fd_sc_hd__buf_4 _253_ (.A(net44),
    .X(rd_data[31]));
 sky130_fd_sc_hd__dfrtp_4 \pipeline_count[0]$_DFFE_PN0P_  (.D(_005_),
    .Q(\pipeline_count[0] ),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \pipeline_count[1]$_DFFE_PN0P_  (.D(_006_),
    .Q(\pipeline_count[1] ),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \pipeline_count[2]$_DFFE_PN0P_  (.D(_007_),
    .Q(\pipeline_count[2] ),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \pipeline_count[3]$_DFFE_PN0P_  (.D(_008_),
    .Q(\pipeline_count[3] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \pipeline_count[4]$_DFFE_PN0P_  (.D(_009_),
    .Q(\pipeline_count[4] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_en_pipe$_DFF_PN0_  (.D(_000_),
    .Q(rd_en_pipe),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[0]$_DFFE_PN0P_  (.D(_010_),
    .Q(\rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[1]$_DFFE_PN0P_  (.D(_011_),
    .Q(\rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[2]$_DFFE_PN0P_  (.D(_012_),
    .Q(\rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[3]$_DFFE_PN0P_  (.D(_013_),
    .Q(\rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[4]$_DFFE_PN0P_  (.D(_014_),
    .Q(\rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_en_pipe[0]$_DFF_PN0_  (.D(_001_),
    .Q(\wr_en_pipe[0] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_en_pipe[1]$_DFF_PN0_  (.D(\wr_en_pipe[0] ),
    .Q(\wr_en_pipe[1] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[0]$_DFFE_PN0P_  (.D(_015_),
    .Q(\wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[1]$_DFFE_PN0P_  (.D(_016_),
    .Q(\wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[2]$_DFFE_PN0P_  (.D(_017_),
    .Q(\wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[3]$_DFFE_PN0P_  (.D(_018_),
    .Q(\wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[4]$_DFFE_PN0P_  (.D(_019_),
    .Q(\wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__buf_6 hold1 (.A(net45),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_47 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rd_en),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(wr_en),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 output3 (.A(net4),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output4 (.A(net5),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output5 (.A(net6),
    .X(data_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output6 (.A(net7),
    .X(data_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output7 (.A(net8),
    .X(data_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output8 (.A(net9),
    .X(data_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output9 (.A(net10),
    .X(data_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net11),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net12),
    .X(full));
 sky130_fd_sc_hd__conb_1 _222__12 (.LO(net13));
 sky130_fd_sc_hd__conb_1 _223__13 (.LO(net14));
 sky130_fd_sc_hd__conb_1 _224__14 (.LO(net15));
 sky130_fd_sc_hd__conb_1 _225__15 (.LO(net16));
 sky130_fd_sc_hd__conb_1 _226__16 (.LO(net17));
 sky130_fd_sc_hd__conb_1 _227__17 (.LO(net18));
 sky130_fd_sc_hd__conb_1 _228__18 (.LO(net19));
 sky130_fd_sc_hd__conb_1 _229__19 (.LO(net20));
 sky130_fd_sc_hd__conb_1 _230__20 (.LO(net21));
 sky130_fd_sc_hd__conb_1 _231__21 (.LO(net22));
 sky130_fd_sc_hd__conb_1 _232__22 (.LO(net23));
 sky130_fd_sc_hd__conb_1 _233__23 (.LO(net24));
 sky130_fd_sc_hd__conb_1 _234__24 (.LO(net25));
 sky130_fd_sc_hd__conb_1 _235__25 (.LO(net26));
 sky130_fd_sc_hd__conb_1 _236__26 (.LO(net27));
 sky130_fd_sc_hd__conb_1 _237__27 (.LO(net28));
 sky130_fd_sc_hd__conb_1 _238__28 (.LO(net29));
 sky130_fd_sc_hd__conb_1 _239__29 (.LO(net30));
 sky130_fd_sc_hd__conb_1 _240__30 (.LO(net31));
 sky130_fd_sc_hd__conb_1 _241__31 (.LO(net32));
 sky130_fd_sc_hd__conb_1 _242__32 (.LO(net33));
 sky130_fd_sc_hd__conb_1 _243__33 (.LO(net34));
 sky130_fd_sc_hd__conb_1 _244__34 (.LO(net35));
 sky130_fd_sc_hd__conb_1 _245__35 (.LO(net36));
 sky130_fd_sc_hd__conb_1 _246__36 (.LO(net37));
 sky130_fd_sc_hd__conb_1 _247__37 (.LO(net38));
 sky130_fd_sc_hd__conb_1 _248__38 (.LO(net39));
 sky130_fd_sc_hd__conb_1 _249__39 (.LO(net40));
 sky130_fd_sc_hd__conb_1 _250__40 (.LO(net41));
 sky130_fd_sc_hd__conb_1 _251__41 (.LO(net42));
 sky130_fd_sc_hd__conb_1 _252__42 (.LO(net43));
 sky130_fd_sc_hd__conb_1 _253__43 (.LO(net44));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net45));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_113 ();
endmodule
