module fir_filter (clk,
    data_out_valid,
    data_valid,
    rst_n,
    data_in,
    data_out);
 input clk;
 output data_out_valid;
 input data_valid;
 input rst_n;
 input [7:0] data_in;
 output [18:0] data_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire \delay_line[0][0] ;
 wire \delay_line[0][1] ;
 wire \delay_line[0][2] ;
 wire \delay_line[0][3] ;
 wire \delay_line[0][4] ;
 wire \delay_line[0][5] ;
 wire \delay_line[0][6] ;
 wire \delay_line[0][7] ;
 wire \delay_line[1][0] ;
 wire \delay_line[1][1] ;
 wire \delay_line[1][2] ;
 wire \delay_line[1][3] ;
 wire \delay_line[1][4] ;
 wire \delay_line[1][5] ;
 wire \delay_line[1][6] ;
 wire \delay_line[1][7] ;
 wire \delay_line[2][0] ;
 wire \delay_line[2][1] ;
 wire \delay_line[2][2] ;
 wire \delay_line[2][3] ;
 wire \delay_line[2][4] ;
 wire \delay_line[2][5] ;
 wire \delay_line[2][6] ;
 wire \delay_line[2][7] ;
 wire \delay_line[3][0] ;
 wire \delay_line[3][1] ;
 wire \delay_line[3][2] ;
 wire \delay_line[3][3] ;
 wire \delay_line[3][4] ;
 wire \delay_line[3][5] ;
 wire \delay_line[3][6] ;
 wire \delay_line[3][7] ;
 wire \mac_result[0] ;
 wire \mac_result[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 INV_X1 _325_ (.A(_270_),
    .ZN(_298_));
 INV_X1 _326_ (.A(_303_),
    .ZN(_299_));
 INV_X1 _327_ (.A(_324_),
    .ZN(_300_));
 BUF_X1 _328_ (.A(data_valid),
    .Z(_052_));
 INV_X2 _329_ (.A(_052_),
    .ZN(_053_));
 CLKBUF_X3 _330_ (.A(_053_),
    .Z(_054_));
 CLKBUF_X3 _331_ (.A(_054_),
    .Z(_055_));
 BUF_X2 _332_ (.A(rst_n),
    .Z(_056_));
 INV_X2 _333_ (.A(_056_),
    .ZN(_057_));
 BUF_X4 _334_ (.A(_057_),
    .Z(_058_));
 NOR2_X1 _335_ (.A1(_055_),
    .A2(_058_),
    .ZN(_000_));
 CLKBUF_X3 _336_ (.A(_052_),
    .Z(_059_));
 NAND2_X1 _337_ (.A1(net1),
    .A2(_059_),
    .ZN(_060_));
 NAND2_X1 _338_ (.A1(\delay_line[0][0] ),
    .A2(_054_),
    .ZN(_061_));
 AOI21_X1 _339_ (.A(_058_),
    .B1(_060_),
    .B2(_061_),
    .ZN(_001_));
 CLKBUF_X3 _340_ (.A(_052_),
    .Z(_062_));
 CLKBUF_X3 _341_ (.A(_062_),
    .Z(_063_));
 NAND2_X1 _342_ (.A1(_063_),
    .A2(net2),
    .ZN(_064_));
 CLKBUF_X3 _343_ (.A(_053_),
    .Z(_065_));
 NAND2_X1 _344_ (.A1(_065_),
    .A2(\delay_line[0][1] ),
    .ZN(_066_));
 AOI21_X1 _345_ (.A(_058_),
    .B1(_064_),
    .B2(_066_),
    .ZN(_002_));
 NAND2_X1 _346_ (.A1(_063_),
    .A2(net3),
    .ZN(_067_));
 NAND2_X1 _347_ (.A1(_065_),
    .A2(\delay_line[0][2] ),
    .ZN(_068_));
 AOI21_X1 _348_ (.A(_058_),
    .B1(_067_),
    .B2(_068_),
    .ZN(_003_));
 NAND2_X1 _349_ (.A1(_063_),
    .A2(net4),
    .ZN(_069_));
 NAND2_X1 _350_ (.A1(_065_),
    .A2(\delay_line[0][3] ),
    .ZN(_070_));
 AOI21_X1 _351_ (.A(_058_),
    .B1(_069_),
    .B2(_070_),
    .ZN(_004_));
 NAND2_X1 _352_ (.A1(_063_),
    .A2(net5),
    .ZN(_071_));
 NAND2_X1 _353_ (.A1(_065_),
    .A2(\delay_line[0][4] ),
    .ZN(_072_));
 AOI21_X1 _354_ (.A(_058_),
    .B1(_071_),
    .B2(_072_),
    .ZN(_005_));
 NAND2_X1 _355_ (.A1(_063_),
    .A2(net6),
    .ZN(_073_));
 NAND2_X1 _356_ (.A1(_065_),
    .A2(\delay_line[0][5] ),
    .ZN(_074_));
 AOI21_X1 _357_ (.A(_058_),
    .B1(_073_),
    .B2(_074_),
    .ZN(_006_));
 NAND2_X1 _358_ (.A1(_063_),
    .A2(net7),
    .ZN(_075_));
 NAND2_X1 _359_ (.A1(_065_),
    .A2(\delay_line[0][6] ),
    .ZN(_076_));
 AOI21_X1 _360_ (.A(_058_),
    .B1(_075_),
    .B2(_076_),
    .ZN(_007_));
 NAND2_X1 _361_ (.A1(_063_),
    .A2(net8),
    .ZN(_077_));
 NAND2_X1 _362_ (.A1(_065_),
    .A2(\delay_line[0][7] ),
    .ZN(_078_));
 AOI21_X1 _363_ (.A(_058_),
    .B1(_077_),
    .B2(_078_),
    .ZN(_008_));
 CLKBUF_X3 _364_ (.A(_057_),
    .Z(_079_));
 NAND2_X1 _365_ (.A1(\delay_line[0][0] ),
    .A2(_059_),
    .ZN(_080_));
 NAND2_X1 _366_ (.A1(_065_),
    .A2(\delay_line[1][0] ),
    .ZN(_081_));
 AOI21_X1 _367_ (.A(_079_),
    .B1(_080_),
    .B2(_081_),
    .ZN(_009_));
 NAND2_X1 _368_ (.A1(_063_),
    .A2(\delay_line[0][1] ),
    .ZN(_082_));
 NAND2_X1 _369_ (.A1(_065_),
    .A2(\delay_line[1][1] ),
    .ZN(_083_));
 AOI21_X1 _370_ (.A(_079_),
    .B1(_082_),
    .B2(_083_),
    .ZN(_010_));
 NAND2_X1 _371_ (.A1(_063_),
    .A2(\delay_line[0][2] ),
    .ZN(_084_));
 CLKBUF_X3 _372_ (.A(_053_),
    .Z(_085_));
 NAND2_X1 _373_ (.A1(_085_),
    .A2(\delay_line[1][2] ),
    .ZN(_086_));
 AOI21_X1 _374_ (.A(_079_),
    .B1(_084_),
    .B2(_086_),
    .ZN(_011_));
 NAND2_X1 _375_ (.A1(_063_),
    .A2(\delay_line[0][3] ),
    .ZN(_087_));
 NAND2_X1 _376_ (.A1(_085_),
    .A2(\delay_line[1][3] ),
    .ZN(_088_));
 AOI21_X1 _377_ (.A(_079_),
    .B1(_087_),
    .B2(_088_),
    .ZN(_012_));
 CLKBUF_X3 _378_ (.A(_062_),
    .Z(_089_));
 NAND2_X1 _379_ (.A1(_089_),
    .A2(\delay_line[0][4] ),
    .ZN(_090_));
 NAND2_X1 _380_ (.A1(_085_),
    .A2(\delay_line[1][4] ),
    .ZN(_091_));
 AOI21_X1 _381_ (.A(_079_),
    .B1(_090_),
    .B2(_091_),
    .ZN(_013_));
 NAND2_X1 _382_ (.A1(_089_),
    .A2(\delay_line[0][5] ),
    .ZN(_092_));
 NAND2_X1 _383_ (.A1(_085_),
    .A2(\delay_line[1][5] ),
    .ZN(_093_));
 AOI21_X1 _384_ (.A(_079_),
    .B1(_092_),
    .B2(_093_),
    .ZN(_014_));
 NAND2_X1 _385_ (.A1(_089_),
    .A2(\delay_line[0][6] ),
    .ZN(_094_));
 NAND2_X1 _386_ (.A1(_085_),
    .A2(\delay_line[1][6] ),
    .ZN(_095_));
 AOI21_X1 _387_ (.A(_079_),
    .B1(_094_),
    .B2(_095_),
    .ZN(_015_));
 NAND2_X1 _388_ (.A1(_089_),
    .A2(\delay_line[0][7] ),
    .ZN(_096_));
 NAND2_X1 _389_ (.A1(_085_),
    .A2(\delay_line[1][7] ),
    .ZN(_097_));
 AOI21_X1 _390_ (.A(_079_),
    .B1(_096_),
    .B2(_097_),
    .ZN(_016_));
 NAND2_X1 _391_ (.A1(_089_),
    .A2(\delay_line[1][0] ),
    .ZN(_098_));
 NAND2_X1 _392_ (.A1(_085_),
    .A2(\delay_line[2][0] ),
    .ZN(_099_));
 AOI21_X1 _393_ (.A(_079_),
    .B1(_098_),
    .B2(_099_),
    .ZN(_017_));
 NAND2_X1 _394_ (.A1(_089_),
    .A2(\delay_line[1][1] ),
    .ZN(_100_));
 NAND2_X1 _395_ (.A1(_085_),
    .A2(\delay_line[2][1] ),
    .ZN(_101_));
 AOI21_X1 _396_ (.A(_079_),
    .B1(_100_),
    .B2(_101_),
    .ZN(_018_));
 CLKBUF_X3 _397_ (.A(_057_),
    .Z(_102_));
 NAND2_X1 _398_ (.A1(_089_),
    .A2(\delay_line[1][2] ),
    .ZN(_103_));
 NAND2_X1 _399_ (.A1(_085_),
    .A2(\delay_line[2][2] ),
    .ZN(_104_));
 AOI21_X1 _400_ (.A(_102_),
    .B1(_103_),
    .B2(_104_),
    .ZN(_019_));
 NAND2_X1 _401_ (.A1(_089_),
    .A2(\delay_line[1][3] ),
    .ZN(_105_));
 NAND2_X1 _402_ (.A1(_085_),
    .A2(\delay_line[2][3] ),
    .ZN(_106_));
 AOI21_X1 _403_ (.A(_102_),
    .B1(_105_),
    .B2(_106_),
    .ZN(_020_));
 NAND2_X1 _404_ (.A1(_089_),
    .A2(\delay_line[1][4] ),
    .ZN(_107_));
 CLKBUF_X3 _405_ (.A(_053_),
    .Z(_108_));
 NAND2_X1 _406_ (.A1(_108_),
    .A2(\delay_line[2][4] ),
    .ZN(_109_));
 AOI21_X1 _407_ (.A(_102_),
    .B1(_107_),
    .B2(_109_),
    .ZN(_021_));
 NAND2_X1 _408_ (.A1(_089_),
    .A2(\delay_line[1][5] ),
    .ZN(_110_));
 NAND2_X1 _409_ (.A1(_108_),
    .A2(\delay_line[2][5] ),
    .ZN(_111_));
 AOI21_X1 _410_ (.A(_102_),
    .B1(_110_),
    .B2(_111_),
    .ZN(_022_));
 CLKBUF_X3 _411_ (.A(_062_),
    .Z(_112_));
 NAND2_X1 _412_ (.A1(_112_),
    .A2(\delay_line[1][6] ),
    .ZN(_113_));
 NAND2_X1 _413_ (.A1(_108_),
    .A2(\delay_line[2][6] ),
    .ZN(_114_));
 AOI21_X1 _414_ (.A(_102_),
    .B1(_113_),
    .B2(_114_),
    .ZN(_023_));
 NAND2_X1 _415_ (.A1(_112_),
    .A2(\delay_line[1][7] ),
    .ZN(_115_));
 NAND2_X1 _416_ (.A1(_108_),
    .A2(\delay_line[2][7] ),
    .ZN(_116_));
 AOI21_X1 _417_ (.A(_102_),
    .B1(_115_),
    .B2(_116_),
    .ZN(_024_));
 NAND2_X1 _418_ (.A1(_112_),
    .A2(\delay_line[2][0] ),
    .ZN(_117_));
 NAND2_X1 _419_ (.A1(_108_),
    .A2(\delay_line[3][0] ),
    .ZN(_118_));
 AOI21_X1 _420_ (.A(_102_),
    .B1(_117_),
    .B2(_118_),
    .ZN(_025_));
 NAND2_X1 _421_ (.A1(_112_),
    .A2(\delay_line[2][1] ),
    .ZN(_119_));
 NAND2_X1 _422_ (.A1(_108_),
    .A2(\delay_line[3][1] ),
    .ZN(_120_));
 AOI21_X1 _423_ (.A(_102_),
    .B1(_119_),
    .B2(_120_),
    .ZN(_026_));
 NAND2_X1 _424_ (.A1(_112_),
    .A2(\delay_line[2][2] ),
    .ZN(_121_));
 NAND2_X1 _425_ (.A1(_108_),
    .A2(\delay_line[3][2] ),
    .ZN(_122_));
 AOI21_X1 _426_ (.A(_102_),
    .B1(_121_),
    .B2(_122_),
    .ZN(_027_));
 NAND2_X1 _427_ (.A1(_112_),
    .A2(\delay_line[2][3] ),
    .ZN(_123_));
 NAND2_X1 _428_ (.A1(_108_),
    .A2(\delay_line[3][3] ),
    .ZN(_124_));
 AOI21_X1 _429_ (.A(_102_),
    .B1(_123_),
    .B2(_124_),
    .ZN(_028_));
 CLKBUF_X3 _430_ (.A(_057_),
    .Z(_125_));
 NAND2_X1 _431_ (.A1(_112_),
    .A2(\delay_line[2][4] ),
    .ZN(_126_));
 NAND2_X1 _432_ (.A1(_108_),
    .A2(\delay_line[3][4] ),
    .ZN(_127_));
 AOI21_X1 _433_ (.A(_125_),
    .B1(_126_),
    .B2(_127_),
    .ZN(_029_));
 NAND2_X1 _434_ (.A1(_112_),
    .A2(\delay_line[2][5] ),
    .ZN(_128_));
 NAND2_X1 _435_ (.A1(_108_),
    .A2(\delay_line[3][5] ),
    .ZN(_129_));
 AOI21_X1 _436_ (.A(_125_),
    .B1(_128_),
    .B2(_129_),
    .ZN(_030_));
 NAND2_X1 _437_ (.A1(_112_),
    .A2(\delay_line[2][6] ),
    .ZN(_130_));
 NAND2_X1 _438_ (.A1(_054_),
    .A2(\delay_line[3][6] ),
    .ZN(_131_));
 AOI21_X1 _439_ (.A(_125_),
    .B1(_130_),
    .B2(_131_),
    .ZN(_031_));
 NAND2_X1 _440_ (.A1(_112_),
    .A2(\delay_line[2][7] ),
    .ZN(_132_));
 NAND2_X1 _441_ (.A1(_054_),
    .A2(\delay_line[3][7] ),
    .ZN(_133_));
 AOI21_X1 _442_ (.A(_125_),
    .B1(_132_),
    .B2(_133_),
    .ZN(_032_));
 NAND2_X1 _443_ (.A1(_059_),
    .A2(\mac_result[0] ),
    .ZN(_134_));
 NAND2_X1 _444_ (.A1(_054_),
    .A2(net9),
    .ZN(_135_));
 AOI21_X1 _445_ (.A(_125_),
    .B1(_134_),
    .B2(_135_),
    .ZN(_033_));
 NAND2_X1 _446_ (.A1(_055_),
    .A2(net10),
    .ZN(_136_));
 INV_X1 _447_ (.A(_311_),
    .ZN(_137_));
 AOI21_X2 _448_ (.A(_304_),
    .B1(_324_),
    .B2(_305_),
    .ZN(_138_));
 BUF_X2 _449_ (.A(_308_),
    .Z(_139_));
 BUF_X2 _450_ (.A(_310_),
    .Z(_140_));
 NAND3_X1 _451_ (.A1(_139_),
    .A2(_140_),
    .A3(_312_),
    .ZN(_141_));
 AOI21_X1 _452_ (.A(_309_),
    .B1(_307_),
    .B2(_140_),
    .ZN(_142_));
 INV_X1 _453_ (.A(_312_),
    .ZN(_143_));
 OAI221_X2 _454_ (.A(_137_),
    .B1(_138_),
    .B2(_141_),
    .C1(_142_),
    .C2(_143_),
    .ZN(_144_));
 BUF_X4 _455_ (.A(_314_),
    .Z(_145_));
 BUF_X1 _456_ (.A(_318_),
    .Z(_146_));
 BUF_X1 _457_ (.A(_320_),
    .Z(_147_));
 BUF_X4 _458_ (.A(_316_),
    .Z(_148_));
 OR2_X1 _459_ (.A1(_148_),
    .A2(_315_),
    .ZN(_149_));
 AND4_X1 _460_ (.A1(_145_),
    .A2(_146_),
    .A3(_147_),
    .A4(_149_),
    .ZN(_150_));
 INV_X1 _461_ (.A(_317_),
    .ZN(_151_));
 AOI21_X1 _462_ (.A(_315_),
    .B1(_313_),
    .B2(_148_),
    .ZN(_152_));
 INV_X1 _463_ (.A(_146_),
    .ZN(_153_));
 OAI21_X1 _464_ (.A(_151_),
    .B1(_152_),
    .B2(_153_),
    .ZN(_154_));
 AOI221_X2 _465_ (.A(_319_),
    .B1(_144_),
    .B2(_150_),
    .C1(_154_),
    .C2(_147_),
    .ZN(_155_));
 XNOR2_X1 _466_ (.A(_322_),
    .B(_155_),
    .ZN(_156_));
 NAND2_X1 _467_ (.A1(_059_),
    .A2(_156_),
    .ZN(_157_));
 AOI21_X1 _468_ (.A(_125_),
    .B1(_136_),
    .B2(_157_),
    .ZN(_034_));
 INV_X1 _469_ (.A(_322_),
    .ZN(_158_));
 AOI21_X4 _470_ (.A(_053_),
    .B1(_321_),
    .B2(_158_),
    .ZN(_159_));
 OR3_X1 _471_ (.A1(_158_),
    .A2(_319_),
    .A3(_321_),
    .ZN(_160_));
 AOI21_X1 _472_ (.A(_057_),
    .B1(_159_),
    .B2(_160_),
    .ZN(_161_));
 NAND2_X1 _473_ (.A1(_147_),
    .A2(_159_),
    .ZN(_162_));
 AOI21_X1 _474_ (.A(_313_),
    .B1(_311_),
    .B2(_145_),
    .ZN(_163_));
 INV_X1 _475_ (.A(_301_),
    .ZN(_164_));
 AOI21_X2 _476_ (.A(_307_),
    .B1(_164_),
    .B2(_139_),
    .ZN(_165_));
 NAND3_X1 _477_ (.A1(_140_),
    .A2(_312_),
    .A3(_145_),
    .ZN(_166_));
 NAND2_X1 _478_ (.A1(_312_),
    .A2(_145_),
    .ZN(_167_));
 INV_X1 _479_ (.A(_309_),
    .ZN(_168_));
 OAI221_X2 _480_ (.A(_163_),
    .B1(_165_),
    .B2(_166_),
    .C1(_167_),
    .C2(_168_),
    .ZN(_169_));
 AND2_X1 _481_ (.A1(_148_),
    .A2(_146_),
    .ZN(_170_));
 AOI221_X2 _482_ (.A(_317_),
    .B1(_169_),
    .B2(_170_),
    .C1(_315_),
    .C2(_146_),
    .ZN(_171_));
 OAI21_X2 _483_ (.A(_161_),
    .B1(_162_),
    .B2(_171_),
    .ZN(_172_));
 INV_X1 _484_ (.A(net11),
    .ZN(_173_));
 AOI21_X1 _485_ (.A(_172_),
    .B1(_173_),
    .B2(_055_),
    .ZN(_035_));
 OAI21_X1 _486_ (.A(_056_),
    .B1(net12),
    .B2(_062_),
    .ZN(_174_));
 INV_X1 _487_ (.A(_321_),
    .ZN(_175_));
 NAND3_X2 _488_ (.A1(_322_),
    .A2(_175_),
    .A3(_155_),
    .ZN(_176_));
 AOI21_X1 _489_ (.A(_174_),
    .B1(_176_),
    .B2(_159_),
    .ZN(_036_));
 INV_X1 _490_ (.A(net13),
    .ZN(_177_));
 AOI21_X1 _491_ (.A(_172_),
    .B1(_177_),
    .B2(_055_),
    .ZN(_037_));
 OAI21_X1 _492_ (.A(_056_),
    .B1(net14),
    .B2(_062_),
    .ZN(_178_));
 AOI21_X1 _493_ (.A(_178_),
    .B1(_176_),
    .B2(_159_),
    .ZN(_038_));
 INV_X1 _494_ (.A(net15),
    .ZN(_179_));
 AOI21_X1 _495_ (.A(_172_),
    .B1(_179_),
    .B2(_055_),
    .ZN(_039_));
 OAI21_X1 _496_ (.A(_056_),
    .B1(net16),
    .B2(_062_),
    .ZN(_180_));
 AOI21_X1 _497_ (.A(_180_),
    .B1(_176_),
    .B2(_159_),
    .ZN(_040_));
 INV_X1 _498_ (.A(net17),
    .ZN(_181_));
 AOI21_X1 _499_ (.A(_172_),
    .B1(_181_),
    .B2(_055_),
    .ZN(_041_));
 OAI21_X1 _500_ (.A(_056_),
    .B1(net18),
    .B2(_062_),
    .ZN(_182_));
 AOI21_X1 _501_ (.A(_182_),
    .B1(_176_),
    .B2(_159_),
    .ZN(_042_));
 NAND2_X1 _502_ (.A1(_059_),
    .A2(\mac_result[1] ),
    .ZN(_183_));
 NAND2_X1 _503_ (.A1(_054_),
    .A2(net19),
    .ZN(_184_));
 AOI21_X1 _504_ (.A(_125_),
    .B1(_183_),
    .B2(_184_),
    .ZN(_043_));
 NOR2_X1 _505_ (.A1(_302_),
    .A2(_054_),
    .ZN(_185_));
 AOI21_X1 _506_ (.A(_185_),
    .B1(net20),
    .B2(_054_),
    .ZN(_186_));
 NOR2_X1 _507_ (.A1(_058_),
    .A2(_186_),
    .ZN(_044_));
 NAND2_X1 _508_ (.A1(_055_),
    .A2(net21),
    .ZN(_187_));
 XNOR2_X1 _509_ (.A(_139_),
    .B(_301_),
    .ZN(_188_));
 NAND2_X1 _510_ (.A1(_059_),
    .A2(_188_),
    .ZN(_189_));
 AOI21_X1 _511_ (.A(_125_),
    .B1(_187_),
    .B2(_189_),
    .ZN(_045_));
 NAND2_X1 _512_ (.A1(_055_),
    .A2(net22),
    .ZN(_190_));
 INV_X1 _513_ (.A(_138_),
    .ZN(_191_));
 AOI21_X1 _514_ (.A(_307_),
    .B1(_191_),
    .B2(_139_),
    .ZN(_192_));
 XNOR2_X1 _515_ (.A(_140_),
    .B(_192_),
    .ZN(_193_));
 NAND2_X1 _516_ (.A1(_059_),
    .A2(_193_),
    .ZN(_194_));
 AOI21_X1 _517_ (.A(_125_),
    .B1(_190_),
    .B2(_194_),
    .ZN(_046_));
 NAND2_X1 _518_ (.A1(_055_),
    .A2(net23),
    .ZN(_195_));
 INV_X1 _519_ (.A(_140_),
    .ZN(_196_));
 OAI21_X1 _520_ (.A(_168_),
    .B1(_165_),
    .B2(_196_),
    .ZN(_197_));
 XNOR2_X1 _521_ (.A(_143_),
    .B(_197_),
    .ZN(_198_));
 NAND2_X1 _522_ (.A1(_059_),
    .A2(_198_),
    .ZN(_199_));
 AOI21_X1 _523_ (.A(_125_),
    .B1(_195_),
    .B2(_199_),
    .ZN(_047_));
 NAND2_X1 _524_ (.A1(_055_),
    .A2(net24),
    .ZN(_200_));
 XOR2_X1 _525_ (.A(_145_),
    .B(_144_),
    .Z(_201_));
 NAND2_X1 _526_ (.A1(_059_),
    .A2(_201_),
    .ZN(_202_));
 AOI21_X1 _527_ (.A(_057_),
    .B1(_200_),
    .B2(_202_),
    .ZN(_048_));
 NAND2_X1 _528_ (.A1(_065_),
    .A2(net25),
    .ZN(_203_));
 XOR2_X1 _529_ (.A(_148_),
    .B(_169_),
    .Z(_204_));
 NAND2_X1 _530_ (.A1(_059_),
    .A2(_204_),
    .ZN(_205_));
 AOI21_X1 _531_ (.A(_057_),
    .B1(_203_),
    .B2(_205_),
    .ZN(_049_));
 NAND3_X1 _532_ (.A1(_145_),
    .A2(_148_),
    .A3(_144_),
    .ZN(_206_));
 NAND2_X1 _533_ (.A1(_152_),
    .A2(_206_),
    .ZN(_207_));
 NAND4_X1 _534_ (.A1(_153_),
    .A2(_062_),
    .A3(_056_),
    .A4(_207_),
    .ZN(_208_));
 NAND3_X1 _535_ (.A1(_146_),
    .A2(_062_),
    .A3(_056_),
    .ZN(_209_));
 NAND2_X1 _536_ (.A1(_054_),
    .A2(net26),
    .ZN(_210_));
 OAI221_X1 _537_ (.A(_208_),
    .B1(_209_),
    .B2(_207_),
    .C1(_210_),
    .C2(_057_),
    .ZN(_050_));
 NAND4_X1 _538_ (.A1(_147_),
    .A2(_062_),
    .A3(_056_),
    .A4(_171_),
    .ZN(_211_));
 OR3_X1 _539_ (.A1(_147_),
    .A2(_053_),
    .A3(_057_),
    .ZN(_212_));
 NAND2_X1 _540_ (.A1(_054_),
    .A2(net27),
    .ZN(_213_));
 OAI221_X1 _541_ (.A(_211_),
    .B1(_212_),
    .B2(_171_),
    .C1(_057_),
    .C2(_213_),
    .ZN(_051_));
 FA_X1 _542_ (.A(\delay_line[0][2] ),
    .B(\delay_line[1][1] ),
    .CI(\delay_line[2][1] ),
    .CO(_266_),
    .S(_267_));
 FA_X1 _543_ (.A(\delay_line[3][2] ),
    .B(_267_),
    .CI(_268_),
    .CO(_269_),
    .S(_270_));
 FA_X1 _544_ (.A(\delay_line[0][1] ),
    .B(\delay_line[1][0] ),
    .CI(\delay_line[2][0] ),
    .CO(_268_),
    .S(_271_));
 FA_X1 _545_ (.A(\delay_line[0][3] ),
    .B(\delay_line[1][2] ),
    .CI(\delay_line[2][2] ),
    .CO(_272_),
    .S(_273_));
 FA_X1 _546_ (.A(\delay_line[3][3] ),
    .B(_273_),
    .CI(_266_),
    .CO(_274_),
    .S(_275_));
 FA_X1 _547_ (.A(\delay_line[0][4] ),
    .B(\delay_line[1][3] ),
    .CI(\delay_line[2][3] ),
    .CO(_276_),
    .S(_277_));
 FA_X1 _548_ (.A(\delay_line[3][4] ),
    .B(_277_),
    .CI(_272_),
    .CO(_278_),
    .S(_279_));
 FA_X1 _549_ (.A(\delay_line[0][5] ),
    .B(\delay_line[1][4] ),
    .CI(\delay_line[2][4] ),
    .CO(_280_),
    .S(_281_));
 FA_X1 _550_ (.A(\delay_line[3][5] ),
    .B(_281_),
    .CI(_276_),
    .CO(_282_),
    .S(_283_));
 FA_X1 _551_ (.A(\delay_line[0][6] ),
    .B(\delay_line[1][5] ),
    .CI(\delay_line[2][5] ),
    .CO(_284_),
    .S(_285_));
 FA_X1 _552_ (.A(\delay_line[3][6] ),
    .B(_285_),
    .CI(_280_),
    .CO(_286_),
    .S(_287_));
 FA_X1 _553_ (.A(\delay_line[0][7] ),
    .B(\delay_line[1][6] ),
    .CI(\delay_line[2][6] ),
    .CO(_288_),
    .S(_289_));
 FA_X1 _554_ (.A(\delay_line[3][7] ),
    .B(_289_),
    .CI(_284_),
    .CO(_290_),
    .S(_291_));
 FA_X1 _555_ (.A(\delay_line[0][7] ),
    .B(\delay_line[1][7] ),
    .CI(\delay_line[2][7] ),
    .CO(_292_),
    .S(_293_));
 FA_X1 _556_ (.A(\delay_line[3][7] ),
    .B(_293_),
    .CI(_288_),
    .CO(_294_),
    .S(_295_));
 FA_X1 _557_ (.A(\delay_line[3][7] ),
    .B(_293_),
    .CI(_292_),
    .CO(_296_),
    .S(_297_));
 FA_X1 _558_ (.A(_298_),
    .B(_299_),
    .CI(_300_),
    .CO(_301_),
    .S(_302_));
 HA_X1 _559_ (.A(_270_),
    .B(_303_),
    .CO(_304_),
    .S(_305_));
 HA_X1 _560_ (.A(\delay_line[3][1] ),
    .B(_271_),
    .CO(_303_),
    .S(_306_));
 HA_X1 _561_ (.A(_275_),
    .B(_269_),
    .CO(_307_),
    .S(_308_));
 HA_X1 _562_ (.A(_279_),
    .B(_274_),
    .CO(_309_),
    .S(_310_));
 HA_X1 _563_ (.A(_283_),
    .B(_278_),
    .CO(_311_),
    .S(_312_));
 HA_X1 _564_ (.A(_287_),
    .B(_282_),
    .CO(_313_),
    .S(_314_));
 HA_X1 _565_ (.A(_291_),
    .B(_286_),
    .CO(_315_),
    .S(_316_));
 HA_X1 _566_ (.A(_295_),
    .B(_290_),
    .CO(_317_),
    .S(_318_));
 HA_X1 _567_ (.A(_297_),
    .B(_294_),
    .CO(_319_),
    .S(_320_));
 HA_X1 _568_ (.A(_297_),
    .B(_296_),
    .CO(_321_),
    .S(_322_));
 HA_X1 _569_ (.A(\delay_line[0][0] ),
    .B(\delay_line[3][0] ),
    .CO(_323_),
    .S(\mac_result[0] ));
 HA_X1 _570_ (.A(_306_),
    .B(_323_),
    .CO(_324_),
    .S(\mac_result[1] ));
 DFF_X1 \data_out_valid$_SDFF_PN0_  (.D(_000_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net28),
    .QN(_265_));
 DFF_X1 \delay_line[0][0]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[0][0] ),
    .QN(_264_));
 DFF_X2 \delay_line[0][1]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[0][1] ),
    .QN(_263_));
 DFF_X1 \delay_line[0][2]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[0][2] ),
    .QN(_262_));
 DFF_X2 \delay_line[0][3]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[0][3] ),
    .QN(_261_));
 DFF_X1 \delay_line[0][4]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[0][4] ),
    .QN(_260_));
 DFF_X2 \delay_line[0][5]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[0][5] ),
    .QN(_259_));
 DFF_X1 \delay_line[0][6]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[0][6] ),
    .QN(_258_));
 DFF_X2 \delay_line[0][7]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[0][7] ),
    .QN(_257_));
 DFF_X1 \delay_line[1][0]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[1][0] ),
    .QN(_256_));
 DFF_X1 \delay_line[1][1]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[1][1] ),
    .QN(_255_));
 DFF_X1 \delay_line[1][2]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[1][2] ),
    .QN(_254_));
 DFF_X1 \delay_line[1][3]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[1][3] ),
    .QN(_253_));
 DFF_X1 \delay_line[1][4]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[1][4] ),
    .QN(_252_));
 DFF_X1 \delay_line[1][5]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[1][5] ),
    .QN(_251_));
 DFF_X1 \delay_line[1][6]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[1][6] ),
    .QN(_250_));
 DFF_X1 \delay_line[1][7]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[1][7] ),
    .QN(_249_));
 DFF_X1 \delay_line[2][0]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[2][0] ),
    .QN(_248_));
 DFF_X1 \delay_line[2][1]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[2][1] ),
    .QN(_247_));
 DFF_X1 \delay_line[2][2]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[2][2] ),
    .QN(_246_));
 DFF_X1 \delay_line[2][3]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[2][3] ),
    .QN(_245_));
 DFF_X1 \delay_line[2][4]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[2][4] ),
    .QN(_244_));
 DFF_X1 \delay_line[2][5]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[2][5] ),
    .QN(_243_));
 DFF_X1 \delay_line[2][6]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[2][6] ),
    .QN(_242_));
 DFF_X1 \delay_line[2][7]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[2][7] ),
    .QN(_241_));
 DFF_X1 \delay_line[3][0]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[3][0] ),
    .QN(_240_));
 DFF_X1 \delay_line[3][1]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\delay_line[3][1] ),
    .QN(_239_));
 DFF_X1 \delay_line[3][2]$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\delay_line[3][2] ),
    .QN(_238_));
 DFF_X1 \delay_line[3][3]$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\delay_line[3][3] ),
    .QN(_237_));
 DFF_X1 \delay_line[3][4]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\delay_line[3][4] ),
    .QN(_236_));
 DFF_X1 \delay_line[3][5]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\delay_line[3][5] ),
    .QN(_235_));
 DFF_X1 \delay_line[3][6]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\delay_line[3][6] ),
    .QN(_234_));
 DFF_X2 \delay_line[3][7]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\delay_line[3][7] ),
    .QN(_233_));
 DFF_X1 \result[0]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net9),
    .QN(_232_));
 DFF_X1 \result[10]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net10),
    .QN(_231_));
 DFF_X1 \result[11]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net11),
    .QN(_230_));
 DFF_X1 \result[12]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net12),
    .QN(_229_));
 DFF_X1 \result[13]$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net13),
    .QN(_228_));
 DFF_X1 \result[14]$_SDFFE_PN0P_  (.D(_038_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net14),
    .QN(_227_));
 DFF_X1 \result[15]$_SDFFE_PN0P_  (.D(_039_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net15),
    .QN(_226_));
 DFF_X1 \result[16]$_SDFFE_PN0P_  (.D(_040_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net16),
    .QN(_225_));
 DFF_X1 \result[17]$_SDFFE_PN0P_  (.D(_041_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net17),
    .QN(_224_));
 DFF_X1 \result[18]$_SDFFE_PN0P_  (.D(_042_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net18),
    .QN(_223_));
 DFF_X1 \result[1]$_SDFFE_PN0P_  (.D(_043_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net19),
    .QN(_222_));
 DFF_X1 \result[2]$_SDFFE_PN0P_  (.D(_044_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net20),
    .QN(_221_));
 DFF_X1 \result[3]$_SDFFE_PN0P_  (.D(_045_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net21),
    .QN(_220_));
 DFF_X1 \result[4]$_SDFFE_PN0P_  (.D(_046_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net22),
    .QN(_219_));
 DFF_X1 \result[5]$_SDFFE_PN0P_  (.D(_047_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net23),
    .QN(_218_));
 DFF_X1 \result[6]$_SDFFE_PN0P_  (.D(_048_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net24),
    .QN(_217_));
 DFF_X1 \result[7]$_SDFFE_PN0P_  (.D(_049_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net25),
    .QN(_216_));
 DFF_X1 \result[8]$_SDFFE_PN0P_  (.D(_050_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net26),
    .QN(_215_));
 DFF_X1 \result[9]$_SDFFE_PN0P_  (.D(_051_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net27),
    .QN(_214_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_111 ();
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[2]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[3]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[5]),
    .Z(net6));
 BUF_X1 input7 (.A(data_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[7]),
    .Z(net8));
 BUF_X1 output9 (.A(net9),
    .Z(data_out[0]));
 BUF_X1 output10 (.A(net10),
    .Z(data_out[10]));
 BUF_X1 output11 (.A(net11),
    .Z(data_out[11]));
 BUF_X1 output12 (.A(net12),
    .Z(data_out[12]));
 BUF_X1 output13 (.A(net13),
    .Z(data_out[13]));
 BUF_X1 output14 (.A(net14),
    .Z(data_out[14]));
 BUF_X1 output15 (.A(net15),
    .Z(data_out[15]));
 BUF_X1 output16 (.A(net16),
    .Z(data_out[16]));
 BUF_X1 output17 (.A(net17),
    .Z(data_out[17]));
 BUF_X1 output18 (.A(net18),
    .Z(data_out[18]));
 BUF_X1 output19 (.A(net19),
    .Z(data_out[1]));
 BUF_X1 output20 (.A(net20),
    .Z(data_out[2]));
 BUF_X1 output21 (.A(net21),
    .Z(data_out[3]));
 BUF_X1 output22 (.A(net22),
    .Z(data_out[4]));
 BUF_X1 output23 (.A(net23),
    .Z(data_out[5]));
 BUF_X1 output24 (.A(net24),
    .Z(data_out[6]));
 BUF_X1 output25 (.A(net25),
    .Z(data_out[7]));
 BUF_X1 output26 (.A(net26),
    .Z(data_out[8]));
 BUF_X1 output27 (.A(net27),
    .Z(data_out[9]));
 BUF_X1 output28 (.A(net28),
    .Z(data_out_valid));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_2_1__leaf_clk));
 INV_X2 clkload2 (.A(clknet_2_3__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X16 FILLER_0_129 ();
 FILLCELL_X8 FILLER_0_145 ();
 FILLCELL_X1 FILLER_0_153 ();
 FILLCELL_X32 FILLER_0_160 ();
 FILLCELL_X8 FILLER_0_192 ();
 FILLCELL_X4 FILLER_0_200 ();
 FILLCELL_X32 FILLER_0_207 ();
 FILLCELL_X4 FILLER_0_239 ();
 FILLCELL_X2 FILLER_0_243 ();
 FILLCELL_X32 FILLER_0_248 ();
 FILLCELL_X32 FILLER_0_280 ();
 FILLCELL_X32 FILLER_0_312 ();
 FILLCELL_X32 FILLER_0_344 ();
 FILLCELL_X32 FILLER_0_376 ();
 FILLCELL_X8 FILLER_0_408 ();
 FILLCELL_X2 FILLER_0_416 ();
 FILLCELL_X1 FILLER_0_418 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X8 FILLER_1_161 ();
 FILLCELL_X2 FILLER_1_169 ();
 FILLCELL_X32 FILLER_1_174 ();
 FILLCELL_X32 FILLER_1_206 ();
 FILLCELL_X32 FILLER_1_238 ();
 FILLCELL_X8 FILLER_1_270 ();
 FILLCELL_X2 FILLER_1_278 ();
 FILLCELL_X1 FILLER_1_280 ();
 FILLCELL_X4 FILLER_1_284 ();
 FILLCELL_X2 FILLER_1_288 ();
 FILLCELL_X1 FILLER_1_290 ();
 FILLCELL_X32 FILLER_1_294 ();
 FILLCELL_X32 FILLER_1_326 ();
 FILLCELL_X32 FILLER_1_358 ();
 FILLCELL_X16 FILLER_1_390 ();
 FILLCELL_X8 FILLER_1_406 ();
 FILLCELL_X4 FILLER_1_414 ();
 FILLCELL_X1 FILLER_1_418 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X2 FILLER_2_417 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X2 FILLER_3_417 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X2 FILLER_4_417 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X2 FILLER_5_417 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X2 FILLER_6_417 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X2 FILLER_7_417 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X2 FILLER_8_417 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X2 FILLER_9_417 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X2 FILLER_10_417 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X2 FILLER_11_417 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X2 FILLER_12_417 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X2 FILLER_13_417 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X2 FILLER_14_417 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X2 FILLER_15_417 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X2 FILLER_16_417 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X2 FILLER_17_417 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X2 FILLER_18_417 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X16 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_212 ();
 FILLCELL_X2 FILLER_19_244 ();
 FILLCELL_X1 FILLER_19_246 ();
 FILLCELL_X32 FILLER_19_250 ();
 FILLCELL_X4 FILLER_19_285 ();
 FILLCELL_X2 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_294 ();
 FILLCELL_X32 FILLER_19_326 ();
 FILLCELL_X32 FILLER_19_358 ();
 FILLCELL_X16 FILLER_19_390 ();
 FILLCELL_X8 FILLER_19_406 ();
 FILLCELL_X4 FILLER_19_414 ();
 FILLCELL_X1 FILLER_19_418 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X16 FILLER_20_129 ();
 FILLCELL_X8 FILLER_20_145 ();
 FILLCELL_X4 FILLER_20_153 ();
 FILLCELL_X2 FILLER_20_157 ();
 FILLCELL_X1 FILLER_20_159 ();
 FILLCELL_X8 FILLER_20_163 ();
 FILLCELL_X2 FILLER_20_171 ();
 FILLCELL_X32 FILLER_20_176 ();
 FILLCELL_X32 FILLER_20_208 ();
 FILLCELL_X4 FILLER_20_240 ();
 FILLCELL_X16 FILLER_20_248 ();
 FILLCELL_X8 FILLER_20_264 ();
 FILLCELL_X4 FILLER_20_272 ();
 FILLCELL_X2 FILLER_20_276 ();
 FILLCELL_X1 FILLER_20_278 ();
 FILLCELL_X8 FILLER_20_283 ();
 FILLCELL_X32 FILLER_20_295 ();
 FILLCELL_X32 FILLER_20_327 ();
 FILLCELL_X32 FILLER_20_359 ();
 FILLCELL_X16 FILLER_20_391 ();
 FILLCELL_X8 FILLER_20_407 ();
 FILLCELL_X4 FILLER_20_415 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X2 FILLER_21_168 ();
 FILLCELL_X1 FILLER_21_170 ();
 FILLCELL_X8 FILLER_21_197 ();
 FILLCELL_X4 FILLER_21_205 ();
 FILLCELL_X2 FILLER_21_209 ();
 FILLCELL_X16 FILLER_21_218 ();
 FILLCELL_X4 FILLER_21_234 ();
 FILLCELL_X8 FILLER_21_257 ();
 FILLCELL_X4 FILLER_21_265 ();
 FILLCELL_X32 FILLER_21_305 ();
 FILLCELL_X32 FILLER_21_337 ();
 FILLCELL_X32 FILLER_21_369 ();
 FILLCELL_X16 FILLER_21_401 ();
 FILLCELL_X2 FILLER_21_417 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X16 FILLER_22_129 ();
 FILLCELL_X8 FILLER_22_145 ();
 FILLCELL_X4 FILLER_22_153 ();
 FILLCELL_X2 FILLER_22_157 ();
 FILLCELL_X16 FILLER_22_176 ();
 FILLCELL_X8 FILLER_22_192 ();
 FILLCELL_X4 FILLER_22_200 ();
 FILLCELL_X2 FILLER_22_204 ();
 FILLCELL_X1 FILLER_22_206 ();
 FILLCELL_X16 FILLER_22_224 ();
 FILLCELL_X2 FILLER_22_240 ();
 FILLCELL_X1 FILLER_22_242 ();
 FILLCELL_X32 FILLER_22_246 ();
 FILLCELL_X1 FILLER_22_278 ();
 FILLCELL_X4 FILLER_22_282 ();
 FILLCELL_X2 FILLER_22_286 ();
 FILLCELL_X1 FILLER_22_288 ();
 FILLCELL_X32 FILLER_22_292 ();
 FILLCELL_X32 FILLER_22_324 ();
 FILLCELL_X32 FILLER_22_356 ();
 FILLCELL_X16 FILLER_22_388 ();
 FILLCELL_X8 FILLER_22_404 ();
 FILLCELL_X4 FILLER_22_412 ();
 FILLCELL_X2 FILLER_22_416 ();
 FILLCELL_X1 FILLER_22_418 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X16 FILLER_23_129 ();
 FILLCELL_X8 FILLER_23_145 ();
 FILLCELL_X4 FILLER_23_153 ();
 FILLCELL_X32 FILLER_23_160 ();
 FILLCELL_X32 FILLER_23_192 ();
 FILLCELL_X32 FILLER_23_224 ();
 FILLCELL_X16 FILLER_23_256 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X2 FILLER_23_417 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X16 FILLER_24_129 ();
 FILLCELL_X8 FILLER_24_145 ();
 FILLCELL_X1 FILLER_24_153 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X16 FILLER_24_225 ();
 FILLCELL_X1 FILLER_24_241 ();
 FILLCELL_X32 FILLER_24_245 ();
 FILLCELL_X4 FILLER_24_284 ();
 FILLCELL_X1 FILLER_24_288 ();
 FILLCELL_X32 FILLER_24_292 ();
 FILLCELL_X32 FILLER_24_324 ();
 FILLCELL_X32 FILLER_24_356 ();
 FILLCELL_X16 FILLER_24_388 ();
 FILLCELL_X8 FILLER_24_404 ();
 FILLCELL_X4 FILLER_24_412 ();
 FILLCELL_X2 FILLER_24_416 ();
 FILLCELL_X1 FILLER_24_418 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X8 FILLER_25_129 ();
 FILLCELL_X2 FILLER_25_137 ();
 FILLCELL_X1 FILLER_25_139 ();
 FILLCELL_X8 FILLER_25_164 ();
 FILLCELL_X1 FILLER_25_172 ();
 FILLCELL_X8 FILLER_25_190 ();
 FILLCELL_X2 FILLER_25_198 ();
 FILLCELL_X16 FILLER_25_217 ();
 FILLCELL_X8 FILLER_25_233 ();
 FILLCELL_X32 FILLER_25_245 ();
 FILLCELL_X1 FILLER_25_277 ();
 FILLCELL_X2 FILLER_25_284 ();
 FILLCELL_X32 FILLER_25_290 ();
 FILLCELL_X32 FILLER_25_322 ();
 FILLCELL_X32 FILLER_25_354 ();
 FILLCELL_X32 FILLER_25_386 ();
 FILLCELL_X1 FILLER_25_418 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X16 FILLER_26_129 ();
 FILLCELL_X8 FILLER_26_145 ();
 FILLCELL_X2 FILLER_26_153 ();
 FILLCELL_X1 FILLER_26_155 ();
 FILLCELL_X16 FILLER_26_161 ();
 FILLCELL_X2 FILLER_26_177 ();
 FILLCELL_X1 FILLER_26_186 ();
 FILLCELL_X16 FILLER_26_190 ();
 FILLCELL_X4 FILLER_26_216 ();
 FILLCELL_X2 FILLER_26_220 ();
 FILLCELL_X8 FILLER_26_242 ();
 FILLCELL_X2 FILLER_26_250 ();
 FILLCELL_X2 FILLER_26_276 ();
 FILLCELL_X1 FILLER_26_278 ();
 FILLCELL_X32 FILLER_26_299 ();
 FILLCELL_X32 FILLER_26_331 ();
 FILLCELL_X32 FILLER_26_363 ();
 FILLCELL_X16 FILLER_26_395 ();
 FILLCELL_X8 FILLER_26_411 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X4 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_160 ();
 FILLCELL_X16 FILLER_27_192 ();
 FILLCELL_X8 FILLER_27_208 ();
 FILLCELL_X4 FILLER_27_216 ();
 FILLCELL_X2 FILLER_27_220 ();
 FILLCELL_X32 FILLER_27_241 ();
 FILLCELL_X1 FILLER_27_273 ();
 FILLCELL_X32 FILLER_27_290 ();
 FILLCELL_X32 FILLER_27_322 ();
 FILLCELL_X32 FILLER_27_354 ();
 FILLCELL_X32 FILLER_27_386 ();
 FILLCELL_X1 FILLER_27_418 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X2 FILLER_28_161 ();
 FILLCELL_X16 FILLER_28_166 ();
 FILLCELL_X4 FILLER_28_182 ();
 FILLCELL_X1 FILLER_28_186 ();
 FILLCELL_X16 FILLER_28_190 ();
 FILLCELL_X2 FILLER_28_206 ();
 FILLCELL_X1 FILLER_28_208 ();
 FILLCELL_X4 FILLER_28_212 ();
 FILLCELL_X2 FILLER_28_216 ();
 FILLCELL_X1 FILLER_28_218 ();
 FILLCELL_X16 FILLER_28_243 ();
 FILLCELL_X8 FILLER_28_259 ();
 FILLCELL_X16 FILLER_28_270 ();
 FILLCELL_X2 FILLER_28_286 ();
 FILLCELL_X1 FILLER_28_295 ();
 FILLCELL_X32 FILLER_28_299 ();
 FILLCELL_X32 FILLER_28_331 ();
 FILLCELL_X32 FILLER_28_363 ();
 FILLCELL_X16 FILLER_28_395 ();
 FILLCELL_X8 FILLER_28_411 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X8 FILLER_29_129 ();
 FILLCELL_X4 FILLER_29_154 ();
 FILLCELL_X2 FILLER_29_158 ();
 FILLCELL_X16 FILLER_29_167 ();
 FILLCELL_X4 FILLER_29_183 ();
 FILLCELL_X1 FILLER_29_187 ();
 FILLCELL_X32 FILLER_29_213 ();
 FILLCELL_X16 FILLER_29_245 ();
 FILLCELL_X2 FILLER_29_261 ();
 FILLCELL_X1 FILLER_29_263 ();
 FILLCELL_X8 FILLER_29_271 ();
 FILLCELL_X2 FILLER_29_279 ();
 FILLCELL_X32 FILLER_29_322 ();
 FILLCELL_X32 FILLER_29_354 ();
 FILLCELL_X32 FILLER_29_386 ();
 FILLCELL_X1 FILLER_29_418 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X16 FILLER_30_129 ();
 FILLCELL_X2 FILLER_30_145 ();
 FILLCELL_X2 FILLER_30_150 ();
 FILLCELL_X8 FILLER_30_157 ();
 FILLCELL_X1 FILLER_30_186 ();
 FILLCELL_X8 FILLER_30_190 ();
 FILLCELL_X4 FILLER_30_198 ();
 FILLCELL_X1 FILLER_30_202 ();
 FILLCELL_X16 FILLER_30_220 ();
 FILLCELL_X4 FILLER_30_236 ();
 FILLCELL_X8 FILLER_30_243 ();
 FILLCELL_X2 FILLER_30_251 ();
 FILLCELL_X16 FILLER_30_270 ();
 FILLCELL_X4 FILLER_30_286 ();
 FILLCELL_X2 FILLER_30_290 ();
 FILLCELL_X1 FILLER_30_292 ();
 FILLCELL_X32 FILLER_30_309 ();
 FILLCELL_X32 FILLER_30_341 ();
 FILLCELL_X32 FILLER_30_373 ();
 FILLCELL_X8 FILLER_30_405 ();
 FILLCELL_X4 FILLER_30_413 ();
 FILLCELL_X2 FILLER_30_417 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X16 FILLER_31_97 ();
 FILLCELL_X8 FILLER_31_113 ();
 FILLCELL_X2 FILLER_31_121 ();
 FILLCELL_X1 FILLER_31_123 ();
 FILLCELL_X4 FILLER_31_141 ();
 FILLCELL_X2 FILLER_31_145 ();
 FILLCELL_X1 FILLER_31_159 ();
 FILLCELL_X32 FILLER_31_165 ();
 FILLCELL_X1 FILLER_31_197 ();
 FILLCELL_X16 FILLER_31_217 ();
 FILLCELL_X8 FILLER_31_233 ();
 FILLCELL_X4 FILLER_31_241 ();
 FILLCELL_X4 FILLER_31_265 ();
 FILLCELL_X1 FILLER_31_269 ();
 FILLCELL_X16 FILLER_31_273 ();
 FILLCELL_X4 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_299 ();
 FILLCELL_X32 FILLER_31_331 ();
 FILLCELL_X32 FILLER_31_363 ();
 FILLCELL_X16 FILLER_31_395 ();
 FILLCELL_X8 FILLER_31_411 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X4 FILLER_32_129 ();
 FILLCELL_X1 FILLER_32_133 ();
 FILLCELL_X2 FILLER_32_151 ();
 FILLCELL_X1 FILLER_32_153 ();
 FILLCELL_X1 FILLER_32_161 ();
 FILLCELL_X16 FILLER_32_165 ();
 FILLCELL_X8 FILLER_32_181 ();
 FILLCELL_X4 FILLER_32_189 ();
 FILLCELL_X2 FILLER_32_193 ();
 FILLCELL_X1 FILLER_32_195 ();
 FILLCELL_X2 FILLER_32_201 ();
 FILLCELL_X1 FILLER_32_203 ();
 FILLCELL_X16 FILLER_32_207 ();
 FILLCELL_X4 FILLER_32_223 ();
 FILLCELL_X1 FILLER_32_227 ();
 FILLCELL_X8 FILLER_32_231 ();
 FILLCELL_X4 FILLER_32_239 ();
 FILLCELL_X2 FILLER_32_243 ();
 FILLCELL_X16 FILLER_32_270 ();
 FILLCELL_X8 FILLER_32_286 ();
 FILLCELL_X32 FILLER_32_302 ();
 FILLCELL_X32 FILLER_32_334 ();
 FILLCELL_X16 FILLER_32_366 ();
 FILLCELL_X2 FILLER_32_382 ();
 FILLCELL_X1 FILLER_32_384 ();
 FILLCELL_X16 FILLER_32_388 ();
 FILLCELL_X8 FILLER_32_404 ();
 FILLCELL_X4 FILLER_32_412 ();
 FILLCELL_X2 FILLER_32_416 ();
 FILLCELL_X1 FILLER_32_418 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X16 FILLER_33_129 ();
 FILLCELL_X2 FILLER_33_161 ();
 FILLCELL_X8 FILLER_33_166 ();
 FILLCELL_X4 FILLER_33_174 ();
 FILLCELL_X2 FILLER_33_178 ();
 FILLCELL_X32 FILLER_33_183 ();
 FILLCELL_X32 FILLER_33_215 ();
 FILLCELL_X8 FILLER_33_247 ();
 FILLCELL_X16 FILLER_33_275 ();
 FILLCELL_X1 FILLER_33_291 ();
 FILLCELL_X2 FILLER_33_309 ();
 FILLCELL_X8 FILLER_33_314 ();
 FILLCELL_X2 FILLER_33_322 ();
 FILLCELL_X1 FILLER_33_324 ();
 FILLCELL_X2 FILLER_33_332 ();
 FILLCELL_X32 FILLER_33_337 ();
 FILLCELL_X32 FILLER_33_369 ();
 FILLCELL_X16 FILLER_33_401 ();
 FILLCELL_X2 FILLER_33_417 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X2 FILLER_34_129 ();
 FILLCELL_X1 FILLER_34_131 ();
 FILLCELL_X2 FILLER_34_148 ();
 FILLCELL_X1 FILLER_34_150 ();
 FILLCELL_X16 FILLER_34_154 ();
 FILLCELL_X1 FILLER_34_170 ();
 FILLCELL_X2 FILLER_34_199 ();
 FILLCELL_X2 FILLER_34_208 ();
 FILLCELL_X2 FILLER_34_226 ();
 FILLCELL_X1 FILLER_34_228 ();
 FILLCELL_X4 FILLER_34_233 ();
 FILLCELL_X2 FILLER_34_237 ();
 FILLCELL_X1 FILLER_34_239 ();
 FILLCELL_X16 FILLER_34_243 ();
 FILLCELL_X8 FILLER_34_259 ();
 FILLCELL_X1 FILLER_34_267 ();
 FILLCELL_X4 FILLER_34_288 ();
 FILLCELL_X4 FILLER_34_298 ();
 FILLCELL_X2 FILLER_34_302 ();
 FILLCELL_X1 FILLER_34_304 ();
 FILLCELL_X32 FILLER_34_339 ();
 FILLCELL_X32 FILLER_34_371 ();
 FILLCELL_X16 FILLER_34_403 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X16 FILLER_35_129 ();
 FILLCELL_X4 FILLER_35_145 ();
 FILLCELL_X1 FILLER_35_149 ();
 FILLCELL_X16 FILLER_35_154 ();
 FILLCELL_X4 FILLER_35_170 ();
 FILLCELL_X8 FILLER_35_191 ();
 FILLCELL_X2 FILLER_35_199 ();
 FILLCELL_X8 FILLER_35_218 ();
 FILLCELL_X32 FILLER_35_243 ();
 FILLCELL_X16 FILLER_35_275 ();
 FILLCELL_X8 FILLER_35_291 ();
 FILLCELL_X4 FILLER_35_299 ();
 FILLCELL_X2 FILLER_35_303 ();
 FILLCELL_X4 FILLER_35_315 ();
 FILLCELL_X1 FILLER_35_319 ();
 FILLCELL_X32 FILLER_35_330 ();
 FILLCELL_X32 FILLER_35_362 ();
 FILLCELL_X16 FILLER_35_394 ();
 FILLCELL_X8 FILLER_35_410 ();
 FILLCELL_X1 FILLER_35_418 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X16 FILLER_36_129 ();
 FILLCELL_X4 FILLER_36_145 ();
 FILLCELL_X2 FILLER_36_149 ();
 FILLCELL_X32 FILLER_36_170 ();
 FILLCELL_X32 FILLER_36_202 ();
 FILLCELL_X16 FILLER_36_250 ();
 FILLCELL_X8 FILLER_36_266 ();
 FILLCELL_X4 FILLER_36_274 ();
 FILLCELL_X2 FILLER_36_278 ();
 FILLCELL_X1 FILLER_36_280 ();
 FILLCELL_X4 FILLER_36_297 ();
 FILLCELL_X2 FILLER_36_301 ();
 FILLCELL_X1 FILLER_36_303 ();
 FILLCELL_X4 FILLER_36_314 ();
 FILLCELL_X2 FILLER_36_321 ();
 FILLCELL_X1 FILLER_36_323 ();
 FILLCELL_X4 FILLER_36_327 ();
 FILLCELL_X1 FILLER_36_335 ();
 FILLCELL_X16 FILLER_36_356 ();
 FILLCELL_X8 FILLER_36_372 ();
 FILLCELL_X32 FILLER_36_383 ();
 FILLCELL_X4 FILLER_36_415 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X1 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_165 ();
 FILLCELL_X32 FILLER_37_197 ();
 FILLCELL_X32 FILLER_37_229 ();
 FILLCELL_X32 FILLER_37_261 ();
 FILLCELL_X32 FILLER_37_293 ();
 FILLCELL_X8 FILLER_37_325 ();
 FILLCELL_X1 FILLER_37_337 ();
 FILLCELL_X16 FILLER_37_358 ();
 FILLCELL_X8 FILLER_37_374 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X2 FILLER_37_417 ();
 FILLCELL_X16 FILLER_38_1 ();
 FILLCELL_X8 FILLER_38_17 ();
 FILLCELL_X1 FILLER_38_25 ();
 FILLCELL_X32 FILLER_38_29 ();
 FILLCELL_X32 FILLER_38_61 ();
 FILLCELL_X32 FILLER_38_93 ();
 FILLCELL_X8 FILLER_38_125 ();
 FILLCELL_X2 FILLER_38_133 ();
 FILLCELL_X1 FILLER_38_135 ();
 FILLCELL_X16 FILLER_38_152 ();
 FILLCELL_X4 FILLER_38_168 ();
 FILLCELL_X1 FILLER_38_172 ();
 FILLCELL_X16 FILLER_38_183 ();
 FILLCELL_X4 FILLER_38_199 ();
 FILLCELL_X1 FILLER_38_203 ();
 FILLCELL_X8 FILLER_38_214 ();
 FILLCELL_X1 FILLER_38_222 ();
 FILLCELL_X16 FILLER_38_228 ();
 FILLCELL_X2 FILLER_38_244 ();
 FILLCELL_X1 FILLER_38_246 ();
 FILLCELL_X8 FILLER_38_257 ();
 FILLCELL_X1 FILLER_38_265 ();
 FILLCELL_X16 FILLER_38_276 ();
 FILLCELL_X8 FILLER_38_292 ();
 FILLCELL_X4 FILLER_38_300 ();
 FILLCELL_X1 FILLER_38_304 ();
 FILLCELL_X8 FILLER_38_317 ();
 FILLCELL_X1 FILLER_38_325 ();
 FILLCELL_X32 FILLER_38_343 ();
 FILLCELL_X16 FILLER_38_375 ();
 FILLCELL_X4 FILLER_38_391 ();
 FILLCELL_X16 FILLER_38_398 ();
 FILLCELL_X4 FILLER_38_414 ();
 FILLCELL_X1 FILLER_38_418 ();
 FILLCELL_X16 FILLER_39_1 ();
 FILLCELL_X8 FILLER_39_17 ();
 FILLCELL_X2 FILLER_39_25 ();
 FILLCELL_X1 FILLER_39_27 ();
 FILLCELL_X32 FILLER_39_31 ();
 FILLCELL_X32 FILLER_39_63 ();
 FILLCELL_X8 FILLER_39_95 ();
 FILLCELL_X1 FILLER_39_103 ();
 FILLCELL_X32 FILLER_39_121 ();
 FILLCELL_X2 FILLER_39_153 ();
 FILLCELL_X8 FILLER_39_165 ();
 FILLCELL_X1 FILLER_39_173 ();
 FILLCELL_X16 FILLER_39_181 ();
 FILLCELL_X8 FILLER_39_197 ();
 FILLCELL_X16 FILLER_39_212 ();
 FILLCELL_X2 FILLER_39_228 ();
 FILLCELL_X8 FILLER_39_240 ();
 FILLCELL_X8 FILLER_39_252 ();
 FILLCELL_X32 FILLER_39_268 ();
 FILLCELL_X2 FILLER_39_300 ();
 FILLCELL_X1 FILLER_39_311 ();
 FILLCELL_X4 FILLER_39_314 ();
 FILLCELL_X2 FILLER_39_321 ();
 FILLCELL_X1 FILLER_39_323 ();
 FILLCELL_X32 FILLER_39_331 ();
 FILLCELL_X32 FILLER_39_363 ();
 FILLCELL_X16 FILLER_39_395 ();
 FILLCELL_X8 FILLER_39_411 ();
 FILLCELL_X16 FILLER_40_1 ();
 FILLCELL_X8 FILLER_40_17 ();
 FILLCELL_X4 FILLER_40_28 ();
 FILLCELL_X2 FILLER_40_32 ();
 FILLCELL_X32 FILLER_40_37 ();
 FILLCELL_X16 FILLER_40_69 ();
 FILLCELL_X2 FILLER_40_85 ();
 FILLCELL_X16 FILLER_40_112 ();
 FILLCELL_X8 FILLER_40_128 ();
 FILLCELL_X2 FILLER_40_136 ();
 FILLCELL_X1 FILLER_40_138 ();
 FILLCELL_X4 FILLER_40_149 ();
 FILLCELL_X2 FILLER_40_153 ();
 FILLCELL_X1 FILLER_40_155 ();
 FILLCELL_X16 FILLER_40_159 ();
 FILLCELL_X4 FILLER_40_175 ();
 FILLCELL_X32 FILLER_40_183 ();
 FILLCELL_X16 FILLER_40_215 ();
 FILLCELL_X1 FILLER_40_231 ();
 FILLCELL_X2 FILLER_40_243 ();
 FILLCELL_X8 FILLER_40_253 ();
 FILLCELL_X4 FILLER_40_261 ();
 FILLCELL_X2 FILLER_40_265 ();
 FILLCELL_X16 FILLER_40_271 ();
 FILLCELL_X8 FILLER_40_287 ();
 FILLCELL_X2 FILLER_40_295 ();
 FILLCELL_X32 FILLER_40_313 ();
 FILLCELL_X32 FILLER_40_345 ();
 FILLCELL_X32 FILLER_40_377 ();
 FILLCELL_X8 FILLER_40_409 ();
 FILLCELL_X2 FILLER_40_417 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X16 FILLER_41_65 ();
 FILLCELL_X2 FILLER_41_81 ();
 FILLCELL_X16 FILLER_41_112 ();
 FILLCELL_X4 FILLER_41_128 ();
 FILLCELL_X2 FILLER_41_132 ();
 FILLCELL_X4 FILLER_41_144 ();
 FILLCELL_X2 FILLER_41_148 ();
 FILLCELL_X16 FILLER_41_153 ();
 FILLCELL_X2 FILLER_41_169 ();
 FILLCELL_X32 FILLER_41_189 ();
 FILLCELL_X8 FILLER_41_221 ();
 FILLCELL_X2 FILLER_41_229 ();
 FILLCELL_X1 FILLER_41_231 ();
 FILLCELL_X32 FILLER_41_273 ();
 FILLCELL_X32 FILLER_41_305 ();
 FILLCELL_X32 FILLER_41_337 ();
 FILLCELL_X32 FILLER_41_369 ();
 FILLCELL_X16 FILLER_41_401 ();
 FILLCELL_X2 FILLER_41_417 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X16 FILLER_42_65 ();
 FILLCELL_X2 FILLER_42_81 ();
 FILLCELL_X16 FILLER_42_112 ();
 FILLCELL_X4 FILLER_42_128 ();
 FILLCELL_X2 FILLER_42_132 ();
 FILLCELL_X1 FILLER_42_134 ();
 FILLCELL_X1 FILLER_42_144 ();
 FILLCELL_X1 FILLER_42_147 ();
 FILLCELL_X1 FILLER_42_153 ();
 FILLCELL_X2 FILLER_42_159 ();
 FILLCELL_X1 FILLER_42_176 ();
 FILLCELL_X2 FILLER_42_194 ();
 FILLCELL_X32 FILLER_42_199 ();
 FILLCELL_X8 FILLER_42_231 ();
 FILLCELL_X2 FILLER_42_239 ();
 FILLCELL_X4 FILLER_42_249 ();
 FILLCELL_X2 FILLER_42_253 ();
 FILLCELL_X2 FILLER_42_261 ();
 FILLCELL_X1 FILLER_42_263 ();
 FILLCELL_X32 FILLER_42_270 ();
 FILLCELL_X32 FILLER_42_302 ();
 FILLCELL_X32 FILLER_42_334 ();
 FILLCELL_X32 FILLER_42_366 ();
 FILLCELL_X16 FILLER_42_398 ();
 FILLCELL_X4 FILLER_42_414 ();
 FILLCELL_X1 FILLER_42_418 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X8 FILLER_43_129 ();
 FILLCELL_X2 FILLER_43_137 ();
 FILLCELL_X2 FILLER_43_152 ();
 FILLCELL_X1 FILLER_43_166 ();
 FILLCELL_X1 FILLER_43_173 ();
 FILLCELL_X1 FILLER_43_177 ();
 FILLCELL_X16 FILLER_43_182 ();
 FILLCELL_X1 FILLER_43_198 ();
 FILLCELL_X16 FILLER_43_212 ();
 FILLCELL_X8 FILLER_43_228 ();
 FILLCELL_X4 FILLER_43_236 ();
 FILLCELL_X2 FILLER_43_240 ();
 FILLCELL_X1 FILLER_43_242 ();
 FILLCELL_X8 FILLER_43_249 ();
 FILLCELL_X1 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_261 ();
 FILLCELL_X32 FILLER_43_293 ();
 FILLCELL_X32 FILLER_43_325 ();
 FILLCELL_X32 FILLER_43_357 ();
 FILLCELL_X16 FILLER_43_389 ();
 FILLCELL_X8 FILLER_43_405 ();
 FILLCELL_X4 FILLER_43_413 ();
 FILLCELL_X2 FILLER_43_417 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X16 FILLER_44_129 ();
 FILLCELL_X4 FILLER_44_145 ();
 FILLCELL_X2 FILLER_44_149 ();
 FILLCELL_X1 FILLER_44_156 ();
 FILLCELL_X8 FILLER_44_169 ();
 FILLCELL_X4 FILLER_44_177 ();
 FILLCELL_X2 FILLER_44_181 ();
 FILLCELL_X4 FILLER_44_203 ();
 FILLCELL_X1 FILLER_44_207 ();
 FILLCELL_X32 FILLER_44_211 ();
 FILLCELL_X32 FILLER_44_243 ();
 FILLCELL_X32 FILLER_44_275 ();
 FILLCELL_X32 FILLER_44_307 ();
 FILLCELL_X32 FILLER_44_339 ();
 FILLCELL_X32 FILLER_44_371 ();
 FILLCELL_X16 FILLER_44_403 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X16 FILLER_45_129 ();
 FILLCELL_X8 FILLER_45_145 ();
 FILLCELL_X1 FILLER_45_153 ();
 FILLCELL_X1 FILLER_45_162 ();
 FILLCELL_X2 FILLER_45_168 ();
 FILLCELL_X32 FILLER_45_182 ();
 FILLCELL_X32 FILLER_45_214 ();
 FILLCELL_X16 FILLER_45_249 ();
 FILLCELL_X4 FILLER_45_265 ();
 FILLCELL_X32 FILLER_45_272 ();
 FILLCELL_X32 FILLER_45_304 ();
 FILLCELL_X32 FILLER_45_336 ();
 FILLCELL_X32 FILLER_45_368 ();
 FILLCELL_X16 FILLER_45_400 ();
 FILLCELL_X2 FILLER_45_416 ();
 FILLCELL_X1 FILLER_45_418 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X16 FILLER_46_129 ();
 FILLCELL_X8 FILLER_46_145 ();
 FILLCELL_X1 FILLER_46_167 ();
 FILLCELL_X16 FILLER_46_171 ();
 FILLCELL_X8 FILLER_46_187 ();
 FILLCELL_X4 FILLER_46_195 ();
 FILLCELL_X2 FILLER_46_199 ();
 FILLCELL_X32 FILLER_46_206 ();
 FILLCELL_X8 FILLER_46_238 ();
 FILLCELL_X4 FILLER_46_246 ();
 FILLCELL_X2 FILLER_46_250 ();
 FILLCELL_X1 FILLER_46_252 ();
 FILLCELL_X32 FILLER_46_274 ();
 FILLCELL_X32 FILLER_46_306 ();
 FILLCELL_X32 FILLER_46_338 ();
 FILLCELL_X32 FILLER_46_370 ();
 FILLCELL_X16 FILLER_46_402 ();
 FILLCELL_X1 FILLER_46_418 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X2 FILLER_47_167 ();
 FILLCELL_X1 FILLER_47_169 ();
 FILLCELL_X8 FILLER_47_173 ();
 FILLCELL_X4 FILLER_47_181 ();
 FILLCELL_X2 FILLER_47_185 ();
 FILLCELL_X1 FILLER_47_187 ();
 FILLCELL_X4 FILLER_47_199 ();
 FILLCELL_X2 FILLER_47_206 ();
 FILLCELL_X1 FILLER_47_208 ();
 FILLCELL_X16 FILLER_47_216 ();
 FILLCELL_X8 FILLER_47_232 ();
 FILLCELL_X4 FILLER_47_240 ();
 FILLCELL_X1 FILLER_47_248 ();
 FILLCELL_X4 FILLER_47_254 ();
 FILLCELL_X1 FILLER_47_258 ();
 FILLCELL_X2 FILLER_47_266 ();
 FILLCELL_X1 FILLER_47_268 ();
 FILLCELL_X32 FILLER_47_272 ();
 FILLCELL_X32 FILLER_47_304 ();
 FILLCELL_X32 FILLER_47_336 ();
 FILLCELL_X32 FILLER_47_368 ();
 FILLCELL_X16 FILLER_47_400 ();
 FILLCELL_X2 FILLER_47_416 ();
 FILLCELL_X1 FILLER_47_418 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X16 FILLER_48_133 ();
 FILLCELL_X1 FILLER_48_149 ();
 FILLCELL_X16 FILLER_48_167 ();
 FILLCELL_X2 FILLER_48_183 ();
 FILLCELL_X1 FILLER_48_185 ();
 FILLCELL_X16 FILLER_48_220 ();
 FILLCELL_X32 FILLER_48_270 ();
 FILLCELL_X32 FILLER_48_302 ();
 FILLCELL_X32 FILLER_48_334 ();
 FILLCELL_X32 FILLER_48_366 ();
 FILLCELL_X16 FILLER_48_398 ();
 FILLCELL_X4 FILLER_48_414 ();
 FILLCELL_X1 FILLER_48_418 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X16 FILLER_49_129 ();
 FILLCELL_X8 FILLER_49_145 ();
 FILLCELL_X1 FILLER_49_153 ();
 FILLCELL_X32 FILLER_49_174 ();
 FILLCELL_X32 FILLER_49_206 ();
 FILLCELL_X4 FILLER_49_238 ();
 FILLCELL_X2 FILLER_49_242 ();
 FILLCELL_X32 FILLER_49_247 ();
 FILLCELL_X32 FILLER_49_279 ();
 FILLCELL_X32 FILLER_49_311 ();
 FILLCELL_X32 FILLER_49_343 ();
 FILLCELL_X32 FILLER_49_375 ();
 FILLCELL_X8 FILLER_49_407 ();
 FILLCELL_X4 FILLER_49_415 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X4 FILLER_50_257 ();
 FILLCELL_X1 FILLER_50_261 ();
 FILLCELL_X32 FILLER_50_265 ();
 FILLCELL_X32 FILLER_50_297 ();
 FILLCELL_X32 FILLER_50_329 ();
 FILLCELL_X32 FILLER_50_361 ();
 FILLCELL_X16 FILLER_50_393 ();
 FILLCELL_X8 FILLER_50_409 ();
 FILLCELL_X2 FILLER_50_417 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X8 FILLER_51_193 ();
 FILLCELL_X2 FILLER_51_201 ();
 FILLCELL_X32 FILLER_51_209 ();
 FILLCELL_X32 FILLER_51_241 ();
 FILLCELL_X32 FILLER_51_273 ();
 FILLCELL_X32 FILLER_51_305 ();
 FILLCELL_X32 FILLER_51_337 ();
 FILLCELL_X32 FILLER_51_369 ();
 FILLCELL_X16 FILLER_51_401 ();
 FILLCELL_X2 FILLER_51_417 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X16 FILLER_52_161 ();
 FILLCELL_X8 FILLER_52_177 ();
 FILLCELL_X2 FILLER_52_185 ();
 FILLCELL_X1 FILLER_52_187 ();
 FILLCELL_X2 FILLER_52_211 ();
 FILLCELL_X1 FILLER_52_213 ();
 FILLCELL_X2 FILLER_52_218 ();
 FILLCELL_X16 FILLER_52_239 ();
 FILLCELL_X4 FILLER_52_255 ();
 FILLCELL_X32 FILLER_52_276 ();
 FILLCELL_X32 FILLER_52_308 ();
 FILLCELL_X32 FILLER_52_340 ();
 FILLCELL_X32 FILLER_52_372 ();
 FILLCELL_X8 FILLER_52_404 ();
 FILLCELL_X4 FILLER_52_412 ();
 FILLCELL_X2 FILLER_52_416 ();
 FILLCELL_X1 FILLER_52_418 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X16 FILLER_53_161 ();
 FILLCELL_X8 FILLER_53_177 ();
 FILLCELL_X4 FILLER_53_185 ();
 FILLCELL_X1 FILLER_53_189 ();
 FILLCELL_X32 FILLER_53_230 ();
 FILLCELL_X32 FILLER_53_262 ();
 FILLCELL_X32 FILLER_53_294 ();
 FILLCELL_X32 FILLER_53_326 ();
 FILLCELL_X32 FILLER_53_358 ();
 FILLCELL_X16 FILLER_53_390 ();
 FILLCELL_X8 FILLER_53_406 ();
 FILLCELL_X4 FILLER_53_414 ();
 FILLCELL_X1 FILLER_53_418 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X8 FILLER_54_193 ();
 FILLCELL_X4 FILLER_54_201 ();
 FILLCELL_X2 FILLER_54_205 ();
 FILLCELL_X1 FILLER_54_207 ();
 FILLCELL_X32 FILLER_54_211 ();
 FILLCELL_X32 FILLER_54_243 ();
 FILLCELL_X32 FILLER_54_275 ();
 FILLCELL_X32 FILLER_54_307 ();
 FILLCELL_X32 FILLER_54_339 ();
 FILLCELL_X32 FILLER_54_371 ();
 FILLCELL_X16 FILLER_54_403 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X4 FILLER_55_161 ();
 FILLCELL_X1 FILLER_55_165 ();
 FILLCELL_X2 FILLER_55_169 ();
 FILLCELL_X1 FILLER_55_171 ();
 FILLCELL_X16 FILLER_55_175 ();
 FILLCELL_X8 FILLER_55_191 ();
 FILLCELL_X2 FILLER_55_199 ();
 FILLCELL_X2 FILLER_55_204 ();
 FILLCELL_X1 FILLER_55_206 ();
 FILLCELL_X2 FILLER_55_210 ();
 FILLCELL_X2 FILLER_55_218 ();
 FILLCELL_X16 FILLER_55_226 ();
 FILLCELL_X2 FILLER_55_242 ();
 FILLCELL_X1 FILLER_55_244 ();
 FILLCELL_X16 FILLER_55_248 ();
 FILLCELL_X1 FILLER_55_264 ();
 FILLCELL_X1 FILLER_55_268 ();
 FILLCELL_X2 FILLER_55_272 ();
 FILLCELL_X1 FILLER_55_274 ();
 FILLCELL_X32 FILLER_55_278 ();
 FILLCELL_X32 FILLER_55_310 ();
 FILLCELL_X32 FILLER_55_342 ();
 FILLCELL_X32 FILLER_55_374 ();
 FILLCELL_X8 FILLER_55_406 ();
 FILLCELL_X4 FILLER_55_414 ();
 FILLCELL_X1 FILLER_55_418 ();
endmodule
