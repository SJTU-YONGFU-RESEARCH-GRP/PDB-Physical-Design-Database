module sine_cosine_generator (clk,
    enable,
    rst_n,
    valid_out,
    cosine_out,
    phase_in,
    sine_out);
 input clk;
 input enable;
 input rst_n;
 output valid_out;
 output [15:0] cosine_out;
 input [15:0] phase_in;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X2 _323_ (.A(net4),
    .Z(_261_));
 INV_X2 _324_ (.A(_261_),
    .ZN(_309_));
 BUF_X2 _325_ (.A(net5),
    .Z(_262_));
 INV_X2 _326_ (.A(_262_),
    .ZN(_310_));
 BUF_X2 _327_ (.A(rst_n),
    .Z(_263_));
 CLKBUF_X3 _328_ (.A(_263_),
    .Z(_264_));
 BUF_X2 _329_ (.A(enable),
    .Z(_265_));
 CLKBUF_X3 _330_ (.A(_265_),
    .Z(_266_));
 OAI21_X1 _331_ (.A(_264_),
    .B1(_266_),
    .B2(net15),
    .ZN(_267_));
 NOR4_X4 _332_ (.A1(net6),
    .A2(net1),
    .A3(net8),
    .A4(net9),
    .ZN(_268_));
 NOR4_X4 _333_ (.A1(net7),
    .A2(net10),
    .A3(net12),
    .A4(net2),
    .ZN(_269_));
 NOR4_X4 _334_ (.A1(net11),
    .A2(net14),
    .A3(net13),
    .A4(net3),
    .ZN(_270_));
 AND3_X1 _335_ (.A1(_268_),
    .A2(_269_),
    .A3(_270_),
    .ZN(_271_));
 CLKBUF_X3 _336_ (.A(_271_),
    .Z(_272_));
 CLKBUF_X3 _337_ (.A(phase_in[15]),
    .Z(_273_));
 INV_X2 _338_ (.A(_273_),
    .ZN(_274_));
 BUF_X4 _339_ (.A(phase_in[14]),
    .Z(_275_));
 BUF_X4 _340_ (.A(_275_),
    .Z(_276_));
 CLKBUF_X3 _341_ (.A(_311_),
    .Z(_277_));
 INV_X1 _342_ (.A(_277_),
    .ZN(_278_));
 NOR3_X2 _343_ (.A1(_274_),
    .A2(_276_),
    .A3(_278_),
    .ZN(_279_));
 CLKBUF_X3 _344_ (.A(_273_),
    .Z(_280_));
 CLKBUF_X3 _345_ (.A(_321_),
    .Z(_281_));
 NAND2_X2 _346_ (.A1(_275_),
    .A2(_281_),
    .ZN(_282_));
 NOR2_X1 _347_ (.A1(_280_),
    .A2(_282_),
    .ZN(_283_));
 OAI21_X1 _348_ (.A(_272_),
    .B1(_279_),
    .B2(_283_),
    .ZN(_284_));
 NAND4_X1 _349_ (.A1(net1),
    .A2(net8),
    .A3(net7),
    .A4(net12),
    .ZN(_285_));
 NAND4_X1 _350_ (.A1(net14),
    .A2(net13),
    .A3(net3),
    .A4(net2),
    .ZN(_023_));
 NOR2_X1 _351_ (.A1(_285_),
    .A2(_023_),
    .ZN(_024_));
 AND4_X1 _352_ (.A1(net6),
    .A2(net10),
    .A3(net9),
    .A4(net11),
    .ZN(_025_));
 NAND3_X2 _353_ (.A1(_279_),
    .A2(_024_),
    .A3(_025_),
    .ZN(_026_));
 NAND3_X1 _354_ (.A1(_265_),
    .A2(_284_),
    .A3(_026_),
    .ZN(_027_));
 CLKBUF_X3 _355_ (.A(_275_),
    .Z(_028_));
 OR2_X1 _356_ (.A1(_317_),
    .A2(_028_),
    .ZN(_029_));
 NAND2_X1 _357_ (.A1(_028_),
    .A2(_261_),
    .ZN(_030_));
 NAND2_X1 _358_ (.A1(_029_),
    .A2(_030_),
    .ZN(_031_));
 CLKBUF_X3 _359_ (.A(_280_),
    .Z(_032_));
 CLKBUF_X3 _360_ (.A(_319_),
    .Z(_033_));
 NAND2_X2 _361_ (.A1(_275_),
    .A2(_033_),
    .ZN(_034_));
 AOI21_X1 _362_ (.A(_032_),
    .B1(_278_),
    .B2(_034_),
    .ZN(_035_));
 BUF_X1 _363_ (.A(_315_),
    .Z(_036_));
 CLKBUF_X3 _364_ (.A(_036_),
    .Z(_037_));
 AND2_X1 _365_ (.A1(_275_),
    .A2(_277_),
    .ZN(_038_));
 NOR2_X1 _366_ (.A1(_037_),
    .A2(_038_),
    .ZN(_039_));
 INV_X1 _367_ (.A(_275_),
    .ZN(_040_));
 CLKBUF_X3 _368_ (.A(_040_),
    .Z(_041_));
 CLKBUF_X3 _369_ (.A(_041_),
    .Z(_042_));
 CLKBUF_X3 _370_ (.A(_281_),
    .Z(_043_));
 NAND3_X1 _371_ (.A1(_280_),
    .A2(_042_),
    .A3(_043_),
    .ZN(_044_));
 NAND2_X1 _372_ (.A1(_039_),
    .A2(_044_),
    .ZN(_045_));
 OAI21_X1 _373_ (.A(_272_),
    .B1(_035_),
    .B2(_045_),
    .ZN(_046_));
 AOI21_X1 _374_ (.A(_027_),
    .B1(_031_),
    .B2(_046_),
    .ZN(_047_));
 NAND2_X1 _375_ (.A1(_274_),
    .A2(_276_),
    .ZN(_048_));
 CLKBUF_X3 _376_ (.A(_033_),
    .Z(_049_));
 NOR2_X1 _377_ (.A1(_049_),
    .A2(_277_),
    .ZN(_050_));
 AND2_X1 _378_ (.A1(_280_),
    .A2(_034_),
    .ZN(_051_));
 NOR2_X1 _379_ (.A1(_050_),
    .A2(_051_),
    .ZN(_052_));
 OAI221_X1 _380_ (.A(_272_),
    .B1(_048_),
    .B2(_049_),
    .C1(_052_),
    .C2(_043_),
    .ZN(_053_));
 AOI21_X1 _381_ (.A(_267_),
    .B1(_047_),
    .B2(_053_),
    .ZN(_000_));
 OAI21_X1 _382_ (.A(_264_),
    .B1(net16),
    .B2(_266_),
    .ZN(_054_));
 OAI21_X1 _383_ (.A(_282_),
    .B1(_310_),
    .B2(_276_),
    .ZN(_055_));
 BUF_X1 _384_ (.A(_312_),
    .Z(_056_));
 NAND2_X1 _385_ (.A1(_275_),
    .A2(_056_),
    .ZN(_057_));
 OAI21_X1 _386_ (.A(_057_),
    .B1(_262_),
    .B2(_276_),
    .ZN(_058_));
 CLKBUF_X3 _387_ (.A(_274_),
    .Z(_059_));
 MUX2_X1 _388_ (.A(_055_),
    .B(_058_),
    .S(_059_),
    .Z(_060_));
 NAND2_X1 _389_ (.A1(_026_),
    .A2(_060_),
    .ZN(_061_));
 CLKBUF_X3 _390_ (.A(_273_),
    .Z(_062_));
 MUX2_X1 _391_ (.A(_277_),
    .B(_037_),
    .S(_275_),
    .Z(_063_));
 NOR3_X1 _392_ (.A1(_062_),
    .A2(_049_),
    .A3(_063_),
    .ZN(_064_));
 NOR2_X1 _393_ (.A1(_059_),
    .A2(_043_),
    .ZN(_065_));
 NAND2_X1 _394_ (.A1(_041_),
    .A2(_037_),
    .ZN(_066_));
 AOI21_X1 _395_ (.A(_064_),
    .B1(_065_),
    .B2(_066_),
    .ZN(_067_));
 INV_X1 _396_ (.A(_067_),
    .ZN(_068_));
 NAND3_X4 _397_ (.A1(_268_),
    .A2(_269_),
    .A3(_270_),
    .ZN(_069_));
 OAI21_X2 _398_ (.A(_033_),
    .B1(_275_),
    .B2(_274_),
    .ZN(_070_));
 NOR3_X2 _399_ (.A1(_036_),
    .A2(_321_),
    .A3(_311_),
    .ZN(_071_));
 AOI21_X4 _400_ (.A(_069_),
    .B1(_070_),
    .B2(_071_),
    .ZN(_072_));
 MUX2_X1 _401_ (.A(_061_),
    .B(_068_),
    .S(_072_),
    .Z(_073_));
 AOI21_X1 _402_ (.A(_054_),
    .B1(_073_),
    .B2(_266_),
    .ZN(_001_));
 INV_X2 _403_ (.A(_263_),
    .ZN(_074_));
 INV_X2 _404_ (.A(_265_),
    .ZN(_075_));
 NAND2_X1 _405_ (.A1(_075_),
    .A2(net17),
    .ZN(_076_));
 XNOR2_X1 _406_ (.A(_028_),
    .B(_261_),
    .ZN(_077_));
 NAND2_X2 _407_ (.A1(_276_),
    .A2(_037_),
    .ZN(_078_));
 NAND2_X1 _408_ (.A1(_041_),
    .A2(_261_),
    .ZN(_079_));
 NAND2_X1 _409_ (.A1(_078_),
    .A2(_079_),
    .ZN(_080_));
 MUX2_X1 _410_ (.A(_077_),
    .B(_080_),
    .S(_280_),
    .Z(_081_));
 NAND4_X2 _411_ (.A1(net6),
    .A2(net11),
    .A3(net14),
    .A4(net13),
    .ZN(_082_));
 NAND3_X2 _412_ (.A1(net3),
    .A2(net2),
    .A3(_311_),
    .ZN(_083_));
 NAND4_X2 _413_ (.A1(net8),
    .A2(net7),
    .A3(net10),
    .A4(net9),
    .ZN(_084_));
 NAND4_X2 _414_ (.A1(_273_),
    .A2(_040_),
    .A3(net1),
    .A4(net12),
    .ZN(_085_));
 NOR4_X4 _415_ (.A1(_082_),
    .A2(_083_),
    .A3(_084_),
    .A4(_085_),
    .ZN(_086_));
 OR2_X1 _416_ (.A1(_086_),
    .A2(_072_),
    .ZN(_087_));
 BUF_X8 _417_ (.A(_087_),
    .Z(_088_));
 OR2_X1 _418_ (.A1(_036_),
    .A2(_277_),
    .ZN(_089_));
 NOR4_X1 _419_ (.A1(_274_),
    .A2(_276_),
    .A3(_281_),
    .A4(_089_),
    .ZN(_090_));
 OAI21_X1 _420_ (.A(_043_),
    .B1(_041_),
    .B2(_062_),
    .ZN(_091_));
 NOR2_X1 _421_ (.A1(_049_),
    .A2(_089_),
    .ZN(_092_));
 AOI21_X1 _422_ (.A(_090_),
    .B1(_091_),
    .B2(_092_),
    .ZN(_093_));
 NAND2_X1 _423_ (.A1(_062_),
    .A2(_078_),
    .ZN(_094_));
 OAI221_X1 _424_ (.A(_094_),
    .B1(_048_),
    .B2(_043_),
    .C1(_028_),
    .C2(_089_),
    .ZN(_095_));
 NAND3_X1 _425_ (.A1(_272_),
    .A2(_093_),
    .A3(_095_),
    .ZN(_096_));
 CLKBUF_X3 _426_ (.A(_280_),
    .Z(_097_));
 OAI21_X1 _427_ (.A(_044_),
    .B1(_034_),
    .B2(_097_),
    .ZN(_098_));
 OAI221_X1 _428_ (.A(_266_),
    .B1(_081_),
    .B2(_088_),
    .C1(_096_),
    .C2(_098_),
    .ZN(_099_));
 AOI21_X1 _429_ (.A(_074_),
    .B1(_076_),
    .B2(_099_),
    .ZN(_002_));
 NOR2_X4 _430_ (.A1(_086_),
    .A2(_072_),
    .ZN(_100_));
 NAND2_X1 _431_ (.A1(_265_),
    .A2(_263_),
    .ZN(_101_));
 INV_X1 _432_ (.A(_101_),
    .ZN(_102_));
 BUF_X4 _433_ (.A(_102_),
    .Z(_022_));
 OR2_X1 _434_ (.A1(_042_),
    .A2(_313_),
    .ZN(_103_));
 NAND2_X1 _435_ (.A1(_097_),
    .A2(_103_),
    .ZN(_104_));
 NAND4_X1 _436_ (.A1(_048_),
    .A2(_100_),
    .A3(_022_),
    .A4(_104_),
    .ZN(_105_));
 CLKBUF_X3 _437_ (.A(_028_),
    .Z(_106_));
 NAND2_X1 _438_ (.A1(_097_),
    .A2(_106_),
    .ZN(_107_));
 NOR3_X1 _439_ (.A1(_049_),
    .A2(_037_),
    .A3(_043_),
    .ZN(_108_));
 NOR2_X1 _440_ (.A1(_037_),
    .A2(_281_),
    .ZN(_109_));
 AND2_X1 _441_ (.A1(_050_),
    .A2(_109_),
    .ZN(_110_));
 NAND2_X1 _442_ (.A1(_059_),
    .A2(_042_),
    .ZN(_111_));
 OAI22_X1 _443_ (.A1(_107_),
    .A2(_108_),
    .B1(_110_),
    .B2(_111_),
    .ZN(_112_));
 NAND3_X1 _444_ (.A1(_272_),
    .A2(_022_),
    .A3(_112_),
    .ZN(_113_));
 NOR2_X4 _445_ (.A1(_265_),
    .A2(_074_),
    .ZN(_114_));
 NAND2_X1 _446_ (.A1(net18),
    .A2(_114_),
    .ZN(_115_));
 NAND3_X1 _447_ (.A1(_105_),
    .A2(_113_),
    .A3(_115_),
    .ZN(_003_));
 CLKBUF_X3 _448_ (.A(_265_),
    .Z(_116_));
 OAI21_X1 _449_ (.A(_264_),
    .B1(net21),
    .B2(_116_),
    .ZN(_117_));
 NAND2_X1 _450_ (.A1(_280_),
    .A2(_041_),
    .ZN(_118_));
 OAI21_X1 _451_ (.A(_118_),
    .B1(_103_),
    .B2(_097_),
    .ZN(_119_));
 NAND2_X1 _452_ (.A1(_100_),
    .A2(_119_),
    .ZN(_120_));
 NOR2_X1 _453_ (.A1(_049_),
    .A2(_037_),
    .ZN(_121_));
 OAI22_X1 _454_ (.A1(_118_),
    .A2(_109_),
    .B1(_121_),
    .B2(_048_),
    .ZN(_122_));
 AND2_X1 _455_ (.A1(_272_),
    .A2(_122_),
    .ZN(_123_));
 NOR2_X1 _456_ (.A1(_027_),
    .A2(_123_),
    .ZN(_124_));
 AOI21_X1 _457_ (.A(_117_),
    .B1(_120_),
    .B2(_124_),
    .ZN(_004_));
 INV_X1 _458_ (.A(_036_),
    .ZN(_125_));
 OAI21_X1 _459_ (.A(_034_),
    .B1(_125_),
    .B2(_028_),
    .ZN(_126_));
 NAND2_X1 _460_ (.A1(_032_),
    .A2(_126_),
    .ZN(_127_));
 INV_X1 _461_ (.A(_281_),
    .ZN(_128_));
 OAI21_X1 _462_ (.A(_078_),
    .B1(_128_),
    .B2(_028_),
    .ZN(_129_));
 NAND2_X1 _463_ (.A1(_059_),
    .A2(_129_),
    .ZN(_130_));
 AOI21_X2 _464_ (.A(_069_),
    .B1(_127_),
    .B2(_130_),
    .ZN(_131_));
 AND2_X1 _465_ (.A1(_041_),
    .A2(_033_),
    .ZN(_132_));
 AOI21_X1 _466_ (.A(_132_),
    .B1(_310_),
    .B2(_106_),
    .ZN(_133_));
 MUX2_X1 _467_ (.A(_056_),
    .B(_133_),
    .S(_059_),
    .Z(_134_));
 OAI221_X1 _468_ (.A(_022_),
    .B1(_131_),
    .B2(_096_),
    .C1(_134_),
    .C2(_088_),
    .ZN(_135_));
 NAND3_X1 _469_ (.A1(_075_),
    .A2(net22),
    .A3(_264_),
    .ZN(_136_));
 NAND2_X1 _470_ (.A1(_135_),
    .A2(_136_),
    .ZN(_005_));
 OAI21_X1 _471_ (.A(_264_),
    .B1(net29),
    .B2(_116_),
    .ZN(_137_));
 OAI21_X1 _472_ (.A(_282_),
    .B1(_278_),
    .B2(_028_),
    .ZN(_138_));
 NAND3_X1 _473_ (.A1(_059_),
    .A2(_272_),
    .A3(_138_),
    .ZN(_139_));
 NAND3_X1 _474_ (.A1(_116_),
    .A2(_026_),
    .A3(_139_),
    .ZN(_140_));
 NOR2_X1 _475_ (.A1(_123_),
    .A2(_140_),
    .ZN(_141_));
 CLKBUF_X3 _476_ (.A(_059_),
    .Z(_142_));
 NOR3_X1 _477_ (.A1(_142_),
    .A2(_106_),
    .A3(_313_),
    .ZN(_143_));
 NAND2_X1 _478_ (.A1(_042_),
    .A2(_277_),
    .ZN(_144_));
 AOI21_X1 _479_ (.A(_097_),
    .B1(_144_),
    .B2(_103_),
    .ZN(_145_));
 OAI21_X1 _480_ (.A(_100_),
    .B1(_143_),
    .B2(_145_),
    .ZN(_146_));
 AOI21_X1 _481_ (.A(_137_),
    .B1(_141_),
    .B2(_146_),
    .ZN(_006_));
 OAI21_X1 _482_ (.A(_264_),
    .B1(net26),
    .B2(_116_),
    .ZN(_147_));
 NOR2_X1 _483_ (.A1(_131_),
    .A2(_140_),
    .ZN(_148_));
 INV_X1 _484_ (.A(_056_),
    .ZN(_149_));
 NAND2_X1 _485_ (.A1(_041_),
    .A2(_149_),
    .ZN(_150_));
 NAND2_X1 _486_ (.A1(_028_),
    .A2(_262_),
    .ZN(_151_));
 AOI21_X1 _487_ (.A(_280_),
    .B1(_150_),
    .B2(_151_),
    .ZN(_152_));
 OAI21_X1 _488_ (.A(_034_),
    .B1(_149_),
    .B2(_106_),
    .ZN(_153_));
 AOI21_X1 _489_ (.A(_152_),
    .B1(_153_),
    .B2(_032_),
    .ZN(_154_));
 OR2_X1 _490_ (.A1(_088_),
    .A2(_154_),
    .ZN(_155_));
 AOI21_X1 _491_ (.A(_147_),
    .B1(_148_),
    .B2(_155_),
    .ZN(_007_));
 OAI21_X1 _492_ (.A(_263_),
    .B1(net19),
    .B2(_116_),
    .ZN(_156_));
 NAND3_X1 _493_ (.A1(_280_),
    .A2(_030_),
    .A3(_066_),
    .ZN(_157_));
 NAND3_X1 _494_ (.A1(_059_),
    .A2(_029_),
    .A3(_078_),
    .ZN(_158_));
 NAND3_X1 _495_ (.A1(_026_),
    .A2(_157_),
    .A3(_158_),
    .ZN(_159_));
 NOR2_X1 _496_ (.A1(_276_),
    .A2(_277_),
    .ZN(_160_));
 NOR2_X1 _497_ (.A1(_033_),
    .A2(_281_),
    .ZN(_161_));
 AOI221_X1 _498_ (.A(_273_),
    .B1(_276_),
    .B2(_125_),
    .C1(_160_),
    .C2(_161_),
    .ZN(_162_));
 OAI21_X1 _499_ (.A(_066_),
    .B1(_161_),
    .B2(_042_),
    .ZN(_163_));
 AOI21_X1 _500_ (.A(_162_),
    .B1(_163_),
    .B2(_032_),
    .ZN(_164_));
 MUX2_X1 _501_ (.A(_159_),
    .B(_164_),
    .S(_072_),
    .Z(_165_));
 AOI21_X1 _502_ (.A(_156_),
    .B1(_165_),
    .B2(_266_),
    .ZN(_008_));
 NAND2_X1 _503_ (.A1(_042_),
    .A2(_043_),
    .ZN(_166_));
 AOI21_X1 _504_ (.A(_051_),
    .B1(_166_),
    .B2(_142_),
    .ZN(_167_));
 MUX2_X1 _505_ (.A(_041_),
    .B(_262_),
    .S(_261_),
    .Z(_168_));
 NOR2_X1 _506_ (.A1(_032_),
    .A2(_168_),
    .ZN(_169_));
 AOI21_X1 _507_ (.A(_132_),
    .B1(_056_),
    .B2(_106_),
    .ZN(_170_));
 AOI21_X1 _508_ (.A(_169_),
    .B1(_170_),
    .B2(_097_),
    .ZN(_171_));
 OAI221_X1 _509_ (.A(_266_),
    .B1(_096_),
    .B2(_167_),
    .C1(_171_),
    .C2(_088_),
    .ZN(_172_));
 NAND2_X1 _510_ (.A1(_075_),
    .A2(net28),
    .ZN(_173_));
 AOI21_X1 _511_ (.A(_074_),
    .B1(_172_),
    .B2(_173_),
    .ZN(_009_));
 NAND3_X1 _512_ (.A1(_097_),
    .A2(_166_),
    .A3(_151_),
    .ZN(_174_));
 MUX2_X1 _513_ (.A(_106_),
    .B(_262_),
    .S(_261_),
    .Z(_175_));
 NAND2_X1 _514_ (.A1(_142_),
    .A2(_175_),
    .ZN(_176_));
 NAND4_X1 _515_ (.A1(_100_),
    .A2(_022_),
    .A3(_174_),
    .A4(_176_),
    .ZN(_177_));
 AOI21_X1 _516_ (.A(_049_),
    .B1(_089_),
    .B2(_042_),
    .ZN(_178_));
 AOI22_X1 _517_ (.A1(_065_),
    .A2(_078_),
    .B1(_178_),
    .B2(_142_),
    .ZN(_179_));
 NAND3_X1 _518_ (.A1(_272_),
    .A2(_022_),
    .A3(_179_),
    .ZN(_180_));
 NAND2_X1 _519_ (.A1(net20),
    .A2(_114_),
    .ZN(_181_));
 NAND3_X1 _520_ (.A1(_177_),
    .A2(_180_),
    .A3(_181_),
    .ZN(_010_));
 NAND2_X1 _521_ (.A1(net31),
    .A2(_114_),
    .ZN(_182_));
 OAI21_X2 _522_ (.A(_079_),
    .B1(_042_),
    .B2(_317_),
    .ZN(_183_));
 OAI21_X1 _523_ (.A(_106_),
    .B1(_049_),
    .B2(_277_),
    .ZN(_184_));
 AOI21_X1 _524_ (.A(_043_),
    .B1(_049_),
    .B2(_142_),
    .ZN(_185_));
 NAND3_X1 _525_ (.A1(_089_),
    .A2(_184_),
    .A3(_185_),
    .ZN(_186_));
 OAI221_X2 _526_ (.A(_022_),
    .B1(_183_),
    .B2(_088_),
    .C1(_186_),
    .C2(_069_),
    .ZN(_187_));
 NAND2_X1 _527_ (.A1(_182_),
    .A2(_187_),
    .ZN(_011_));
 NAND3_X1 _528_ (.A1(_075_),
    .A2(net32),
    .A3(_264_),
    .ZN(_188_));
 MUX2_X1 _529_ (.A(_277_),
    .B(_281_),
    .S(_273_),
    .Z(_189_));
 NAND2_X1 _530_ (.A1(_276_),
    .A2(_189_),
    .ZN(_190_));
 NAND2_X1 _531_ (.A1(_062_),
    .A2(_125_),
    .ZN(_191_));
 MUX2_X2 _532_ (.A(_281_),
    .B(_033_),
    .S(_275_),
    .Z(_192_));
 OAI21_X1 _533_ (.A(_191_),
    .B1(_192_),
    .B2(_032_),
    .ZN(_193_));
 NAND3_X1 _534_ (.A1(_072_),
    .A2(_190_),
    .A3(_193_),
    .ZN(_194_));
 NAND2_X1 _535_ (.A1(_022_),
    .A2(_194_),
    .ZN(_195_));
 NAND2_X1 _536_ (.A1(_106_),
    .A2(_310_),
    .ZN(_196_));
 NAND3_X1 _537_ (.A1(_032_),
    .A2(_196_),
    .A3(_150_),
    .ZN(_197_));
 OAI21_X1 _538_ (.A(_151_),
    .B1(_043_),
    .B2(_106_),
    .ZN(_198_));
 OAI21_X1 _539_ (.A(_197_),
    .B1(_198_),
    .B2(_097_),
    .ZN(_199_));
 NOR2_X1 _540_ (.A1(_088_),
    .A2(_199_),
    .ZN(_200_));
 OAI21_X1 _541_ (.A(_188_),
    .B1(_195_),
    .B2(_200_),
    .ZN(_012_));
 NAND2_X1 _542_ (.A1(net33),
    .A2(_114_),
    .ZN(_201_));
 NAND2_X1 _543_ (.A1(_062_),
    .A2(_192_),
    .ZN(_202_));
 NAND2_X1 _544_ (.A1(_072_),
    .A2(_202_),
    .ZN(_203_));
 NAND2_X1 _545_ (.A1(_059_),
    .A2(_037_),
    .ZN(_204_));
 AOI21_X1 _546_ (.A(_069_),
    .B1(_190_),
    .B2(_204_),
    .ZN(_205_));
 NOR2_X1 _547_ (.A1(_142_),
    .A2(_261_),
    .ZN(_206_));
 AOI21_X1 _548_ (.A(_206_),
    .B1(_039_),
    .B2(_142_),
    .ZN(_207_));
 OAI221_X2 _549_ (.A(_022_),
    .B1(_203_),
    .B2(_205_),
    .C1(_207_),
    .C2(_088_),
    .ZN(_208_));
 NAND2_X1 _550_ (.A1(_201_),
    .A2(_208_),
    .ZN(_013_));
 AOI21_X1 _551_ (.A(_062_),
    .B1(_039_),
    .B2(_161_),
    .ZN(_209_));
 NAND2_X1 _552_ (.A1(_042_),
    .A2(_313_),
    .ZN(_210_));
 AOI221_X2 _553_ (.A(_075_),
    .B1(_271_),
    .B2(_209_),
    .C1(_210_),
    .C2(_100_),
    .ZN(_211_));
 NOR2_X1 _554_ (.A1(_142_),
    .A2(_075_),
    .ZN(_212_));
 OAI21_X1 _555_ (.A(_263_),
    .B1(net34),
    .B2(_116_),
    .ZN(_213_));
 NOR3_X1 _556_ (.A1(_211_),
    .A2(_212_),
    .A3(_213_),
    .ZN(_014_));
 NAND3_X1 _557_ (.A1(_075_),
    .A2(net36),
    .A3(_264_),
    .ZN(_214_));
 OAI21_X1 _558_ (.A(_142_),
    .B1(_037_),
    .B2(_192_),
    .ZN(_215_));
 NAND3_X1 _559_ (.A1(_072_),
    .A2(_190_),
    .A3(_215_),
    .ZN(_216_));
 NAND2_X1 _560_ (.A1(_022_),
    .A2(_216_),
    .ZN(_217_));
 MUX2_X1 _561_ (.A(_049_),
    .B(_043_),
    .S(_028_),
    .Z(_218_));
 NAND2_X1 _562_ (.A1(_032_),
    .A2(_218_),
    .ZN(_219_));
 OAI21_X1 _563_ (.A(_282_),
    .B1(_262_),
    .B2(_106_),
    .ZN(_220_));
 OAI21_X1 _564_ (.A(_219_),
    .B1(_220_),
    .B2(_097_),
    .ZN(_221_));
 NOR2_X1 _565_ (.A1(_088_),
    .A2(_221_),
    .ZN(_222_));
 OAI21_X1 _566_ (.A(_214_),
    .B1(_217_),
    .B2(_222_),
    .ZN(_015_));
 OAI21_X1 _567_ (.A(_263_),
    .B1(net37),
    .B2(_116_),
    .ZN(_223_));
 NAND3_X1 _568_ (.A1(_097_),
    .A2(_100_),
    .A3(_210_),
    .ZN(_224_));
 NAND2_X1 _569_ (.A1(_116_),
    .A2(_026_),
    .ZN(_225_));
 AOI21_X1 _570_ (.A(_142_),
    .B1(_109_),
    .B2(_184_),
    .ZN(_226_));
 AOI21_X1 _571_ (.A(_225_),
    .B1(_226_),
    .B2(_272_),
    .ZN(_227_));
 AOI21_X1 _572_ (.A(_223_),
    .B1(_224_),
    .B2(_227_),
    .ZN(_016_));
 OAI21_X1 _573_ (.A(_263_),
    .B1(net38),
    .B2(_116_),
    .ZN(_228_));
 AOI21_X1 _574_ (.A(_062_),
    .B1(_034_),
    .B2(_150_),
    .ZN(_229_));
 NAND2_X1 _575_ (.A1(_041_),
    .A2(_262_),
    .ZN(_230_));
 AND3_X1 _576_ (.A1(_062_),
    .A2(_230_),
    .A3(_057_),
    .ZN(_231_));
 OR3_X1 _577_ (.A1(_086_),
    .A2(_229_),
    .A3(_231_),
    .ZN(_232_));
 NOR3_X2 _578_ (.A1(_273_),
    .A2(_276_),
    .A3(_033_),
    .ZN(_233_));
 NOR2_X1 _579_ (.A1(_274_),
    .A2(_192_),
    .ZN(_234_));
 NOR4_X2 _580_ (.A1(_273_),
    .A2(_041_),
    .A3(_281_),
    .A4(_277_),
    .ZN(_235_));
 NOR3_X1 _581_ (.A1(_233_),
    .A2(_234_),
    .A3(_235_),
    .ZN(_236_));
 NOR2_X1 _582_ (.A1(_037_),
    .A2(_236_),
    .ZN(_237_));
 MUX2_X1 _583_ (.A(_232_),
    .B(_237_),
    .S(_072_),
    .Z(_238_));
 AOI21_X1 _584_ (.A(_228_),
    .B1(_238_),
    .B2(_266_),
    .ZN(_017_));
 OAI21_X1 _585_ (.A(_264_),
    .B1(net45),
    .B2(_266_),
    .ZN(_239_));
 OAI21_X1 _586_ (.A(_190_),
    .B1(_125_),
    .B2(_059_),
    .ZN(_240_));
 AOI221_X2 _587_ (.A(_203_),
    .B1(_240_),
    .B2(_271_),
    .C1(_114_),
    .C2(net45),
    .ZN(_241_));
 NAND2_X1 _588_ (.A1(_280_),
    .A2(_313_),
    .ZN(_242_));
 OR2_X1 _589_ (.A1(_062_),
    .A2(_038_),
    .ZN(_243_));
 AOI221_X1 _590_ (.A(_088_),
    .B1(_242_),
    .B2(_243_),
    .C1(_114_),
    .C2(net45),
    .ZN(_244_));
 NOR3_X1 _591_ (.A1(_239_),
    .A2(_241_),
    .A3(_244_),
    .ZN(_018_));
 NOR2_X1 _592_ (.A1(_191_),
    .A2(_192_),
    .ZN(_245_));
 NOR4_X1 _593_ (.A1(_069_),
    .A2(_233_),
    .A3(_235_),
    .A4(_245_),
    .ZN(_246_));
 AOI22_X1 _594_ (.A1(net42),
    .A2(_114_),
    .B1(_246_),
    .B2(_102_),
    .ZN(_247_));
 NOR2_X1 _595_ (.A1(_042_),
    .A2(_056_),
    .ZN(_248_));
 NOR3_X1 _596_ (.A1(_032_),
    .A2(_132_),
    .A3(_248_),
    .ZN(_249_));
 OR3_X1 _597_ (.A1(_101_),
    .A2(_231_),
    .A3(_249_),
    .ZN(_250_));
 OAI21_X1 _598_ (.A(_247_),
    .B1(_250_),
    .B2(_088_),
    .ZN(_019_));
 OAI21_X1 _599_ (.A(_263_),
    .B1(net35),
    .B2(_116_),
    .ZN(_251_));
 OR4_X1 _600_ (.A1(_062_),
    .A2(_033_),
    .A3(_281_),
    .A4(_038_),
    .ZN(_252_));
 NAND3_X1 _601_ (.A1(_272_),
    .A2(_191_),
    .A3(_252_),
    .ZN(_253_));
 OAI21_X1 _602_ (.A(_191_),
    .B1(_183_),
    .B2(_032_),
    .ZN(_254_));
 MUX2_X1 _603_ (.A(_253_),
    .B(_254_),
    .S(_100_),
    .Z(_255_));
 AOI21_X1 _604_ (.A(_251_),
    .B1(_255_),
    .B2(_266_),
    .ZN(_020_));
 OAI21_X1 _605_ (.A(_125_),
    .B1(_233_),
    .B2(_235_),
    .ZN(_256_));
 NOR2_X1 _606_ (.A1(_069_),
    .A2(_234_),
    .ZN(_257_));
 NOR2_X1 _607_ (.A1(_229_),
    .A2(_234_),
    .ZN(_258_));
 AOI221_X2 _608_ (.A(_075_),
    .B1(_256_),
    .B2(_257_),
    .C1(_258_),
    .C2(_100_),
    .ZN(_259_));
 OAI21_X1 _609_ (.A(_264_),
    .B1(net44),
    .B2(_266_),
    .ZN(_260_));
 NOR2_X1 _610_ (.A1(_259_),
    .A2(_260_),
    .ZN(_021_));
 HA_X1 _611_ (.A(_309_),
    .B(_310_),
    .CO(_311_),
    .S(_312_));
 HA_X1 _612_ (.A(_309_),
    .B(_310_),
    .CO(_313_),
    .S(_314_));
 HA_X1 _613_ (.A(_309_),
    .B(net5),
    .CO(_315_),
    .S(_316_));
 HA_X1 _614_ (.A(_309_),
    .B(net5),
    .CO(_317_),
    .S(_318_));
 HA_X1 _615_ (.A(net4),
    .B(_310_),
    .CO(_319_),
    .S(_320_));
 HA_X1 _616_ (.A(net4),
    .B(net5),
    .CO(_321_),
    .S(_322_));
 BUF_X1 _617_ (.A(net29),
    .Z(net23));
 BUF_X1 _618_ (.A(net26),
    .Z(net24));
 BUF_X1 _619_ (.A(net26),
    .Z(net25));
 BUF_X1 _620_ (.A(net19),
    .Z(net27));
 BUF_X1 _621_ (.A(net20),
    .Z(net30));
 BUF_X1 _622_ (.A(net45),
    .Z(net39));
 BUF_X1 _623_ (.A(net42),
    .Z(net40));
 BUF_X1 _624_ (.A(net42),
    .Z(net41));
 BUF_X1 _625_ (.A(net35),
    .Z(net43));
 BUF_X1 _626_ (.A(net36),
    .Z(net46));
 DFF_X1 \cosine_out[0]$_SDFFE_PN0P_  (.D(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net15),
    .QN(_308_));
 DFF_X1 \cosine_out[10]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net16),
    .QN(_307_));
 DFF_X1 \cosine_out[11]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net17),
    .QN(_306_));
 DFF_X1 \cosine_out[12]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net18),
    .QN(_305_));
 DFF_X1 \cosine_out[15]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net21),
    .QN(_304_));
 DFF_X1 \cosine_out[1]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net22),
    .QN(_303_));
 DFF_X1 \cosine_out[2]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net29),
    .QN(_302_));
 DFF_X1 \cosine_out[5]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net26),
    .QN(_301_));
 DFF_X1 \cosine_out[6]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net19),
    .QN(_300_));
 DFF_X1 \cosine_out[7]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net28),
    .QN(_299_));
 DFF_X1 \cosine_out[9]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net20),
    .QN(_298_));
 DFF_X1 \sine_out[0]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net31),
    .QN(_297_));
 DFF_X1 \sine_out[10]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net32),
    .QN(_296_));
 DFF_X1 \sine_out[11]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net33),
    .QN(_295_));
 DFF_X1 \sine_out[12]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net34),
    .QN(_294_));
 DFF_X1 \sine_out[14]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net36),
    .QN(_293_));
 DFF_X1 \sine_out[15]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net37),
    .QN(_292_));
 DFF_X1 \sine_out[1]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net38),
    .QN(_291_));
 DFF_X2 \sine_out[2]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net45),
    .QN(_290_));
 DFF_X1 \sine_out[5]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net42),
    .QN(_289_));
 DFF_X1 \sine_out[6]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net35),
    .QN(_288_));
 DFF_X1 \sine_out[7]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net44),
    .QN(_287_));
 DFF_X1 \valid_out$_SDFF_PN0_  (.D(_022_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net47),
    .QN(_286_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_65 ();
 BUF_X2 input1 (.A(phase_in[0]),
    .Z(net1));
 BUF_X2 input2 (.A(phase_in[10]),
    .Z(net2));
 CLKBUF_X2 input3 (.A(phase_in[11]),
    .Z(net3));
 BUF_X1 input4 (.A(phase_in[12]),
    .Z(net4));
 BUF_X2 input5 (.A(phase_in[13]),
    .Z(net5));
 CLKBUF_X2 input6 (.A(phase_in[1]),
    .Z(net6));
 BUF_X2 input7 (.A(phase_in[2]),
    .Z(net7));
 CLKBUF_X2 input8 (.A(phase_in[3]),
    .Z(net8));
 CLKBUF_X2 input9 (.A(phase_in[4]),
    .Z(net9));
 CLKBUF_X2 input10 (.A(phase_in[5]),
    .Z(net10));
 CLKBUF_X2 input11 (.A(phase_in[6]),
    .Z(net11));
 BUF_X2 input12 (.A(phase_in[7]),
    .Z(net12));
 CLKBUF_X2 input13 (.A(phase_in[8]),
    .Z(net13));
 CLKBUF_X2 input14 (.A(phase_in[9]),
    .Z(net14));
 BUF_X1 output15 (.A(net15),
    .Z(cosine_out[0]));
 BUF_X1 output16 (.A(net16),
    .Z(cosine_out[10]));
 BUF_X1 output17 (.A(net17),
    .Z(cosine_out[11]));
 BUF_X1 output18 (.A(net18),
    .Z(cosine_out[12]));
 BUF_X1 output19 (.A(net19),
    .Z(cosine_out[13]));
 BUF_X1 output20 (.A(net20),
    .Z(cosine_out[14]));
 BUF_X1 output21 (.A(net21),
    .Z(cosine_out[15]));
 BUF_X1 output22 (.A(net22),
    .Z(cosine_out[1]));
 BUF_X1 output23 (.A(net23),
    .Z(cosine_out[2]));
 BUF_X1 output24 (.A(net24),
    .Z(cosine_out[3]));
 BUF_X1 output25 (.A(net25),
    .Z(cosine_out[4]));
 BUF_X1 output26 (.A(net26),
    .Z(cosine_out[5]));
 BUF_X1 output27 (.A(net27),
    .Z(cosine_out[6]));
 BUF_X1 output28 (.A(net28),
    .Z(cosine_out[7]));
 BUF_X1 output29 (.A(net29),
    .Z(cosine_out[8]));
 BUF_X1 output30 (.A(net30),
    .Z(cosine_out[9]));
 BUF_X1 output31 (.A(net31),
    .Z(sine_out[0]));
 BUF_X1 output32 (.A(net32),
    .Z(sine_out[10]));
 BUF_X1 output33 (.A(net33),
    .Z(sine_out[11]));
 BUF_X1 output34 (.A(net34),
    .Z(sine_out[12]));
 BUF_X1 output35 (.A(net35),
    .Z(sine_out[13]));
 BUF_X1 output36 (.A(net36),
    .Z(sine_out[14]));
 BUF_X1 output37 (.A(net37),
    .Z(sine_out[15]));
 BUF_X1 output38 (.A(net38),
    .Z(sine_out[1]));
 BUF_X1 output39 (.A(net39),
    .Z(sine_out[2]));
 BUF_X1 output40 (.A(net40),
    .Z(sine_out[3]));
 BUF_X1 output41 (.A(net41),
    .Z(sine_out[4]));
 BUF_X1 output42 (.A(net42),
    .Z(sine_out[5]));
 BUF_X1 output43 (.A(net43),
    .Z(sine_out[6]));
 BUF_X1 output44 (.A(net44),
    .Z(sine_out[7]));
 BUF_X1 output45 (.A(net45),
    .Z(sine_out[8]));
 BUF_X1 output46 (.A(net46),
    .Z(sine_out[9]));
 BUF_X1 output47 (.A(net47),
    .Z(valid_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_33 ();
 FILLCELL_X2 FILLER_0_41 ();
 FILLCELL_X1 FILLER_0_43 ();
 FILLCELL_X32 FILLER_0_56 ();
 FILLCELL_X16 FILLER_0_88 ();
 FILLCELL_X8 FILLER_0_104 ();
 FILLCELL_X4 FILLER_0_112 ();
 FILLCELL_X2 FILLER_0_116 ();
 FILLCELL_X32 FILLER_0_133 ();
 FILLCELL_X2 FILLER_0_165 ();
 FILLCELL_X1 FILLER_0_167 ();
 FILLCELL_X32 FILLER_0_177 ();
 FILLCELL_X32 FILLER_0_209 ();
 FILLCELL_X8 FILLER_0_241 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X8 FILLER_1_33 ();
 FILLCELL_X4 FILLER_1_41 ();
 FILLCELL_X1 FILLER_1_45 ();
 FILLCELL_X32 FILLER_1_50 ();
 FILLCELL_X32 FILLER_1_82 ();
 FILLCELL_X32 FILLER_1_114 ();
 FILLCELL_X2 FILLER_1_146 ();
 FILLCELL_X32 FILLER_1_151 ();
 FILLCELL_X32 FILLER_1_183 ();
 FILLCELL_X32 FILLER_1_215 ();
 FILLCELL_X2 FILLER_1_247 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X16 FILLER_2_225 ();
 FILLCELL_X8 FILLER_2_241 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X4 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_150 ();
 FILLCELL_X32 FILLER_3_182 ();
 FILLCELL_X32 FILLER_3_214 ();
 FILLCELL_X2 FILLER_3_246 ();
 FILLCELL_X1 FILLER_3_248 ();
 FILLCELL_X4 FILLER_4_1 ();
 FILLCELL_X2 FILLER_4_5 ();
 FILLCELL_X1 FILLER_4_7 ();
 FILLCELL_X8 FILLER_4_12 ();
 FILLCELL_X2 FILLER_4_20 ();
 FILLCELL_X1 FILLER_4_22 ();
 FILLCELL_X32 FILLER_4_50 ();
 FILLCELL_X16 FILLER_4_82 ();
 FILLCELL_X8 FILLER_4_98 ();
 FILLCELL_X2 FILLER_4_106 ();
 FILLCELL_X8 FILLER_4_125 ();
 FILLCELL_X4 FILLER_4_133 ();
 FILLCELL_X1 FILLER_4_137 ();
 FILLCELL_X1 FILLER_4_142 ();
 FILLCELL_X32 FILLER_4_147 ();
 FILLCELL_X32 FILLER_4_179 ();
 FILLCELL_X32 FILLER_4_211 ();
 FILLCELL_X4 FILLER_4_243 ();
 FILLCELL_X2 FILLER_4_247 ();
 FILLCELL_X4 FILLER_5_13 ();
 FILLCELL_X4 FILLER_5_26 ();
 FILLCELL_X1 FILLER_5_30 ();
 FILLCELL_X2 FILLER_5_37 ();
 FILLCELL_X1 FILLER_5_39 ();
 FILLCELL_X32 FILLER_5_63 ();
 FILLCELL_X32 FILLER_5_95 ();
 FILLCELL_X16 FILLER_5_127 ();
 FILLCELL_X4 FILLER_5_143 ();
 FILLCELL_X2 FILLER_5_147 ();
 FILLCELL_X16 FILLER_5_168 ();
 FILLCELL_X8 FILLER_5_184 ();
 FILLCELL_X4 FILLER_5_192 ();
 FILLCELL_X1 FILLER_5_196 ();
 FILLCELL_X32 FILLER_5_217 ();
 FILLCELL_X1 FILLER_6_1 ();
 FILLCELL_X16 FILLER_6_25 ();
 FILLCELL_X8 FILLER_6_41 ();
 FILLCELL_X16 FILLER_6_67 ();
 FILLCELL_X4 FILLER_6_83 ();
 FILLCELL_X2 FILLER_6_87 ();
 FILLCELL_X4 FILLER_6_102 ();
 FILLCELL_X2 FILLER_6_110 ();
 FILLCELL_X32 FILLER_6_117 ();
 FILLCELL_X4 FILLER_6_149 ();
 FILLCELL_X2 FILLER_6_153 ();
 FILLCELL_X16 FILLER_6_169 ();
 FILLCELL_X8 FILLER_6_185 ();
 FILLCELL_X4 FILLER_6_193 ();
 FILLCELL_X2 FILLER_6_197 ();
 FILLCELL_X1 FILLER_6_199 ();
 FILLCELL_X4 FILLER_6_203 ();
 FILLCELL_X8 FILLER_6_211 ();
 FILLCELL_X4 FILLER_6_219 ();
 FILLCELL_X1 FILLER_6_223 ();
 FILLCELL_X4 FILLER_6_241 ();
 FILLCELL_X1 FILLER_6_245 ();
 FILLCELL_X4 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_9 ();
 FILLCELL_X2 FILLER_7_13 ();
 FILLCELL_X4 FILLER_7_19 ();
 FILLCELL_X4 FILLER_7_34 ();
 FILLCELL_X2 FILLER_7_38 ();
 FILLCELL_X1 FILLER_7_40 ();
 FILLCELL_X32 FILLER_7_44 ();
 FILLCELL_X8 FILLER_7_76 ();
 FILLCELL_X8 FILLER_7_88 ();
 FILLCELL_X1 FILLER_7_96 ();
 FILLCELL_X1 FILLER_7_116 ();
 FILLCELL_X16 FILLER_7_130 ();
 FILLCELL_X4 FILLER_7_146 ();
 FILLCELL_X2 FILLER_7_150 ();
 FILLCELL_X32 FILLER_7_163 ();
 FILLCELL_X16 FILLER_7_195 ();
 FILLCELL_X8 FILLER_7_216 ();
 FILLCELL_X1 FILLER_7_224 ();
 FILLCELL_X1 FILLER_7_229 ();
 FILLCELL_X8 FILLER_7_234 ();
 FILLCELL_X4 FILLER_7_242 ();
 FILLCELL_X2 FILLER_7_246 ();
 FILLCELL_X1 FILLER_7_248 ();
 FILLCELL_X4 FILLER_8_1 ();
 FILLCELL_X2 FILLER_8_5 ();
 FILLCELL_X8 FILLER_8_11 ();
 FILLCELL_X4 FILLER_8_19 ();
 FILLCELL_X2 FILLER_8_23 ();
 FILLCELL_X1 FILLER_8_25 ();
 FILLCELL_X32 FILLER_8_53 ();
 FILLCELL_X4 FILLER_8_85 ();
 FILLCELL_X2 FILLER_8_89 ();
 FILLCELL_X1 FILLER_8_91 ();
 FILLCELL_X4 FILLER_8_101 ();
 FILLCELL_X1 FILLER_8_121 ();
 FILLCELL_X2 FILLER_8_133 ();
 FILLCELL_X1 FILLER_8_135 ();
 FILLCELL_X1 FILLER_8_140 ();
 FILLCELL_X2 FILLER_8_144 ();
 FILLCELL_X8 FILLER_8_161 ();
 FILLCELL_X2 FILLER_8_169 ();
 FILLCELL_X1 FILLER_8_171 ();
 FILLCELL_X16 FILLER_8_175 ();
 FILLCELL_X1 FILLER_8_191 ();
 FILLCELL_X2 FILLER_8_197 ();
 FILLCELL_X8 FILLER_8_204 ();
 FILLCELL_X4 FILLER_8_212 ();
 FILLCELL_X1 FILLER_8_216 ();
 FILLCELL_X4 FILLER_8_234 ();
 FILLCELL_X2 FILLER_8_238 ();
 FILLCELL_X1 FILLER_8_240 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_33 ();
 FILLCELL_X1 FILLER_9_37 ();
 FILLCELL_X32 FILLER_9_43 ();
 FILLCELL_X4 FILLER_9_75 ();
 FILLCELL_X2 FILLER_9_79 ();
 FILLCELL_X1 FILLER_9_81 ();
 FILLCELL_X8 FILLER_9_90 ();
 FILLCELL_X1 FILLER_9_98 ();
 FILLCELL_X16 FILLER_9_104 ();
 FILLCELL_X4 FILLER_9_120 ();
 FILLCELL_X2 FILLER_9_124 ();
 FILLCELL_X4 FILLER_9_129 ();
 FILLCELL_X1 FILLER_9_133 ();
 FILLCELL_X1 FILLER_9_137 ();
 FILLCELL_X2 FILLER_9_141 ();
 FILLCELL_X1 FILLER_9_143 ();
 FILLCELL_X4 FILLER_9_147 ();
 FILLCELL_X2 FILLER_9_151 ();
 FILLCELL_X32 FILLER_9_157 ();
 FILLCELL_X1 FILLER_9_189 ();
 FILLCELL_X16 FILLER_9_193 ();
 FILLCELL_X8 FILLER_9_209 ();
 FILLCELL_X2 FILLER_9_217 ();
 FILLCELL_X1 FILLER_9_219 ();
 FILLCELL_X8 FILLER_9_228 ();
 FILLCELL_X4 FILLER_9_236 ();
 FILLCELL_X1 FILLER_9_240 ();
 FILLCELL_X2 FILLER_9_244 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X16 FILLER_10_33 ();
 FILLCELL_X4 FILLER_10_49 ();
 FILLCELL_X2 FILLER_10_53 ();
 FILLCELL_X1 FILLER_10_55 ();
 FILLCELL_X16 FILLER_10_63 ();
 FILLCELL_X8 FILLER_10_79 ();
 FILLCELL_X1 FILLER_10_87 ();
 FILLCELL_X4 FILLER_10_130 ();
 FILLCELL_X2 FILLER_10_134 ();
 FILLCELL_X2 FILLER_10_139 ();
 FILLCELL_X1 FILLER_10_141 ();
 FILLCELL_X1 FILLER_10_151 ();
 FILLCELL_X1 FILLER_10_165 ();
 FILLCELL_X8 FILLER_10_173 ();
 FILLCELL_X2 FILLER_10_181 ();
 FILLCELL_X4 FILLER_10_186 ();
 FILLCELL_X2 FILLER_10_190 ();
 FILLCELL_X16 FILLER_10_217 ();
 FILLCELL_X4 FILLER_10_233 ();
 FILLCELL_X2 FILLER_10_237 ();
 FILLCELL_X1 FILLER_10_239 ();
 FILLCELL_X2 FILLER_10_243 ();
 FILLCELL_X1 FILLER_10_245 ();
 FILLCELL_X4 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_5 ();
 FILLCELL_X32 FILLER_11_14 ();
 FILLCELL_X16 FILLER_11_46 ();
 FILLCELL_X8 FILLER_11_62 ();
 FILLCELL_X2 FILLER_11_77 ();
 FILLCELL_X1 FILLER_11_79 ();
 FILLCELL_X8 FILLER_11_85 ();
 FILLCELL_X4 FILLER_11_93 ();
 FILLCELL_X2 FILLER_11_97 ();
 FILLCELL_X8 FILLER_11_104 ();
 FILLCELL_X4 FILLER_11_112 ();
 FILLCELL_X1 FILLER_11_122 ();
 FILLCELL_X1 FILLER_11_126 ();
 FILLCELL_X1 FILLER_11_131 ();
 FILLCELL_X2 FILLER_11_136 ();
 FILLCELL_X2 FILLER_11_146 ();
 FILLCELL_X2 FILLER_11_152 ();
 FILLCELL_X4 FILLER_11_161 ();
 FILLCELL_X1 FILLER_11_165 ();
 FILLCELL_X32 FILLER_11_177 ();
 FILLCELL_X32 FILLER_11_209 ();
 FILLCELL_X8 FILLER_11_241 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_33 ();
 FILLCELL_X8 FILLER_12_49 ();
 FILLCELL_X4 FILLER_12_57 ();
 FILLCELL_X2 FILLER_12_61 ();
 FILLCELL_X1 FILLER_12_63 ();
 FILLCELL_X8 FILLER_12_84 ();
 FILLCELL_X4 FILLER_12_92 ();
 FILLCELL_X1 FILLER_12_96 ();
 FILLCELL_X1 FILLER_12_107 ();
 FILLCELL_X4 FILLER_12_110 ();
 FILLCELL_X1 FILLER_12_114 ();
 FILLCELL_X16 FILLER_12_130 ();
 FILLCELL_X8 FILLER_12_146 ();
 FILLCELL_X1 FILLER_12_154 ();
 FILLCELL_X4 FILLER_12_158 ();
 FILLCELL_X8 FILLER_12_167 ();
 FILLCELL_X4 FILLER_12_175 ();
 FILLCELL_X8 FILLER_12_182 ();
 FILLCELL_X2 FILLER_12_190 ();
 FILLCELL_X4 FILLER_12_195 ();
 FILLCELL_X16 FILLER_12_203 ();
 FILLCELL_X4 FILLER_12_219 ();
 FILLCELL_X2 FILLER_12_223 ();
 FILLCELL_X2 FILLER_12_229 ();
 FILLCELL_X8 FILLER_12_235 ();
 FILLCELL_X2 FILLER_12_246 ();
 FILLCELL_X1 FILLER_12_248 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X16 FILLER_13_65 ();
 FILLCELL_X2 FILLER_13_81 ();
 FILLCELL_X1 FILLER_13_83 ();
 FILLCELL_X8 FILLER_13_92 ();
 FILLCELL_X4 FILLER_13_100 ();
 FILLCELL_X2 FILLER_13_104 ();
 FILLCELL_X1 FILLER_13_106 ();
 FILLCELL_X16 FILLER_13_117 ();
 FILLCELL_X4 FILLER_13_133 ();
 FILLCELL_X1 FILLER_13_144 ();
 FILLCELL_X2 FILLER_13_149 ();
 FILLCELL_X8 FILLER_13_155 ();
 FILLCELL_X4 FILLER_13_163 ();
 FILLCELL_X2 FILLER_13_167 ();
 FILLCELL_X4 FILLER_13_182 ();
 FILLCELL_X4 FILLER_13_190 ();
 FILLCELL_X2 FILLER_13_194 ();
 FILLCELL_X1 FILLER_13_196 ();
 FILLCELL_X1 FILLER_13_201 ();
 FILLCELL_X2 FILLER_13_219 ();
 FILLCELL_X2 FILLER_13_241 ();
 FILLCELL_X1 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_5 ();
 FILLCELL_X8 FILLER_14_37 ();
 FILLCELL_X2 FILLER_14_45 ();
 FILLCELL_X2 FILLER_14_57 ();
 FILLCELL_X4 FILLER_14_64 ();
 FILLCELL_X2 FILLER_14_68 ();
 FILLCELL_X1 FILLER_14_70 ();
 FILLCELL_X2 FILLER_14_78 ();
 FILLCELL_X1 FILLER_14_80 ();
 FILLCELL_X1 FILLER_14_89 ();
 FILLCELL_X8 FILLER_14_94 ();
 FILLCELL_X2 FILLER_14_102 ();
 FILLCELL_X1 FILLER_14_104 ();
 FILLCELL_X1 FILLER_14_113 ();
 FILLCELL_X1 FILLER_14_118 ();
 FILLCELL_X4 FILLER_14_121 ();
 FILLCELL_X2 FILLER_14_128 ();
 FILLCELL_X1 FILLER_14_130 ();
 FILLCELL_X2 FILLER_14_136 ();
 FILLCELL_X32 FILLER_14_148 ();
 FILLCELL_X1 FILLER_14_180 ();
 FILLCELL_X32 FILLER_14_196 ();
 FILLCELL_X16 FILLER_14_228 ();
 FILLCELL_X4 FILLER_14_244 ();
 FILLCELL_X1 FILLER_14_248 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X8 FILLER_15_33 ();
 FILLCELL_X2 FILLER_15_41 ();
 FILLCELL_X1 FILLER_15_43 ();
 FILLCELL_X4 FILLER_15_54 ();
 FILLCELL_X1 FILLER_15_75 ();
 FILLCELL_X2 FILLER_15_79 ();
 FILLCELL_X1 FILLER_15_81 ();
 FILLCELL_X4 FILLER_15_97 ();
 FILLCELL_X1 FILLER_15_101 ();
 FILLCELL_X2 FILLER_15_110 ();
 FILLCELL_X1 FILLER_15_112 ();
 FILLCELL_X8 FILLER_15_117 ();
 FILLCELL_X4 FILLER_15_125 ();
 FILLCELL_X4 FILLER_15_131 ();
 FILLCELL_X2 FILLER_15_135 ();
 FILLCELL_X1 FILLER_15_137 ();
 FILLCELL_X2 FILLER_15_146 ();
 FILLCELL_X4 FILLER_15_152 ();
 FILLCELL_X2 FILLER_15_156 ();
 FILLCELL_X8 FILLER_15_161 ();
 FILLCELL_X16 FILLER_15_173 ();
 FILLCELL_X2 FILLER_15_189 ();
 FILLCELL_X1 FILLER_15_191 ();
 FILLCELL_X32 FILLER_15_196 ();
 FILLCELL_X16 FILLER_15_228 ();
 FILLCELL_X4 FILLER_15_244 ();
 FILLCELL_X1 FILLER_15_248 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X16 FILLER_16_33 ();
 FILLCELL_X8 FILLER_16_49 ();
 FILLCELL_X4 FILLER_16_57 ();
 FILLCELL_X2 FILLER_16_61 ();
 FILLCELL_X16 FILLER_16_67 ();
 FILLCELL_X8 FILLER_16_83 ();
 FILLCELL_X4 FILLER_16_103 ();
 FILLCELL_X1 FILLER_16_107 ();
 FILLCELL_X8 FILLER_16_115 ();
 FILLCELL_X4 FILLER_16_123 ();
 FILLCELL_X2 FILLER_16_127 ();
 FILLCELL_X8 FILLER_16_133 ();
 FILLCELL_X1 FILLER_16_141 ();
 FILLCELL_X8 FILLER_16_145 ();
 FILLCELL_X4 FILLER_16_153 ();
 FILLCELL_X1 FILLER_16_157 ();
 FILLCELL_X4 FILLER_16_162 ();
 FILLCELL_X1 FILLER_16_166 ();
 FILLCELL_X32 FILLER_16_171 ();
 FILLCELL_X32 FILLER_16_203 ();
 FILLCELL_X8 FILLER_16_235 ();
 FILLCELL_X4 FILLER_16_243 ();
 FILLCELL_X2 FILLER_16_247 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X16 FILLER_17_33 ();
 FILLCELL_X4 FILLER_17_49 ();
 FILLCELL_X1 FILLER_17_53 ();
 FILLCELL_X4 FILLER_17_64 ();
 FILLCELL_X8 FILLER_17_71 ();
 FILLCELL_X2 FILLER_17_79 ();
 FILLCELL_X8 FILLER_17_91 ();
 FILLCELL_X4 FILLER_17_99 ();
 FILLCELL_X2 FILLER_17_103 ();
 FILLCELL_X1 FILLER_17_109 ();
 FILLCELL_X4 FILLER_17_115 ();
 FILLCELL_X1 FILLER_17_126 ();
 FILLCELL_X4 FILLER_17_132 ();
 FILLCELL_X2 FILLER_17_136 ();
 FILLCELL_X1 FILLER_17_138 ();
 FILLCELL_X16 FILLER_17_152 ();
 FILLCELL_X1 FILLER_17_168 ();
 FILLCELL_X4 FILLER_17_172 ();
 FILLCELL_X2 FILLER_17_176 ();
 FILLCELL_X1 FILLER_17_178 ();
 FILLCELL_X2 FILLER_17_187 ();
 FILLCELL_X2 FILLER_17_206 ();
 FILLCELL_X8 FILLER_17_212 ();
 FILLCELL_X2 FILLER_17_237 ();
 FILLCELL_X1 FILLER_17_239 ();
 FILLCELL_X2 FILLER_17_243 ();
 FILLCELL_X1 FILLER_17_245 ();
 FILLCELL_X16 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_17 ();
 FILLCELL_X2 FILLER_18_21 ();
 FILLCELL_X1 FILLER_18_23 ();
 FILLCELL_X16 FILLER_18_28 ();
 FILLCELL_X8 FILLER_18_44 ();
 FILLCELL_X1 FILLER_18_52 ();
 FILLCELL_X16 FILLER_18_66 ();
 FILLCELL_X2 FILLER_18_82 ();
 FILLCELL_X4 FILLER_18_105 ();
 FILLCELL_X1 FILLER_18_109 ();
 FILLCELL_X1 FILLER_18_117 ();
 FILLCELL_X2 FILLER_18_133 ();
 FILLCELL_X4 FILLER_18_147 ();
 FILLCELL_X1 FILLER_18_151 ();
 FILLCELL_X4 FILLER_18_156 ();
 FILLCELL_X1 FILLER_18_160 ();
 FILLCELL_X1 FILLER_18_164 ();
 FILLCELL_X2 FILLER_18_190 ();
 FILLCELL_X2 FILLER_18_196 ();
 FILLCELL_X1 FILLER_18_198 ();
 FILLCELL_X4 FILLER_18_203 ();
 FILLCELL_X8 FILLER_18_228 ();
 FILLCELL_X4 FILLER_18_236 ();
 FILLCELL_X2 FILLER_18_240 ();
 FILLCELL_X1 FILLER_18_242 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X16 FILLER_19_65 ();
 FILLCELL_X4 FILLER_19_81 ();
 FILLCELL_X2 FILLER_19_94 ();
 FILLCELL_X1 FILLER_19_96 ();
 FILLCELL_X16 FILLER_19_101 ();
 FILLCELL_X2 FILLER_19_117 ();
 FILLCELL_X1 FILLER_19_119 ();
 FILLCELL_X4 FILLER_19_123 ();
 FILLCELL_X2 FILLER_19_131 ();
 FILLCELL_X1 FILLER_19_133 ();
 FILLCELL_X1 FILLER_19_137 ();
 FILLCELL_X16 FILLER_19_145 ();
 FILLCELL_X4 FILLER_19_161 ();
 FILLCELL_X2 FILLER_19_165 ();
 FILLCELL_X1 FILLER_19_167 ();
 FILLCELL_X4 FILLER_19_172 ();
 FILLCELL_X2 FILLER_19_176 ();
 FILLCELL_X1 FILLER_19_178 ();
 FILLCELL_X8 FILLER_19_182 ();
 FILLCELL_X4 FILLER_19_190 ();
 FILLCELL_X32 FILLER_19_197 ();
 FILLCELL_X16 FILLER_19_229 ();
 FILLCELL_X4 FILLER_19_245 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X16 FILLER_20_65 ();
 FILLCELL_X8 FILLER_20_81 ();
 FILLCELL_X4 FILLER_20_89 ();
 FILLCELL_X1 FILLER_20_100 ();
 FILLCELL_X2 FILLER_20_105 ();
 FILLCELL_X1 FILLER_20_107 ();
 FILLCELL_X4 FILLER_20_117 ();
 FILLCELL_X2 FILLER_20_121 ();
 FILLCELL_X4 FILLER_20_126 ();
 FILLCELL_X2 FILLER_20_130 ();
 FILLCELL_X1 FILLER_20_132 ();
 FILLCELL_X2 FILLER_20_139 ();
 FILLCELL_X2 FILLER_20_145 ();
 FILLCELL_X8 FILLER_20_153 ();
 FILLCELL_X4 FILLER_20_161 ();
 FILLCELL_X2 FILLER_20_165 ();
 FILLCELL_X2 FILLER_20_170 ();
 FILLCELL_X1 FILLER_20_172 ();
 FILLCELL_X8 FILLER_20_180 ();
 FILLCELL_X4 FILLER_20_188 ();
 FILLCELL_X2 FILLER_20_192 ();
 FILLCELL_X8 FILLER_20_198 ();
 FILLCELL_X2 FILLER_20_206 ();
 FILLCELL_X8 FILLER_20_212 ();
 FILLCELL_X4 FILLER_20_237 ();
 FILLCELL_X2 FILLER_20_241 ();
 FILLCELL_X2 FILLER_20_246 ();
 FILLCELL_X1 FILLER_20_248 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X4 FILLER_21_65 ();
 FILLCELL_X8 FILLER_21_84 ();
 FILLCELL_X1 FILLER_21_92 ();
 FILLCELL_X8 FILLER_21_105 ();
 FILLCELL_X4 FILLER_21_113 ();
 FILLCELL_X4 FILLER_21_123 ();
 FILLCELL_X1 FILLER_21_127 ();
 FILLCELL_X16 FILLER_21_131 ();
 FILLCELL_X4 FILLER_21_147 ();
 FILLCELL_X2 FILLER_21_151 ();
 FILLCELL_X8 FILLER_21_157 ();
 FILLCELL_X2 FILLER_21_165 ();
 FILLCELL_X1 FILLER_21_167 ();
 FILLCELL_X4 FILLER_21_171 ();
 FILLCELL_X8 FILLER_21_183 ();
 FILLCELL_X2 FILLER_21_191 ();
 FILLCELL_X1 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_201 ();
 FILLCELL_X4 FILLER_21_233 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X8 FILLER_22_65 ();
 FILLCELL_X2 FILLER_22_73 ();
 FILLCELL_X1 FILLER_22_75 ();
 FILLCELL_X1 FILLER_22_84 ();
 FILLCELL_X2 FILLER_22_90 ();
 FILLCELL_X1 FILLER_22_103 ();
 FILLCELL_X4 FILLER_22_115 ();
 FILLCELL_X2 FILLER_22_119 ();
 FILLCELL_X8 FILLER_22_138 ();
 FILLCELL_X8 FILLER_22_158 ();
 FILLCELL_X8 FILLER_22_182 ();
 FILLCELL_X1 FILLER_22_190 ();
 FILLCELL_X8 FILLER_22_216 ();
 FILLCELL_X2 FILLER_22_244 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X16 FILLER_23_65 ();
 FILLCELL_X1 FILLER_23_81 ();
 FILLCELL_X4 FILLER_23_86 ();
 FILLCELL_X1 FILLER_23_90 ();
 FILLCELL_X8 FILLER_23_95 ();
 FILLCELL_X2 FILLER_23_103 ();
 FILLCELL_X16 FILLER_23_110 ();
 FILLCELL_X8 FILLER_23_126 ();
 FILLCELL_X8 FILLER_23_138 ();
 FILLCELL_X32 FILLER_23_158 ();
 FILLCELL_X32 FILLER_23_190 ();
 FILLCELL_X16 FILLER_23_222 ();
 FILLCELL_X8 FILLER_23_238 ();
 FILLCELL_X2 FILLER_23_246 ();
 FILLCELL_X1 FILLER_23_248 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X8 FILLER_24_97 ();
 FILLCELL_X4 FILLER_24_105 ();
 FILLCELL_X2 FILLER_24_109 ();
 FILLCELL_X2 FILLER_24_115 ();
 FILLCELL_X16 FILLER_24_120 ();
 FILLCELL_X4 FILLER_24_136 ();
 FILLCELL_X32 FILLER_24_143 ();
 FILLCELL_X2 FILLER_24_175 ();
 FILLCELL_X4 FILLER_24_181 ();
 FILLCELL_X2 FILLER_24_189 ();
 FILLCELL_X1 FILLER_24_191 ();
 FILLCELL_X32 FILLER_24_216 ();
 FILLCELL_X1 FILLER_24_248 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X16 FILLER_25_97 ();
 FILLCELL_X8 FILLER_25_113 ();
 FILLCELL_X4 FILLER_25_121 ();
 FILLCELL_X2 FILLER_25_125 ();
 FILLCELL_X1 FILLER_25_127 ();
 FILLCELL_X8 FILLER_25_131 ();
 FILLCELL_X4 FILLER_25_139 ();
 FILLCELL_X1 FILLER_25_143 ();
 FILLCELL_X32 FILLER_25_147 ();
 FILLCELL_X8 FILLER_25_179 ();
 FILLCELL_X32 FILLER_25_207 ();
 FILLCELL_X8 FILLER_25_239 ();
 FILLCELL_X2 FILLER_25_247 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X8 FILLER_26_97 ();
 FILLCELL_X2 FILLER_26_105 ();
 FILLCELL_X8 FILLER_26_114 ();
 FILLCELL_X2 FILLER_26_122 ();
 FILLCELL_X1 FILLER_26_124 ();
 FILLCELL_X8 FILLER_26_129 ();
 FILLCELL_X2 FILLER_26_141 ();
 FILLCELL_X1 FILLER_26_143 ();
 FILLCELL_X4 FILLER_26_148 ();
 FILLCELL_X2 FILLER_26_152 ();
 FILLCELL_X32 FILLER_26_158 ();
 FILLCELL_X32 FILLER_26_190 ();
 FILLCELL_X2 FILLER_26_222 ();
 FILLCELL_X1 FILLER_26_224 ();
 FILLCELL_X16 FILLER_26_231 ();
 FILLCELL_X2 FILLER_26_247 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X4 FILLER_27_114 ();
 FILLCELL_X2 FILLER_27_118 ();
 FILLCELL_X4 FILLER_27_137 ();
 FILLCELL_X16 FILLER_27_158 ();
 FILLCELL_X2 FILLER_27_174 ();
 FILLCELL_X1 FILLER_27_176 ();
 FILLCELL_X32 FILLER_27_181 ();
 FILLCELL_X32 FILLER_27_213 ();
 FILLCELL_X4 FILLER_27_245 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X8 FILLER_28_161 ();
 FILLCELL_X2 FILLER_28_169 ();
 FILLCELL_X1 FILLER_28_171 ();
 FILLCELL_X32 FILLER_28_189 ();
 FILLCELL_X16 FILLER_28_221 ();
 FILLCELL_X8 FILLER_28_237 ();
 FILLCELL_X4 FILLER_28_245 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X8 FILLER_29_161 ();
 FILLCELL_X4 FILLER_29_169 ();
 FILLCELL_X2 FILLER_29_173 ();
 FILLCELL_X1 FILLER_29_175 ();
 FILLCELL_X32 FILLER_29_179 ();
 FILLCELL_X32 FILLER_29_211 ();
 FILLCELL_X4 FILLER_29_243 ();
 FILLCELL_X2 FILLER_29_247 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X16 FILLER_30_97 ();
 FILLCELL_X4 FILLER_30_113 ();
 FILLCELL_X2 FILLER_30_117 ();
 FILLCELL_X4 FILLER_30_125 ();
 FILLCELL_X2 FILLER_30_129 ();
 FILLCELL_X1 FILLER_30_131 ();
 FILLCELL_X4 FILLER_30_149 ();
 FILLCELL_X2 FILLER_30_153 ();
 FILLCELL_X1 FILLER_30_155 ();
 FILLCELL_X32 FILLER_30_162 ();
 FILLCELL_X32 FILLER_30_194 ();
 FILLCELL_X16 FILLER_30_226 ();
 FILLCELL_X4 FILLER_30_242 ();
 FILLCELL_X2 FILLER_30_246 ();
 FILLCELL_X1 FILLER_30_248 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X8 FILLER_31_97 ();
 FILLCELL_X4 FILLER_31_105 ();
 FILLCELL_X16 FILLER_31_129 ();
 FILLCELL_X2 FILLER_31_145 ();
 FILLCELL_X1 FILLER_31_147 ();
 FILLCELL_X32 FILLER_31_171 ();
 FILLCELL_X32 FILLER_31_203 ();
 FILLCELL_X8 FILLER_31_235 ();
 FILLCELL_X4 FILLER_31_243 ();
 FILLCELL_X2 FILLER_31_247 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X8 FILLER_32_97 ();
 FILLCELL_X4 FILLER_32_105 ();
 FILLCELL_X8 FILLER_32_115 ();
 FILLCELL_X1 FILLER_32_123 ();
 FILLCELL_X8 FILLER_32_127 ();
 FILLCELL_X4 FILLER_32_135 ();
 FILLCELL_X2 FILLER_32_139 ();
 FILLCELL_X16 FILLER_32_144 ();
 FILLCELL_X2 FILLER_32_160 ();
 FILLCELL_X8 FILLER_32_171 ();
 FILLCELL_X4 FILLER_32_179 ();
 FILLCELL_X2 FILLER_32_183 ();
 FILLCELL_X1 FILLER_32_185 ();
 FILLCELL_X32 FILLER_32_189 ();
 FILLCELL_X16 FILLER_32_221 ();
 FILLCELL_X8 FILLER_32_237 ();
 FILLCELL_X4 FILLER_32_245 ();
endmodule
