module toggle_register (clk,
    enable,
    load_en,
    rst_n,
    data_out,
    load_data,
    toggle_mask);
 input clk;
 input enable;
 input load_en;
 input rst_n;
 output [7:0] data_out;
 input [7:0] load_data;
 input [7:0] toggle_mask;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire _37_;
 wire _38_;
 wire _39_;
 wire _40_;
 wire _41_;
 wire _42_;
 wire _43_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 CLKBUF_X3 _44_ (.A(rst_n),
    .Z(_08_));
 INV_X2 _45_ (.A(net9),
    .ZN(_09_));
 BUF_X4 _46_ (.A(_09_),
    .Z(_10_));
 OAI21_X1 _47_ (.A(_08_),
    .B1(net1),
    .B2(_10_),
    .ZN(_11_));
 BUF_X8 _48_ (.A(enable),
    .Z(_12_));
 NAND2_X1 _49_ (.A1(_12_),
    .A2(net10),
    .ZN(_13_));
 XOR2_X1 _50_ (.A(net18),
    .B(_13_),
    .Z(_14_));
 AOI21_X1 _51_ (.A(_11_),
    .B1(_14_),
    .B2(_10_),
    .ZN(_00_));
 OAI21_X1 _52_ (.A(_08_),
    .B1(net2),
    .B2(_10_),
    .ZN(_15_));
 NAND2_X1 _53_ (.A1(_12_),
    .A2(net11),
    .ZN(_16_));
 XOR2_X1 _54_ (.A(net19),
    .B(_16_),
    .Z(_17_));
 AOI21_X1 _55_ (.A(_15_),
    .B1(_17_),
    .B2(_10_),
    .ZN(_01_));
 OAI21_X1 _56_ (.A(_08_),
    .B1(net3),
    .B2(_09_),
    .ZN(_18_));
 NAND2_X1 _57_ (.A1(_12_),
    .A2(net12),
    .ZN(_19_));
 XOR2_X1 _58_ (.A(net20),
    .B(_19_),
    .Z(_20_));
 AOI21_X1 _59_ (.A(_18_),
    .B1(_20_),
    .B2(_10_),
    .ZN(_02_));
 OAI21_X1 _60_ (.A(_08_),
    .B1(net4),
    .B2(_09_),
    .ZN(_21_));
 NAND2_X1 _61_ (.A1(_12_),
    .A2(net13),
    .ZN(_22_));
 XOR2_X1 _62_ (.A(net21),
    .B(_22_),
    .Z(_23_));
 AOI21_X1 _63_ (.A(_21_),
    .B1(_23_),
    .B2(_10_),
    .ZN(_03_));
 OAI21_X1 _64_ (.A(_08_),
    .B1(net5),
    .B2(_09_),
    .ZN(_24_));
 NAND2_X1 _65_ (.A1(_12_),
    .A2(net14),
    .ZN(_25_));
 XOR2_X1 _66_ (.A(net22),
    .B(_25_),
    .Z(_26_));
 AOI21_X1 _67_ (.A(_24_),
    .B1(_26_),
    .B2(_10_),
    .ZN(_04_));
 OAI21_X1 _68_ (.A(_08_),
    .B1(net6),
    .B2(_09_),
    .ZN(_27_));
 NAND2_X1 _69_ (.A1(_12_),
    .A2(net15),
    .ZN(_28_));
 XOR2_X1 _70_ (.A(net23),
    .B(_28_),
    .Z(_29_));
 AOI21_X1 _71_ (.A(_27_),
    .B1(_29_),
    .B2(_10_),
    .ZN(_05_));
 OAI21_X1 _72_ (.A(_08_),
    .B1(net7),
    .B2(_09_),
    .ZN(_30_));
 NAND2_X1 _73_ (.A1(_12_),
    .A2(net16),
    .ZN(_31_));
 XOR2_X1 _74_ (.A(net24),
    .B(_31_),
    .Z(_32_));
 AOI21_X1 _75_ (.A(_30_),
    .B1(_32_),
    .B2(_10_),
    .ZN(_06_));
 OAI21_X1 _76_ (.A(_08_),
    .B1(net8),
    .B2(_09_),
    .ZN(_33_));
 NAND2_X1 _77_ (.A1(_12_),
    .A2(net17),
    .ZN(_34_));
 XOR2_X1 _78_ (.A(net25),
    .B(_34_),
    .Z(_35_));
 AOI21_X1 _79_ (.A(_33_),
    .B1(_35_),
    .B2(_10_),
    .ZN(_07_));
 DFF_X1 \data_out[0]$_SDFFE_PN0P_  (.D(_00_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net18),
    .QN(_43_));
 DFF_X1 \data_out[1]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net19),
    .QN(_42_));
 DFF_X1 \data_out[2]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net20),
    .QN(_41_));
 DFF_X1 \data_out[3]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net21),
    .QN(_40_));
 DFF_X1 \data_out[4]$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net22),
    .QN(_39_));
 DFF_X1 \data_out[5]$_SDFFE_PN0P_  (.D(_05_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net23),
    .QN(_38_));
 DFF_X1 \data_out[6]$_SDFFE_PN0P_  (.D(_06_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net24),
    .QN(_37_));
 DFF_X1 \data_out[7]$_SDFFE_PN0P_  (.D(_07_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net25),
    .QN(_36_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_59 ();
 BUF_X1 input1 (.A(load_data[0]),
    .Z(net1));
 BUF_X1 input2 (.A(load_data[1]),
    .Z(net2));
 BUF_X1 input3 (.A(load_data[2]),
    .Z(net3));
 BUF_X1 input4 (.A(load_data[3]),
    .Z(net4));
 BUF_X1 input5 (.A(load_data[4]),
    .Z(net5));
 BUF_X1 input6 (.A(load_data[5]),
    .Z(net6));
 BUF_X1 input7 (.A(load_data[6]),
    .Z(net7));
 BUF_X1 input8 (.A(load_data[7]),
    .Z(net8));
 BUF_X1 input9 (.A(load_en),
    .Z(net9));
 BUF_X1 input10 (.A(toggle_mask[0]),
    .Z(net10));
 BUF_X1 input11 (.A(toggle_mask[1]),
    .Z(net11));
 BUF_X1 input12 (.A(toggle_mask[2]),
    .Z(net12));
 BUF_X1 input13 (.A(toggle_mask[3]),
    .Z(net13));
 BUF_X1 input14 (.A(toggle_mask[4]),
    .Z(net14));
 BUF_X1 input15 (.A(toggle_mask[5]),
    .Z(net15));
 BUF_X1 input16 (.A(toggle_mask[6]),
    .Z(net16));
 BUF_X1 input17 (.A(toggle_mask[7]),
    .Z(net17));
 BUF_X1 output18 (.A(net18),
    .Z(data_out[0]));
 BUF_X1 output19 (.A(net19),
    .Z(data_out[1]));
 BUF_X1 output20 (.A(net20),
    .Z(data_out[2]));
 BUF_X1 output21 (.A(net21),
    .Z(data_out[3]));
 BUF_X1 output22 (.A(net22),
    .Z(data_out[4]));
 BUF_X1 output23 (.A(net23),
    .Z(data_out[5]));
 BUF_X1 output24 (.A(net24),
    .Z(data_out[6]));
 BUF_X1 output25 (.A(net25),
    .Z(data_out[7]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_73 ();
 FILLCELL_X2 FILLER_0_77 ();
 FILLCELL_X16 FILLER_0_82 ();
 FILLCELL_X8 FILLER_0_98 ();
 FILLCELL_X1 FILLER_0_106 ();
 FILLCELL_X4 FILLER_0_110 ();
 FILLCELL_X1 FILLER_0_117 ();
 FILLCELL_X32 FILLER_0_121 ();
 FILLCELL_X32 FILLER_0_153 ();
 FILLCELL_X32 FILLER_0_185 ();
 FILLCELL_X4 FILLER_0_217 ();
 FILLCELL_X1 FILLER_0_221 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X8 FILLER_1_97 ();
 FILLCELL_X4 FILLER_1_105 ();
 FILLCELL_X2 FILLER_1_109 ();
 FILLCELL_X1 FILLER_1_111 ();
 FILLCELL_X32 FILLER_1_115 ();
 FILLCELL_X32 FILLER_1_147 ();
 FILLCELL_X32 FILLER_1_179 ();
 FILLCELL_X8 FILLER_1_211 ();
 FILLCELL_X2 FILLER_1_219 ();
 FILLCELL_X1 FILLER_1_221 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X16 FILLER_2_193 ();
 FILLCELL_X8 FILLER_2_209 ();
 FILLCELL_X4 FILLER_2_217 ();
 FILLCELL_X1 FILLER_2_221 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X16 FILLER_3_193 ();
 FILLCELL_X8 FILLER_3_209 ();
 FILLCELL_X4 FILLER_3_217 ();
 FILLCELL_X1 FILLER_3_221 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X16 FILLER_4_193 ();
 FILLCELL_X8 FILLER_4_209 ();
 FILLCELL_X4 FILLER_4_217 ();
 FILLCELL_X1 FILLER_4_221 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X16 FILLER_5_193 ();
 FILLCELL_X8 FILLER_5_209 ();
 FILLCELL_X4 FILLER_5_217 ();
 FILLCELL_X1 FILLER_5_221 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X16 FILLER_6_193 ();
 FILLCELL_X8 FILLER_6_209 ();
 FILLCELL_X4 FILLER_6_217 ();
 FILLCELL_X1 FILLER_6_221 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X16 FILLER_7_193 ();
 FILLCELL_X8 FILLER_7_209 ();
 FILLCELL_X4 FILLER_7_217 ();
 FILLCELL_X1 FILLER_7_221 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X8 FILLER_8_97 ();
 FILLCELL_X2 FILLER_8_105 ();
 FILLCELL_X1 FILLER_8_107 ();
 FILLCELL_X32 FILLER_8_113 ();
 FILLCELL_X32 FILLER_8_145 ();
 FILLCELL_X32 FILLER_8_177 ();
 FILLCELL_X8 FILLER_8_209 ();
 FILLCELL_X4 FILLER_8_217 ();
 FILLCELL_X1 FILLER_8_221 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X16 FILLER_9_193 ();
 FILLCELL_X8 FILLER_9_209 ();
 FILLCELL_X4 FILLER_9_217 ();
 FILLCELL_X1 FILLER_9_221 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X2 FILLER_10_9 ();
 FILLCELL_X4 FILLER_10_14 ();
 FILLCELL_X2 FILLER_10_18 ();
 FILLCELL_X16 FILLER_10_26 ();
 FILLCELL_X4 FILLER_10_42 ();
 FILLCELL_X2 FILLER_10_46 ();
 FILLCELL_X1 FILLER_10_48 ();
 FILLCELL_X32 FILLER_10_52 ();
 FILLCELL_X16 FILLER_10_84 ();
 FILLCELL_X8 FILLER_10_100 ();
 FILLCELL_X2 FILLER_10_112 ();
 FILLCELL_X32 FILLER_10_121 ();
 FILLCELL_X32 FILLER_10_153 ();
 FILLCELL_X32 FILLER_10_185 ();
 FILLCELL_X4 FILLER_10_217 ();
 FILLCELL_X1 FILLER_10_221 ();
 FILLCELL_X1 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_19 ();
 FILLCELL_X32 FILLER_11_25 ();
 FILLCELL_X32 FILLER_11_57 ();
 FILLCELL_X16 FILLER_11_89 ();
 FILLCELL_X4 FILLER_11_105 ();
 FILLCELL_X2 FILLER_11_113 ();
 FILLCELL_X32 FILLER_11_121 ();
 FILLCELL_X16 FILLER_11_153 ();
 FILLCELL_X8 FILLER_11_169 ();
 FILLCELL_X1 FILLER_11_177 ();
 FILLCELL_X2 FILLER_11_199 ();
 FILLCELL_X4 FILLER_11_207 ();
 FILLCELL_X2 FILLER_11_217 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_5 ();
 FILLCELL_X4 FILLER_12_9 ();
 FILLCELL_X2 FILLER_12_13 ();
 FILLCELL_X1 FILLER_12_15 ();
 FILLCELL_X32 FILLER_12_20 ();
 FILLCELL_X32 FILLER_12_52 ();
 FILLCELL_X16 FILLER_12_84 ();
 FILLCELL_X2 FILLER_12_100 ();
 FILLCELL_X1 FILLER_12_102 ();
 FILLCELL_X32 FILLER_12_120 ();
 FILLCELL_X32 FILLER_12_152 ();
 FILLCELL_X16 FILLER_12_184 ();
 FILLCELL_X8 FILLER_12_200 ();
 FILLCELL_X1 FILLER_12_208 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X16 FILLER_13_193 ();
 FILLCELL_X8 FILLER_13_209 ();
 FILLCELL_X4 FILLER_13_217 ();
 FILLCELL_X1 FILLER_13_221 ();
 FILLCELL_X1 FILLER_14_4 ();
 FILLCELL_X32 FILLER_14_39 ();
 FILLCELL_X32 FILLER_14_71 ();
 FILLCELL_X32 FILLER_14_103 ();
 FILLCELL_X32 FILLER_14_135 ();
 FILLCELL_X16 FILLER_14_167 ();
 FILLCELL_X2 FILLER_14_183 ();
 FILLCELL_X1 FILLER_14_185 ();
 FILLCELL_X2 FILLER_14_217 ();
 FILLCELL_X2 FILLER_15_1 ();
 FILLCELL_X1 FILLER_15_3 ();
 FILLCELL_X16 FILLER_15_10 ();
 FILLCELL_X4 FILLER_15_26 ();
 FILLCELL_X1 FILLER_15_30 ();
 FILLCELL_X32 FILLER_15_37 ();
 FILLCELL_X2 FILLER_15_69 ();
 FILLCELL_X1 FILLER_15_71 ();
 FILLCELL_X16 FILLER_15_77 ();
 FILLCELL_X2 FILLER_15_93 ();
 FILLCELL_X4 FILLER_15_102 ();
 FILLCELL_X1 FILLER_15_106 ();
 FILLCELL_X16 FILLER_15_112 ();
 FILLCELL_X8 FILLER_15_128 ();
 FILLCELL_X4 FILLER_15_136 ();
 FILLCELL_X32 FILLER_15_145 ();
 FILLCELL_X32 FILLER_15_177 ();
 FILLCELL_X2 FILLER_15_209 ();
 FILLCELL_X2 FILLER_15_217 ();
 FILLCELL_X4 FILLER_16_4 ();
 FILLCELL_X32 FILLER_16_12 ();
 FILLCELL_X32 FILLER_16_44 ();
 FILLCELL_X16 FILLER_16_76 ();
 FILLCELL_X8 FILLER_16_92 ();
 FILLCELL_X2 FILLER_16_100 ();
 FILLCELL_X1 FILLER_16_102 ();
 FILLCELL_X32 FILLER_16_107 ();
 FILLCELL_X32 FILLER_16_139 ();
 FILLCELL_X32 FILLER_16_171 ();
 FILLCELL_X16 FILLER_16_203 ();
 FILLCELL_X2 FILLER_16_219 ();
 FILLCELL_X1 FILLER_16_221 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_9 ();
 FILLCELL_X1 FILLER_17_13 ();
 FILLCELL_X32 FILLER_17_18 ();
 FILLCELL_X32 FILLER_17_50 ();
 FILLCELL_X16 FILLER_17_82 ();
 FILLCELL_X4 FILLER_17_98 ();
 FILLCELL_X32 FILLER_17_106 ();
 FILLCELL_X4 FILLER_17_138 ();
 FILLCELL_X16 FILLER_17_146 ();
 FILLCELL_X8 FILLER_17_162 ();
 FILLCELL_X4 FILLER_17_170 ();
 FILLCELL_X2 FILLER_17_174 ();
 FILLCELL_X1 FILLER_17_176 ();
 FILLCELL_X2 FILLER_17_198 ();
 FILLCELL_X1 FILLER_17_200 ();
 FILLCELL_X2 FILLER_17_207 ();
 FILLCELL_X4 FILLER_17_215 ();
 FILLCELL_X1 FILLER_18_1 ();
 FILLCELL_X8 FILLER_18_5 ();
 FILLCELL_X16 FILLER_18_36 ();
 FILLCELL_X8 FILLER_18_52 ();
 FILLCELL_X4 FILLER_18_60 ();
 FILLCELL_X16 FILLER_18_67 ();
 FILLCELL_X8 FILLER_18_83 ();
 FILLCELL_X4 FILLER_18_91 ();
 FILLCELL_X2 FILLER_18_95 ();
 FILLCELL_X32 FILLER_18_114 ();
 FILLCELL_X32 FILLER_18_146 ();
 FILLCELL_X32 FILLER_18_178 ();
 FILLCELL_X8 FILLER_18_210 ();
 FILLCELL_X4 FILLER_18_218 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X8 FILLER_19_97 ();
 FILLCELL_X4 FILLER_19_105 ();
 FILLCELL_X1 FILLER_19_109 ();
 FILLCELL_X32 FILLER_19_119 ();
 FILLCELL_X32 FILLER_19_151 ();
 FILLCELL_X32 FILLER_19_183 ();
 FILLCELL_X4 FILLER_19_215 ();
 FILLCELL_X2 FILLER_19_219 ();
 FILLCELL_X1 FILLER_19_221 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X16 FILLER_20_193 ();
 FILLCELL_X8 FILLER_20_209 ();
 FILLCELL_X4 FILLER_20_217 ();
 FILLCELL_X1 FILLER_20_221 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X16 FILLER_21_193 ();
 FILLCELL_X8 FILLER_21_209 ();
 FILLCELL_X4 FILLER_21_217 ();
 FILLCELL_X1 FILLER_21_221 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X16 FILLER_22_193 ();
 FILLCELL_X8 FILLER_22_209 ();
 FILLCELL_X4 FILLER_22_217 ();
 FILLCELL_X1 FILLER_22_221 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X16 FILLER_23_193 ();
 FILLCELL_X8 FILLER_23_209 ();
 FILLCELL_X4 FILLER_23_217 ();
 FILLCELL_X1 FILLER_23_221 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X16 FILLER_24_193 ();
 FILLCELL_X8 FILLER_24_209 ();
 FILLCELL_X4 FILLER_24_217 ();
 FILLCELL_X1 FILLER_24_221 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X16 FILLER_25_193 ();
 FILLCELL_X8 FILLER_25_209 ();
 FILLCELL_X4 FILLER_25_217 ();
 FILLCELL_X1 FILLER_25_221 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X16 FILLER_26_193 ();
 FILLCELL_X8 FILLER_26_209 ();
 FILLCELL_X4 FILLER_26_217 ();
 FILLCELL_X1 FILLER_26_221 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X16 FILLER_27_193 ();
 FILLCELL_X8 FILLER_27_209 ();
 FILLCELL_X4 FILLER_27_217 ();
 FILLCELL_X1 FILLER_27_221 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X16 FILLER_28_193 ();
 FILLCELL_X8 FILLER_28_209 ();
 FILLCELL_X4 FILLER_28_217 ();
 FILLCELL_X1 FILLER_28_221 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X16 FILLER_29_33 ();
 FILLCELL_X8 FILLER_29_49 ();
 FILLCELL_X4 FILLER_29_57 ();
 FILLCELL_X2 FILLER_29_61 ();
 FILLCELL_X32 FILLER_29_66 ();
 FILLCELL_X4 FILLER_29_98 ();
 FILLCELL_X2 FILLER_29_102 ();
 FILLCELL_X4 FILLER_29_107 ();
 FILLCELL_X1 FILLER_29_114 ();
 FILLCELL_X4 FILLER_29_118 ();
 FILLCELL_X2 FILLER_29_122 ();
 FILLCELL_X32 FILLER_29_127 ();
 FILLCELL_X32 FILLER_29_159 ();
 FILLCELL_X16 FILLER_29_191 ();
 FILLCELL_X8 FILLER_29_207 ();
 FILLCELL_X4 FILLER_29_215 ();
 FILLCELL_X2 FILLER_29_219 ();
 FILLCELL_X1 FILLER_29_221 ();
endmodule
