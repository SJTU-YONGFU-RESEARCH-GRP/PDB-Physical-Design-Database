module alu (clk,
    overflow_flag,
    rst_n,
    zero_flag,
    a,
    b,
    op_code,
    result);
 input clk;
 output overflow_flag;
 input rst_n;
 output zero_flag;
 input [7:0] a;
 input [7:0] b;
 input [2:0] op_code;
 output [7:0] result;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net30;

 sky130_fd_sc_hd__inv_1 _305_ (.A(_270_),
    .Y(_210_));
 sky130_fd_sc_hd__clkbuf_2 _306_ (.A(_269_),
    .X(_211_));
 sky130_fd_sc_hd__nand2b_1 _307_ (.A_N(_211_),
    .B(_262_),
    .Y(_212_));
 sky130_fd_sc_hd__buf_2 _308_ (.A(_277_),
    .X(_213_));
 sky130_fd_sc_hd__a21oi_1 _309_ (.A1(_210_),
    .A2(_212_),
    .B1(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__clkbuf_2 _310_ (.A(_261_),
    .X(_215_));
 sky130_fd_sc_hd__or3_1 _311_ (.A(_215_),
    .B(_211_),
    .C(_213_),
    .X(_216_));
 sky130_fd_sc_hd__o21ba_1 _312_ (.A1(_243_),
    .A2(_240_),
    .B1_N(_254_),
    .X(_217_));
 sky130_fd_sc_hd__nor2_1 _313_ (.A(_216_),
    .B(_217_),
    .Y(_218_));
 sky130_fd_sc_hd__or3_1 _314_ (.A(_278_),
    .B(_286_),
    .C(_294_),
    .X(_219_));
 sky130_fd_sc_hd__nor2b_1 _315_ (.A(_286_),
    .B_N(_285_),
    .Y(_220_));
 sky130_fd_sc_hd__o21bai_1 _316_ (.A1(_293_),
    .A2(_220_),
    .B1_N(_294_),
    .Y(_221_));
 sky130_fd_sc_hd__o31a_1 _317_ (.A1(_214_),
    .A2(_218_),
    .A3(_219_),
    .B1(_221_),
    .X(_222_));
 sky130_fd_sc_hd__xnor2_1 _318_ (.A(_301_),
    .B(_222_),
    .Y(_223_));
 sky130_fd_sc_hd__inv_1 _319_ (.A(_285_),
    .Y(_224_));
 sky130_fd_sc_hd__nor3_1 _320_ (.A(_278_),
    .B(_214_),
    .C(_218_),
    .Y(_225_));
 sky130_fd_sc_hd__xnor2_1 _321_ (.A(_224_),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__inv_1 _322_ (.A(_211_),
    .Y(_227_));
 sky130_fd_sc_hd__o21bai_1 _323_ (.A1(_215_),
    .A2(_241_),
    .B1_N(_262_),
    .Y(_001_));
 sky130_fd_sc_hd__a21oi_1 _324_ (.A1(_227_),
    .A2(_001_),
    .B1(_270_),
    .Y(_002_));
 sky130_fd_sc_hd__xnor2_1 _325_ (.A(_213_),
    .B(_002_),
    .Y(_003_));
 sky130_fd_sc_hd__nor2_1 _326_ (.A(_215_),
    .B(_217_),
    .Y(_004_));
 sky130_fd_sc_hd__nor2_1 _327_ (.A(_262_),
    .B(_004_),
    .Y(_005_));
 sky130_fd_sc_hd__xnor2_1 _328_ (.A(_211_),
    .B(_005_),
    .Y(_006_));
 sky130_fd_sc_hd__inv_1 _329_ (.A(_242_),
    .Y(_007_));
 sky130_fd_sc_hd__buf_2 _330_ (.A(net19),
    .X(_008_));
 sky130_fd_sc_hd__buf_2 _331_ (.A(op_code[1]),
    .X(_009_));
 sky130_fd_sc_hd__clkinvlp_4 _332_ (.A(net18),
    .Y(_010_));
 sky130_fd_sc_hd__or3_1 _333_ (.A(_008_),
    .B(_009_),
    .C(_010_),
    .X(_011_));
 sky130_fd_sc_hd__xor2_1 _334_ (.A(_215_),
    .B(_241_),
    .X(_012_));
 sky130_fd_sc_hd__nor4_1 _335_ (.A(_247_),
    .B(_007_),
    .C(_011_),
    .D(_012_),
    .Y(_013_));
 sky130_fd_sc_hd__nand4b_1 _336_ (.A_N(_226_),
    .B(_003_),
    .C(_006_),
    .D(_013_),
    .Y(_014_));
 sky130_fd_sc_hd__a21oi_1 _337_ (.A1(_278_),
    .A2(_224_),
    .B1(_286_),
    .Y(_015_));
 sky130_fd_sc_hd__o31ai_1 _338_ (.A1(_213_),
    .A2(_285_),
    .A3(_002_),
    .B1(_015_),
    .Y(_016_));
 sky130_fd_sc_hd__xnor2_1 _339_ (.A(_293_),
    .B(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__buf_2 _340_ (.A(net12),
    .X(_018_));
 sky130_fd_sc_hd__buf_2 _341_ (.A(_018_),
    .X(_019_));
 sky130_fd_sc_hd__clkbuf_4 _342_ (.A(net11),
    .X(_020_));
 sky130_fd_sc_hd__buf_2 _343_ (.A(_020_),
    .X(_021_));
 sky130_fd_sc_hd__buf_6 _344_ (.A(net10),
    .X(_022_));
 sky130_fd_sc_hd__buf_6 _345_ (.A(_022_),
    .X(_023_));
 sky130_fd_sc_hd__inv_1 _346_ (.A(net6),
    .Y(_274_));
 sky130_fd_sc_hd__clkbuf_4 _347_ (.A(_023_),
    .X(_024_));
 sky130_fd_sc_hd__nand2_1 _348_ (.A(_024_),
    .B(net5),
    .Y(_025_));
 sky130_fd_sc_hd__o21ai_2 _349_ (.A1(_023_),
    .A2(_274_),
    .B1(_025_),
    .Y(_026_));
 sky130_fd_sc_hd__inv_1 _350_ (.A(net7),
    .Y(_282_));
 sky130_fd_sc_hd__nor2_1 _351_ (.A(_024_),
    .B(net8),
    .Y(_027_));
 sky130_fd_sc_hd__a211oi_1 _352_ (.A1(_024_),
    .A2(_282_),
    .B1(_027_),
    .C1(_020_),
    .Y(_028_));
 sky130_fd_sc_hd__nor3b_1 _353_ (.A(net2),
    .B(net4),
    .C_N(_023_),
    .Y(_029_));
 sky130_fd_sc_hd__nor3_1 _354_ (.A(net3),
    .B(_024_),
    .C(net5),
    .Y(_030_));
 sky130_fd_sc_hd__a21oi_1 _355_ (.A1(net3),
    .A2(_024_),
    .B1(net4),
    .Y(_031_));
 sky130_fd_sc_hd__o22ai_1 _356_ (.A1(_029_),
    .A2(_030_),
    .B1(_031_),
    .B2(_021_),
    .Y(_032_));
 sky130_fd_sc_hd__a2111oi_1 _357_ (.A1(_021_),
    .A2(_026_),
    .B1(_028_),
    .C1(_032_),
    .D1(_249_),
    .Y(_033_));
 sky130_fd_sc_hd__nor2_1 _358_ (.A(_020_),
    .B(_018_),
    .Y(_034_));
 sky130_fd_sc_hd__mux2i_4 _359_ (.A0(net4),
    .A1(net3),
    .S(_024_),
    .Y(_035_));
 sky130_fd_sc_hd__nand2b_2 _360_ (.A_N(_018_),
    .B(_020_),
    .Y(_036_));
 sky130_fd_sc_hd__and3b_1 _361_ (.A_N(_009_),
    .B(net18),
    .C(net19),
    .X(_037_));
 sky130_fd_sc_hd__buf_2 _362_ (.A(_037_),
    .X(_038_));
 sky130_fd_sc_hd__nand2_1 _363_ (.A(_249_),
    .B(_019_),
    .Y(_039_));
 sky130_fd_sc_hd__o211ai_1 _364_ (.A1(_035_),
    .A2(_036_),
    .B1(_038_),
    .C1(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__clkinv_2 _365_ (.A(_018_),
    .Y(_259_));
 sky130_fd_sc_hd__nor3_1 _366_ (.A(_021_),
    .B(_259_),
    .C(_035_),
    .Y(_041_));
 sky130_fd_sc_hd__a211oi_1 _367_ (.A1(_026_),
    .A2(_034_),
    .B1(_040_),
    .C1(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__mux4_1 _368_ (.A0(net7),
    .A1(net6),
    .A2(net3),
    .A3(net2),
    .S0(_023_),
    .S1(_018_),
    .X(_043_));
 sky130_fd_sc_hd__inv_1 _369_ (.A(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__mux2i_4 _370_ (.A0(net5),
    .A1(net4),
    .S(_024_),
    .Y(_045_));
 sky130_fd_sc_hd__nor2b_1 _371_ (.A(_023_),
    .B_N(net9),
    .Y(_046_));
 sky130_fd_sc_hd__a211oi_1 _372_ (.A1(_024_),
    .A2(net8),
    .B1(_046_),
    .C1(_018_),
    .Y(_047_));
 sky130_fd_sc_hd__a211o_1 _373_ (.A1(_019_),
    .A2(_045_),
    .B1(_047_),
    .C1(_021_),
    .X(_048_));
 sky130_fd_sc_hd__o2111ai_1 _374_ (.A1(_019_),
    .A2(_033_),
    .B1(_042_),
    .C1(_044_),
    .D1(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__mux2i_1 _375_ (.A0(net8),
    .A1(net9),
    .S(_022_),
    .Y(_050_));
 sky130_fd_sc_hd__mux2i_4 _376_ (.A0(net6),
    .A1(net7),
    .S(_022_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _377_ (.A(_020_),
    .Y(_252_));
 sky130_fd_sc_hd__mux2i_2 _378_ (.A0(_050_),
    .A1(_051_),
    .S(_252_),
    .Y(_052_));
 sky130_fd_sc_hd__nand3b_2 _379_ (.A_N(net18),
    .B(_009_),
    .C(net19),
    .Y(_053_));
 sky130_fd_sc_hd__nor2b_1 _380_ (.A(_022_),
    .B_N(net8),
    .Y(_054_));
 sky130_fd_sc_hd__o21ai_0 _381_ (.A1(net9),
    .A2(_054_),
    .B1(_034_),
    .Y(_055_));
 sky130_fd_sc_hd__nand2b_1 _382_ (.A_N(_022_),
    .B(net9),
    .Y(_056_));
 sky130_fd_sc_hd__mux2i_1 _383_ (.A0(net7),
    .A1(net8),
    .S(_022_),
    .Y(_057_));
 sky130_fd_sc_hd__mux2_1 _384_ (.A0(_056_),
    .A1(_057_),
    .S(_252_),
    .X(_058_));
 sky130_fd_sc_hd__nand4bb_1 _385_ (.A_N(_052_),
    .B_N(_053_),
    .C(_055_),
    .D(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__nor2_1 _386_ (.A(_259_),
    .B(_046_),
    .Y(_060_));
 sky130_fd_sc_hd__mux2_1 _387_ (.A0(net5),
    .A1(net6),
    .S(_022_),
    .X(_061_));
 sky130_fd_sc_hd__nor2_1 _388_ (.A(_018_),
    .B(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__o32ai_1 _389_ (.A1(_020_),
    .A2(_060_),
    .A3(_062_),
    .B1(_036_),
    .B2(_057_),
    .Y(_063_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(net4),
    .A1(net5),
    .S(_023_),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(net2),
    .A1(net3),
    .S(_023_),
    .X(_065_));
 sky130_fd_sc_hd__mux2i_2 _392_ (.A0(_064_),
    .A1(_065_),
    .S(_252_),
    .Y(_066_));
 sky130_fd_sc_hd__nand2_1 _393_ (.A(_020_),
    .B(_061_),
    .Y(_067_));
 sky130_fd_sc_hd__inv_1 _394_ (.A(net4),
    .Y(_258_));
 sky130_fd_sc_hd__nor2_1 _395_ (.A(net3),
    .B(_023_),
    .Y(_068_));
 sky130_fd_sc_hd__a211o_1 _396_ (.A1(_023_),
    .A2(_258_),
    .B1(_068_),
    .C1(_020_),
    .X(_069_));
 sky130_fd_sc_hd__a31oi_1 _397_ (.A1(_066_),
    .A2(_067_),
    .A3(_069_),
    .B1(_018_),
    .Y(_070_));
 sky130_fd_sc_hd__nor2_1 _398_ (.A(_018_),
    .B(_064_),
    .Y(_071_));
 sky130_fd_sc_hd__mux2_1 _399_ (.A0(net8),
    .A1(net9),
    .S(_023_),
    .X(_072_));
 sky130_fd_sc_hd__nor2_1 _400_ (.A(_259_),
    .B(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__o32ai_1 _401_ (.A1(_020_),
    .A2(_071_),
    .A3(_073_),
    .B1(_036_),
    .B2(_051_),
    .Y(_074_));
 sky130_fd_sc_hd__or4_1 _402_ (.A(_059_),
    .B(_063_),
    .C(_070_),
    .D(_074_),
    .X(_075_));
 sky130_fd_sc_hd__buf_2 _403_ (.A(_008_),
    .X(_076_));
 sky130_fd_sc_hd__buf_2 _404_ (.A(net18),
    .X(_077_));
 sky130_fd_sc_hd__nand2_1 _405_ (.A(_009_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__inv_1 _406_ (.A(_009_),
    .Y(_079_));
 sky130_fd_sc_hd__nand2_1 _407_ (.A(_079_),
    .B(_010_),
    .Y(_080_));
 sky130_fd_sc_hd__or4_1 _408_ (.A(_243_),
    .B(_285_),
    .C(_293_),
    .D(_301_),
    .X(_081_));
 sky130_fd_sc_hd__nor3_1 _409_ (.A(_247_),
    .B(_216_),
    .C(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__mux2i_1 _410_ (.A0(_078_),
    .A1(_080_),
    .S(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__nand4_1 _411_ (.A(_253_),
    .B(_260_),
    .C(_268_),
    .D(_276_),
    .Y(_084_));
 sky130_fd_sc_hd__nor2b_1 _412_ (.A(_008_),
    .B_N(_009_),
    .Y(_085_));
 sky130_fd_sc_hd__nand2_1 _413_ (.A(_077_),
    .B(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__nand4_1 _414_ (.A(_246_),
    .B(_284_),
    .C(_292_),
    .D(_300_),
    .Y(_087_));
 sky130_fd_sc_hd__nor4_1 _415_ (.A(_272_),
    .B(_280_),
    .C(_288_),
    .D(_296_),
    .Y(_088_));
 sky130_fd_sc_hd__nor3_1 _416_ (.A(_264_),
    .B(_236_),
    .C(_302_),
    .Y(_089_));
 sky130_fd_sc_hd__nor2_1 _417_ (.A(_077_),
    .B(_256_),
    .Y(_090_));
 sky130_fd_sc_hd__nand4_1 _418_ (.A(_088_),
    .B(_085_),
    .C(_089_),
    .D(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__o31ai_1 _419_ (.A1(_084_),
    .A2(_086_),
    .A3(_087_),
    .B1(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__a21oi_1 _420_ (.A1(_076_),
    .A2(_083_),
    .B1(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__and3_1 _421_ (.A(_049_),
    .B(_075_),
    .C(_093_),
    .X(_094_));
 sky130_fd_sc_hd__and3_1 _422_ (.A(_237_),
    .B(_215_),
    .C(_211_),
    .X(_095_));
 sky130_fd_sc_hd__a21o_1 _423_ (.A1(_264_),
    .A2(_211_),
    .B1(_272_),
    .X(_096_));
 sky130_fd_sc_hd__o21ai_1 _424_ (.A1(_095_),
    .A2(_096_),
    .B1(_213_),
    .Y(_097_));
 sky130_fd_sc_hd__nor2_1 _425_ (.A(_280_),
    .B(_288_),
    .Y(_098_));
 sky130_fd_sc_hd__o21ai_0 _426_ (.A1(_288_),
    .A2(_285_),
    .B1(_293_),
    .Y(_099_));
 sky130_fd_sc_hd__a21o_1 _427_ (.A1(_097_),
    .A2(_098_),
    .B1(_099_),
    .X(_100_));
 sky130_fd_sc_hd__nand3b_1 _428_ (.A_N(_293_),
    .B(_097_),
    .C(_098_),
    .Y(_101_));
 sky130_fd_sc_hd__o311ai_2 _429_ (.A1(_288_),
    .A2(_285_),
    .A3(_293_),
    .B1(_100_),
    .C1(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__inv_1 _430_ (.A(_301_),
    .Y(_103_));
 sky130_fd_sc_hd__nor3_1 _431_ (.A(_280_),
    .B(_288_),
    .C(_213_),
    .Y(_104_));
 sky130_fd_sc_hd__inv_1 _432_ (.A(_296_),
    .Y(_105_));
 sky130_fd_sc_hd__o21ai_0 _433_ (.A1(_099_),
    .A2(_104_),
    .B1(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__a211oi_1 _434_ (.A1(_236_),
    .A2(_243_),
    .B1(_256_),
    .C1(_264_),
    .Y(_107_));
 sky130_fd_sc_hd__o21ai_0 _435_ (.A1(_215_),
    .A2(_264_),
    .B1(_211_),
    .Y(_108_));
 sky130_fd_sc_hd__o21ai_0 _436_ (.A1(_107_),
    .A2(_108_),
    .B1(_088_),
    .Y(_109_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(_106_),
    .B(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__xnor2_1 _438_ (.A(_103_),
    .B(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__nor3_2 _439_ (.A(_008_),
    .B(_009_),
    .C(net18),
    .Y(_112_));
 sky130_fd_sc_hd__xnor2_1 _440_ (.A(_237_),
    .B(_215_),
    .Y(_113_));
 sky130_fd_sc_hd__nand2_1 _441_ (.A(_112_),
    .B(_113_),
    .Y(_114_));
 sky130_fd_sc_hd__or3_1 _442_ (.A(_238_),
    .B(_247_),
    .C(_114_),
    .X(_115_));
 sky130_fd_sc_hd__nor2_1 _443_ (.A(_215_),
    .B(_264_),
    .Y(_116_));
 sky130_fd_sc_hd__nor2_1 _444_ (.A(_107_),
    .B(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__xnor2_1 _445_ (.A(_227_),
    .B(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__or2_0 _446_ (.A(_095_),
    .B(_096_),
    .X(_119_));
 sky130_fd_sc_hd__xor2_1 _447_ (.A(_213_),
    .B(_119_),
    .X(_120_));
 sky130_fd_sc_hd__nor3_1 _448_ (.A(_115_),
    .B(_118_),
    .C(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__inv_1 _449_ (.A(_272_),
    .Y(_122_));
 sky130_fd_sc_hd__o21ai_0 _450_ (.A1(_107_),
    .A2(_108_),
    .B1(_122_),
    .Y(_123_));
 sky130_fd_sc_hd__a21oi_1 _451_ (.A1(_213_),
    .A2(_123_),
    .B1(_280_),
    .Y(_124_));
 sky130_fd_sc_hd__xnor2_1 _452_ (.A(_224_),
    .B(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__nand4_1 _453_ (.A(_102_),
    .B(_111_),
    .C(_121_),
    .D(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__o311ai_0 _454_ (.A1(_223_),
    .A2(_014_),
    .A3(_017_),
    .B1(_094_),
    .C1(_126_),
    .Y(_000_));
 sky130_fd_sc_hd__buf_2 _455_ (.A(_079_),
    .X(_127_));
 sky130_fd_sc_hd__nor2_1 _456_ (.A(_077_),
    .B(_236_),
    .Y(_128_));
 sky130_fd_sc_hd__a21oi_1 _457_ (.A1(_077_),
    .A2(_246_),
    .B1(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__buf_2 _458_ (.A(_009_),
    .X(_130_));
 sky130_fd_sc_hd__mux2i_1 _459_ (.A0(_247_),
    .A1(_129_),
    .S(_130_),
    .Y(_131_));
 sky130_fd_sc_hd__nor2_1 _460_ (.A(_076_),
    .B(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__nor2_1 _461_ (.A(_019_),
    .B(_066_),
    .Y(_133_));
 sky130_fd_sc_hd__a21oi_1 _462_ (.A1(_019_),
    .A2(_052_),
    .B1(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__and3_1 _463_ (.A(_127_),
    .B(_249_),
    .C(_034_),
    .X(_135_));
 sky130_fd_sc_hd__a21oi_1 _464_ (.A1(_130_),
    .A2(_082_),
    .B1(_135_),
    .Y(_136_));
 sky130_fd_sc_hd__nand2_1 _465_ (.A(_076_),
    .B(_077_),
    .Y(_137_));
 sky130_fd_sc_hd__o22ai_1 _466_ (.A1(_053_),
    .A2(_134_),
    .B1(_136_),
    .B2(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__a311o_1 _467_ (.A1(_127_),
    .A2(_010_),
    .A3(_247_),
    .B1(_132_),
    .C1(_138_),
    .X(_228_));
 sky130_fd_sc_hd__inv_1 _468_ (.A(net2),
    .Y(_244_));
 sky130_fd_sc_hd__a21oi_1 _469_ (.A1(_244_),
    .A2(_024_),
    .B1(_068_),
    .Y(_139_));
 sky130_fd_sc_hd__nand3_1 _470_ (.A(_034_),
    .B(_139_),
    .C(_038_),
    .Y(_140_));
 sky130_fd_sc_hd__buf_2 _471_ (.A(_077_),
    .X(_141_));
 sky130_fd_sc_hd__a21oi_1 _472_ (.A1(_141_),
    .A2(_253_),
    .B1(_090_),
    .Y(_142_));
 sky130_fd_sc_hd__a21oi_1 _473_ (.A1(_141_),
    .A2(_242_),
    .B1(_076_),
    .Y(_143_));
 sky130_fd_sc_hd__a21oi_1 _474_ (.A1(_010_),
    .A2(_243_),
    .B1(_143_),
    .Y(_144_));
 sky130_fd_sc_hd__nor2_1 _475_ (.A(_130_),
    .B(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__a21oi_1 _476_ (.A1(_085_),
    .A2(_142_),
    .B1(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__and3_1 _477_ (.A(_259_),
    .B(_067_),
    .C(_069_),
    .X(_147_));
 sky130_fd_sc_hd__a211o_1 _478_ (.A1(_019_),
    .A2(_058_),
    .B1(_147_),
    .C1(_053_),
    .X(_148_));
 sky130_fd_sc_hd__or3_2 _479_ (.A(_008_),
    .B(_009_),
    .C(_077_),
    .X(_149_));
 sky130_fd_sc_hd__nor2_1 _480_ (.A(_238_),
    .B(_149_),
    .Y(_150_));
 sky130_fd_sc_hd__a31oi_1 _481_ (.A1(_140_),
    .A2(_146_),
    .A3(_148_),
    .B1(_150_),
    .Y(_229_));
 sky130_fd_sc_hd__nand2_1 _482_ (.A(_141_),
    .B(_260_),
    .Y(_151_));
 sky130_fd_sc_hd__o211ai_1 _483_ (.A1(_141_),
    .A2(_264_),
    .B1(_151_),
    .C1(_130_),
    .Y(_152_));
 sky130_fd_sc_hd__nand3_1 _484_ (.A(_127_),
    .B(_141_),
    .C(_012_),
    .Y(_153_));
 sky130_fd_sc_hd__a21oi_1 _485_ (.A1(_152_),
    .A2(_153_),
    .B1(_076_),
    .Y(_154_));
 sky130_fd_sc_hd__nand2b_1 _486_ (.A_N(_215_),
    .B(_008_),
    .Y(_155_));
 sky130_fd_sc_hd__nor2b_1 _487_ (.A(_249_),
    .B_N(_020_),
    .Y(_156_));
 sky130_fd_sc_hd__a21o_1 _488_ (.A1(_252_),
    .A2(_035_),
    .B1(_156_),
    .X(_157_));
 sky130_fd_sc_hd__nor3_1 _489_ (.A(_019_),
    .B(_137_),
    .C(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__a21oi_1 _490_ (.A1(_010_),
    .A2(_155_),
    .B1(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__nand2b_1 _491_ (.A_N(_053_),
    .B(_074_),
    .Y(_160_));
 sky130_fd_sc_hd__o21ai_0 _492_ (.A1(_130_),
    .A2(_159_),
    .B1(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__o21a_1 _493_ (.A1(_154_),
    .A2(_161_),
    .B1(_114_),
    .X(_230_));
 sky130_fd_sc_hd__nor2b_1 _494_ (.A(_053_),
    .B_N(_063_),
    .Y(_162_));
 sky130_fd_sc_hd__nor2_1 _495_ (.A(_021_),
    .B(_045_),
    .Y(_163_));
 sky130_fd_sc_hd__a21oi_1 _496_ (.A1(_021_),
    .A2(_139_),
    .B1(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__nand2_1 _497_ (.A(_259_),
    .B(_038_),
    .Y(_165_));
 sky130_fd_sc_hd__a21oi_1 _498_ (.A1(_009_),
    .A2(_122_),
    .B1(_008_),
    .Y(_166_));
 sky130_fd_sc_hd__a21oi_1 _499_ (.A1(_127_),
    .A2(_211_),
    .B1(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__o22a_1 _500_ (.A1(_268_),
    .A2(_086_),
    .B1(_167_),
    .B2(_141_),
    .X(_168_));
 sky130_fd_sc_hd__o221ai_1 _501_ (.A1(_006_),
    .A2(_011_),
    .B1(_164_),
    .B2(_165_),
    .C1(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__o22a_1 _502_ (.A1(_149_),
    .A2(_118_),
    .B1(_162_),
    .B2(_169_),
    .X(_231_));
 sky130_fd_sc_hd__a21boi_0 _503_ (.A1(_259_),
    .A2(_026_),
    .B1_N(_039_),
    .Y(_170_));
 sky130_fd_sc_hd__o22ai_1 _504_ (.A1(_035_),
    .A2(_036_),
    .B1(_170_),
    .B2(_021_),
    .Y(_171_));
 sky130_fd_sc_hd__inv_1 _505_ (.A(_280_),
    .Y(_172_));
 sky130_fd_sc_hd__a21oi_1 _506_ (.A1(_130_),
    .A2(_172_),
    .B1(_008_),
    .Y(_173_));
 sky130_fd_sc_hd__a21oi_1 _507_ (.A1(_127_),
    .A2(_213_),
    .B1(_173_),
    .Y(_174_));
 sky130_fd_sc_hd__nor2_1 _508_ (.A(_019_),
    .B(_053_),
    .Y(_175_));
 sky130_fd_sc_hd__nand2_1 _509_ (.A(_052_),
    .B(_175_),
    .Y(_176_));
 sky130_fd_sc_hd__o221ai_1 _510_ (.A1(_276_),
    .A2(_086_),
    .B1(_174_),
    .B2(_141_),
    .C1(_176_),
    .Y(_177_));
 sky130_fd_sc_hd__nor2_1 _511_ (.A(_003_),
    .B(_011_),
    .Y(_178_));
 sky130_fd_sc_hd__a211oi_1 _512_ (.A1(_038_),
    .A2(_171_),
    .B1(_177_),
    .C1(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__nor2_1 _513_ (.A(_149_),
    .B(_120_),
    .Y(_180_));
 sky130_fd_sc_hd__nor2_1 _514_ (.A(_179_),
    .B(_180_),
    .Y(_232_));
 sky130_fd_sc_hd__nor3_2 _515_ (.A(_076_),
    .B(_130_),
    .C(_010_),
    .Y(_181_));
 sky130_fd_sc_hd__o22ai_2 _516_ (.A1(_021_),
    .A2(_044_),
    .B1(_036_),
    .B2(_045_),
    .Y(_182_));
 sky130_fd_sc_hd__inv_1 _517_ (.A(_288_),
    .Y(_183_));
 sky130_fd_sc_hd__a21oi_1 _518_ (.A1(_130_),
    .A2(_183_),
    .B1(_008_),
    .Y(_184_));
 sky130_fd_sc_hd__a21oi_1 _519_ (.A1(_127_),
    .A2(_285_),
    .B1(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__nand2b_1 _520_ (.A_N(_058_),
    .B(_175_),
    .Y(_186_));
 sky130_fd_sc_hd__o221ai_1 _521_ (.A1(_284_),
    .A2(_086_),
    .B1(_185_),
    .B2(_141_),
    .C1(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__a221oi_1 _522_ (.A1(_226_),
    .A2(_181_),
    .B1(_182_),
    .B2(_038_),
    .C1(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__a21oi_1 _523_ (.A1(_112_),
    .A2(_125_),
    .B1(_188_),
    .Y(_233_));
 sky130_fd_sc_hd__a21oi_1 _524_ (.A1(_021_),
    .A2(_026_),
    .B1(_028_),
    .Y(_189_));
 sky130_fd_sc_hd__mux2i_1 _525_ (.A0(_189_),
    .A1(_157_),
    .S(_019_),
    .Y(_190_));
 sky130_fd_sc_hd__nor3_1 _526_ (.A(_077_),
    .B(_021_),
    .C(_019_),
    .Y(_191_));
 sky130_fd_sc_hd__nand2b_1 _527_ (.A_N(_008_),
    .B(_077_),
    .Y(_192_));
 sky130_fd_sc_hd__nor2_1 _528_ (.A(_292_),
    .B(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__a31oi_1 _529_ (.A1(_076_),
    .A2(_072_),
    .A3(_191_),
    .B1(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__a21oi_1 _530_ (.A1(_130_),
    .A2(_105_),
    .B1(_076_),
    .Y(_195_));
 sky130_fd_sc_hd__a21oi_1 _531_ (.A1(_127_),
    .A2(_293_),
    .B1(_195_),
    .Y(_196_));
 sky130_fd_sc_hd__o22ai_1 _532_ (.A1(_127_),
    .A2(_194_),
    .B1(_196_),
    .B2(_141_),
    .Y(_197_));
 sky130_fd_sc_hd__a221oi_1 _533_ (.A1(_181_),
    .A2(_017_),
    .B1(_190_),
    .B2(_038_),
    .C1(_197_),
    .Y(_198_));
 sky130_fd_sc_hd__a21oi_1 _534_ (.A1(_102_),
    .A2(_112_),
    .B1(_198_),
    .Y(_234_));
 sky130_fd_sc_hd__o21ai_1 _535_ (.A1(_252_),
    .A2(_044_),
    .B1(_048_),
    .Y(_199_));
 sky130_fd_sc_hd__nor2_1 _536_ (.A(_300_),
    .B(_192_),
    .Y(_200_));
 sky130_fd_sc_hd__a31oi_1 _537_ (.A1(_076_),
    .A2(_046_),
    .A3(_191_),
    .B1(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__inv_1 _538_ (.A(_302_),
    .Y(_202_));
 sky130_fd_sc_hd__a21oi_1 _539_ (.A1(_130_),
    .A2(_202_),
    .B1(_076_),
    .Y(_203_));
 sky130_fd_sc_hd__a21oi_1 _540_ (.A1(_127_),
    .A2(_301_),
    .B1(_203_),
    .Y(_204_));
 sky130_fd_sc_hd__o22ai_1 _541_ (.A1(_127_),
    .A2(_201_),
    .B1(_204_),
    .B2(_141_),
    .Y(_205_));
 sky130_fd_sc_hd__a221oi_1 _542_ (.A1(_223_),
    .A2(_181_),
    .B1(_199_),
    .B2(_038_),
    .C1(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__a21oi_1 _543_ (.A1(_111_),
    .A2(_112_),
    .B1(_206_),
    .Y(_235_));
 sky130_fd_sc_hd__inv_1 _544_ (.A(net9),
    .Y(_298_));
 sky130_fd_sc_hd__xnor2_1 _545_ (.A(_298_),
    .B(_222_),
    .Y(_207_));
 sky130_fd_sc_hd__a21oi_1 _546_ (.A1(_105_),
    .A2(_100_),
    .B1(_149_),
    .Y(_208_));
 sky130_fd_sc_hd__a21oi_1 _547_ (.A1(_181_),
    .A2(_207_),
    .B1(_208_),
    .Y(_209_));
 sky130_fd_sc_hd__o22ai_1 _548_ (.A1(_202_),
    .A2(_149_),
    .B1(_209_),
    .B2(_103_),
    .Y(_304_));
 sky130_fd_sc_hd__inv_1 _549_ (.A(net3),
    .Y(_239_));
 sky130_fd_sc_hd__inv_1 _550_ (.A(net5),
    .Y(_266_));
 sky130_fd_sc_hd__inv_1 _551_ (.A(net8),
    .Y(_290_));
 sky130_fd_sc_hd__inv_1 _552_ (.A(_024_),
    .Y(_245_));
 sky130_fd_sc_hd__inv_1 _553_ (.A(net13),
    .Y(_267_));
 sky130_fd_sc_hd__inv_1 _554_ (.A(net14),
    .Y(_275_));
 sky130_fd_sc_hd__inv_1 _555_ (.A(net15),
    .Y(_283_));
 sky130_fd_sc_hd__inv_1 _556_ (.A(net16),
    .Y(_291_));
 sky130_fd_sc_hd__inv_1 _557_ (.A(net17),
    .Y(_299_));
 sky130_fd_sc_hd__fa_1 _558_ (.A(net3),
    .B(net11),
    .CIN(_236_),
    .COUT(_237_),
    .SUM(_238_));
 sky130_fd_sc_hd__fa_1 _559_ (.A(_239_),
    .B(net11),
    .CIN(_240_),
    .COUT(_241_),
    .SUM(_242_));
 sky130_fd_sc_hd__ha_1 _560_ (.A(_244_),
    .B(_245_),
    .COUT(_246_),
    .SUM(_247_));
 sky130_fd_sc_hd__ha_1 _561_ (.A(_244_),
    .B(net10),
    .COUT(_240_),
    .SUM(_248_));
 sky130_fd_sc_hd__ha_1 _562_ (.A(net2),
    .B(_245_),
    .COUT(_249_),
    .SUM(_250_));
 sky130_fd_sc_hd__ha_1 _563_ (.A(net2),
    .B(net10),
    .COUT(_236_),
    .SUM(_251_));
 sky130_fd_sc_hd__ha_1 _564_ (.A(_239_),
    .B(_252_),
    .COUT(_253_),
    .SUM(_243_));
 sky130_fd_sc_hd__ha_1 _565_ (.A(net3),
    .B(_252_),
    .COUT(_254_),
    .SUM(_255_));
 sky130_fd_sc_hd__ha_1 _566_ (.A(net3),
    .B(net11),
    .COUT(_256_),
    .SUM(_257_));
 sky130_fd_sc_hd__ha_1 _567_ (.A(_258_),
    .B(_259_),
    .COUT(_260_),
    .SUM(_261_));
 sky130_fd_sc_hd__ha_1 _568_ (.A(net4),
    .B(_259_),
    .COUT(_262_),
    .SUM(_263_));
 sky130_fd_sc_hd__ha_2 _569_ (.A(net4),
    .B(net12),
    .COUT(_264_),
    .SUM(_265_));
 sky130_fd_sc_hd__ha_1 _570_ (.A(_266_),
    .B(_267_),
    .COUT(_268_),
    .SUM(_269_));
 sky130_fd_sc_hd__ha_1 _571_ (.A(net5),
    .B(_267_),
    .COUT(_270_),
    .SUM(_271_));
 sky130_fd_sc_hd__ha_1 _572_ (.A(net5),
    .B(net13),
    .COUT(_272_),
    .SUM(_273_));
 sky130_fd_sc_hd__ha_1 _573_ (.A(_274_),
    .B(_275_),
    .COUT(_276_),
    .SUM(_277_));
 sky130_fd_sc_hd__ha_1 _574_ (.A(net6),
    .B(_275_),
    .COUT(_278_),
    .SUM(_279_));
 sky130_fd_sc_hd__ha_1 _575_ (.A(net6),
    .B(net14),
    .COUT(_280_),
    .SUM(_281_));
 sky130_fd_sc_hd__ha_2 _576_ (.A(_282_),
    .B(_283_),
    .COUT(_284_),
    .SUM(_285_));
 sky130_fd_sc_hd__ha_1 _577_ (.A(net7),
    .B(_283_),
    .COUT(_286_),
    .SUM(_287_));
 sky130_fd_sc_hd__ha_2 _578_ (.A(net7),
    .B(net15),
    .COUT(_288_),
    .SUM(_289_));
 sky130_fd_sc_hd__ha_2 _579_ (.A(_290_),
    .B(_291_),
    .COUT(_292_),
    .SUM(_293_));
 sky130_fd_sc_hd__ha_1 _580_ (.A(net8),
    .B(_291_),
    .COUT(_294_),
    .SUM(_295_));
 sky130_fd_sc_hd__ha_1 _581_ (.A(net8),
    .B(net16),
    .COUT(_296_),
    .SUM(_297_));
 sky130_fd_sc_hd__ha_1 _582_ (.A(_298_),
    .B(_299_),
    .COUT(_300_),
    .SUM(_301_));
 sky130_fd_sc_hd__ha_1 _583_ (.A(net9),
    .B(net17),
    .COUT(_302_),
    .SUM(_303_));
 sky130_fd_sc_hd__dfrtp_1 \overflow_flag$_DFF_PN0_  (.D(_304_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[0]$_DFF_PN0_  (.D(_228_),
    .Q(net21),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[1]$_DFF_PN0_  (.D(_229_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[2]$_DFF_PN0_  (.D(_230_),
    .Q(net23),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[3]$_DFF_PN0_  (.D(_231_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[4]$_DFF_PN0_  (.D(_232_),
    .Q(net25),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[5]$_DFF_PN0_  (.D(_233_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[6]$_DFF_PN0_  (.D(_234_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[7]$_DFF_PN0_  (.D(_235_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \zero_flag$_DFF_PN0_  (.D(_000_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 hold1 (.A(net30),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_47 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(a[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(a[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input3 (.A(a[2]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input4 (.A(a[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input5 (.A(a[4]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input6 (.A(a[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(a[6]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input8 (.A(a[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(b[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(b[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(b[2]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(b[3]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(b[4]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(b[5]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(b[6]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(b[7]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(op_code[0]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(op_code[2]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(overflow_flag));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(result[0]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(result[1]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(result[2]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(result[3]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(result[4]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(result[5]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(result[6]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(result[7]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(zero_flag));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net30));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_124 ();
endmodule
