module register_file (clk,
    read_en1,
    read_en2,
    rst_n,
    write_en,
    read_addr1,
    read_addr2,
    read_data1,
    read_data2,
    write_addr,
    write_data);
 input clk;
 input read_en1;
 input read_en2;
 input rst_n;
 input write_en;
 input [4:0] read_addr1;
 input [4:0] read_addr2;
 output [31:0] read_data1;
 output [31:0] read_data2;
 input [4:0] write_addr;
 input [31:0] write_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire \registers[0][0] ;
 wire \registers[0][10] ;
 wire \registers[0][11] ;
 wire \registers[0][12] ;
 wire \registers[0][13] ;
 wire \registers[0][14] ;
 wire \registers[0][15] ;
 wire \registers[0][16] ;
 wire \registers[0][17] ;
 wire \registers[0][18] ;
 wire \registers[0][19] ;
 wire \registers[0][1] ;
 wire \registers[0][20] ;
 wire \registers[0][21] ;
 wire \registers[0][22] ;
 wire \registers[0][23] ;
 wire \registers[0][24] ;
 wire \registers[0][25] ;
 wire \registers[0][26] ;
 wire \registers[0][27] ;
 wire \registers[0][28] ;
 wire \registers[0][29] ;
 wire \registers[0][2] ;
 wire \registers[0][30] ;
 wire \registers[0][31] ;
 wire \registers[0][3] ;
 wire \registers[0][4] ;
 wire \registers[0][5] ;
 wire \registers[0][6] ;
 wire \registers[0][7] ;
 wire \registers[0][8] ;
 wire \registers[0][9] ;
 wire \registers[10][0] ;
 wire \registers[10][10] ;
 wire \registers[10][11] ;
 wire \registers[10][12] ;
 wire \registers[10][13] ;
 wire \registers[10][14] ;
 wire \registers[10][15] ;
 wire \registers[10][16] ;
 wire \registers[10][17] ;
 wire \registers[10][18] ;
 wire \registers[10][19] ;
 wire \registers[10][1] ;
 wire \registers[10][20] ;
 wire \registers[10][21] ;
 wire \registers[10][22] ;
 wire \registers[10][23] ;
 wire \registers[10][24] ;
 wire \registers[10][25] ;
 wire \registers[10][26] ;
 wire \registers[10][27] ;
 wire \registers[10][28] ;
 wire \registers[10][29] ;
 wire \registers[10][2] ;
 wire \registers[10][30] ;
 wire \registers[10][31] ;
 wire \registers[10][3] ;
 wire \registers[10][4] ;
 wire \registers[10][5] ;
 wire \registers[10][6] ;
 wire \registers[10][7] ;
 wire \registers[10][8] ;
 wire \registers[10][9] ;
 wire \registers[11][0] ;
 wire \registers[11][10] ;
 wire \registers[11][11] ;
 wire \registers[11][12] ;
 wire \registers[11][13] ;
 wire \registers[11][14] ;
 wire \registers[11][15] ;
 wire \registers[11][16] ;
 wire \registers[11][17] ;
 wire \registers[11][18] ;
 wire \registers[11][19] ;
 wire \registers[11][1] ;
 wire \registers[11][20] ;
 wire \registers[11][21] ;
 wire \registers[11][22] ;
 wire \registers[11][23] ;
 wire \registers[11][24] ;
 wire \registers[11][25] ;
 wire \registers[11][26] ;
 wire \registers[11][27] ;
 wire \registers[11][28] ;
 wire \registers[11][29] ;
 wire \registers[11][2] ;
 wire \registers[11][30] ;
 wire \registers[11][31] ;
 wire \registers[11][3] ;
 wire \registers[11][4] ;
 wire \registers[11][5] ;
 wire \registers[11][6] ;
 wire \registers[11][7] ;
 wire \registers[11][8] ;
 wire \registers[11][9] ;
 wire \registers[12][0] ;
 wire \registers[12][10] ;
 wire \registers[12][11] ;
 wire \registers[12][12] ;
 wire \registers[12][13] ;
 wire \registers[12][14] ;
 wire \registers[12][15] ;
 wire \registers[12][16] ;
 wire \registers[12][17] ;
 wire \registers[12][18] ;
 wire \registers[12][19] ;
 wire \registers[12][1] ;
 wire \registers[12][20] ;
 wire \registers[12][21] ;
 wire \registers[12][22] ;
 wire \registers[12][23] ;
 wire \registers[12][24] ;
 wire \registers[12][25] ;
 wire \registers[12][26] ;
 wire \registers[12][27] ;
 wire \registers[12][28] ;
 wire \registers[12][29] ;
 wire \registers[12][2] ;
 wire \registers[12][30] ;
 wire \registers[12][31] ;
 wire \registers[12][3] ;
 wire \registers[12][4] ;
 wire \registers[12][5] ;
 wire \registers[12][6] ;
 wire \registers[12][7] ;
 wire \registers[12][8] ;
 wire \registers[12][9] ;
 wire \registers[13][0] ;
 wire \registers[13][10] ;
 wire \registers[13][11] ;
 wire \registers[13][12] ;
 wire \registers[13][13] ;
 wire \registers[13][14] ;
 wire \registers[13][15] ;
 wire \registers[13][16] ;
 wire \registers[13][17] ;
 wire \registers[13][18] ;
 wire \registers[13][19] ;
 wire \registers[13][1] ;
 wire \registers[13][20] ;
 wire \registers[13][21] ;
 wire \registers[13][22] ;
 wire \registers[13][23] ;
 wire \registers[13][24] ;
 wire \registers[13][25] ;
 wire \registers[13][26] ;
 wire \registers[13][27] ;
 wire \registers[13][28] ;
 wire \registers[13][29] ;
 wire \registers[13][2] ;
 wire \registers[13][30] ;
 wire \registers[13][31] ;
 wire \registers[13][3] ;
 wire \registers[13][4] ;
 wire \registers[13][5] ;
 wire \registers[13][6] ;
 wire \registers[13][7] ;
 wire \registers[13][8] ;
 wire \registers[13][9] ;
 wire \registers[14][0] ;
 wire \registers[14][10] ;
 wire \registers[14][11] ;
 wire \registers[14][12] ;
 wire \registers[14][13] ;
 wire \registers[14][14] ;
 wire \registers[14][15] ;
 wire \registers[14][16] ;
 wire \registers[14][17] ;
 wire \registers[14][18] ;
 wire \registers[14][19] ;
 wire \registers[14][1] ;
 wire \registers[14][20] ;
 wire \registers[14][21] ;
 wire \registers[14][22] ;
 wire \registers[14][23] ;
 wire \registers[14][24] ;
 wire \registers[14][25] ;
 wire \registers[14][26] ;
 wire \registers[14][27] ;
 wire \registers[14][28] ;
 wire \registers[14][29] ;
 wire \registers[14][2] ;
 wire \registers[14][30] ;
 wire \registers[14][31] ;
 wire \registers[14][3] ;
 wire \registers[14][4] ;
 wire \registers[14][5] ;
 wire \registers[14][6] ;
 wire \registers[14][7] ;
 wire \registers[14][8] ;
 wire \registers[14][9] ;
 wire \registers[15][0] ;
 wire \registers[15][10] ;
 wire \registers[15][11] ;
 wire \registers[15][12] ;
 wire \registers[15][13] ;
 wire \registers[15][14] ;
 wire \registers[15][15] ;
 wire \registers[15][16] ;
 wire \registers[15][17] ;
 wire \registers[15][18] ;
 wire \registers[15][19] ;
 wire \registers[15][1] ;
 wire \registers[15][20] ;
 wire \registers[15][21] ;
 wire \registers[15][22] ;
 wire \registers[15][23] ;
 wire \registers[15][24] ;
 wire \registers[15][25] ;
 wire \registers[15][26] ;
 wire \registers[15][27] ;
 wire \registers[15][28] ;
 wire \registers[15][29] ;
 wire \registers[15][2] ;
 wire \registers[15][30] ;
 wire \registers[15][31] ;
 wire \registers[15][3] ;
 wire \registers[15][4] ;
 wire \registers[15][5] ;
 wire \registers[15][6] ;
 wire \registers[15][7] ;
 wire \registers[15][8] ;
 wire \registers[15][9] ;
 wire \registers[16][0] ;
 wire \registers[16][10] ;
 wire \registers[16][11] ;
 wire \registers[16][12] ;
 wire \registers[16][13] ;
 wire \registers[16][14] ;
 wire \registers[16][15] ;
 wire \registers[16][16] ;
 wire \registers[16][17] ;
 wire \registers[16][18] ;
 wire \registers[16][19] ;
 wire \registers[16][1] ;
 wire \registers[16][20] ;
 wire \registers[16][21] ;
 wire \registers[16][22] ;
 wire \registers[16][23] ;
 wire \registers[16][24] ;
 wire \registers[16][25] ;
 wire \registers[16][26] ;
 wire \registers[16][27] ;
 wire \registers[16][28] ;
 wire \registers[16][29] ;
 wire \registers[16][2] ;
 wire \registers[16][30] ;
 wire \registers[16][31] ;
 wire \registers[16][3] ;
 wire \registers[16][4] ;
 wire \registers[16][5] ;
 wire \registers[16][6] ;
 wire \registers[16][7] ;
 wire \registers[16][8] ;
 wire \registers[16][9] ;
 wire \registers[17][0] ;
 wire \registers[17][10] ;
 wire \registers[17][11] ;
 wire \registers[17][12] ;
 wire \registers[17][13] ;
 wire \registers[17][14] ;
 wire \registers[17][15] ;
 wire \registers[17][16] ;
 wire \registers[17][17] ;
 wire \registers[17][18] ;
 wire \registers[17][19] ;
 wire \registers[17][1] ;
 wire \registers[17][20] ;
 wire \registers[17][21] ;
 wire \registers[17][22] ;
 wire \registers[17][23] ;
 wire \registers[17][24] ;
 wire \registers[17][25] ;
 wire \registers[17][26] ;
 wire \registers[17][27] ;
 wire \registers[17][28] ;
 wire \registers[17][29] ;
 wire \registers[17][2] ;
 wire \registers[17][30] ;
 wire \registers[17][31] ;
 wire \registers[17][3] ;
 wire \registers[17][4] ;
 wire \registers[17][5] ;
 wire \registers[17][6] ;
 wire \registers[17][7] ;
 wire \registers[17][8] ;
 wire \registers[17][9] ;
 wire \registers[18][0] ;
 wire \registers[18][10] ;
 wire \registers[18][11] ;
 wire \registers[18][12] ;
 wire \registers[18][13] ;
 wire \registers[18][14] ;
 wire \registers[18][15] ;
 wire \registers[18][16] ;
 wire \registers[18][17] ;
 wire \registers[18][18] ;
 wire \registers[18][19] ;
 wire \registers[18][1] ;
 wire \registers[18][20] ;
 wire \registers[18][21] ;
 wire \registers[18][22] ;
 wire \registers[18][23] ;
 wire \registers[18][24] ;
 wire \registers[18][25] ;
 wire \registers[18][26] ;
 wire \registers[18][27] ;
 wire \registers[18][28] ;
 wire \registers[18][29] ;
 wire \registers[18][2] ;
 wire \registers[18][30] ;
 wire \registers[18][31] ;
 wire \registers[18][3] ;
 wire \registers[18][4] ;
 wire \registers[18][5] ;
 wire \registers[18][6] ;
 wire \registers[18][7] ;
 wire \registers[18][8] ;
 wire \registers[18][9] ;
 wire \registers[19][0] ;
 wire \registers[19][10] ;
 wire \registers[19][11] ;
 wire \registers[19][12] ;
 wire \registers[19][13] ;
 wire \registers[19][14] ;
 wire \registers[19][15] ;
 wire \registers[19][16] ;
 wire \registers[19][17] ;
 wire \registers[19][18] ;
 wire \registers[19][19] ;
 wire \registers[19][1] ;
 wire \registers[19][20] ;
 wire \registers[19][21] ;
 wire \registers[19][22] ;
 wire \registers[19][23] ;
 wire \registers[19][24] ;
 wire \registers[19][25] ;
 wire \registers[19][26] ;
 wire \registers[19][27] ;
 wire \registers[19][28] ;
 wire \registers[19][29] ;
 wire \registers[19][2] ;
 wire \registers[19][30] ;
 wire \registers[19][31] ;
 wire \registers[19][3] ;
 wire \registers[19][4] ;
 wire \registers[19][5] ;
 wire \registers[19][6] ;
 wire \registers[19][7] ;
 wire \registers[19][8] ;
 wire \registers[19][9] ;
 wire \registers[1][0] ;
 wire \registers[1][10] ;
 wire \registers[1][11] ;
 wire \registers[1][12] ;
 wire \registers[1][13] ;
 wire \registers[1][14] ;
 wire \registers[1][15] ;
 wire \registers[1][16] ;
 wire \registers[1][17] ;
 wire \registers[1][18] ;
 wire \registers[1][19] ;
 wire \registers[1][1] ;
 wire \registers[1][20] ;
 wire \registers[1][21] ;
 wire \registers[1][22] ;
 wire \registers[1][23] ;
 wire \registers[1][24] ;
 wire \registers[1][25] ;
 wire \registers[1][26] ;
 wire \registers[1][27] ;
 wire \registers[1][28] ;
 wire \registers[1][29] ;
 wire \registers[1][2] ;
 wire \registers[1][30] ;
 wire \registers[1][31] ;
 wire \registers[1][3] ;
 wire \registers[1][4] ;
 wire \registers[1][5] ;
 wire \registers[1][6] ;
 wire \registers[1][7] ;
 wire \registers[1][8] ;
 wire \registers[1][9] ;
 wire \registers[20][0] ;
 wire \registers[20][10] ;
 wire \registers[20][11] ;
 wire \registers[20][12] ;
 wire \registers[20][13] ;
 wire \registers[20][14] ;
 wire \registers[20][15] ;
 wire \registers[20][16] ;
 wire \registers[20][17] ;
 wire \registers[20][18] ;
 wire \registers[20][19] ;
 wire \registers[20][1] ;
 wire \registers[20][20] ;
 wire \registers[20][21] ;
 wire \registers[20][22] ;
 wire \registers[20][23] ;
 wire \registers[20][24] ;
 wire \registers[20][25] ;
 wire \registers[20][26] ;
 wire \registers[20][27] ;
 wire \registers[20][28] ;
 wire \registers[20][29] ;
 wire \registers[20][2] ;
 wire \registers[20][30] ;
 wire \registers[20][31] ;
 wire \registers[20][3] ;
 wire \registers[20][4] ;
 wire \registers[20][5] ;
 wire \registers[20][6] ;
 wire \registers[20][7] ;
 wire \registers[20][8] ;
 wire \registers[20][9] ;
 wire \registers[21][0] ;
 wire \registers[21][10] ;
 wire \registers[21][11] ;
 wire \registers[21][12] ;
 wire \registers[21][13] ;
 wire \registers[21][14] ;
 wire \registers[21][15] ;
 wire \registers[21][16] ;
 wire \registers[21][17] ;
 wire \registers[21][18] ;
 wire \registers[21][19] ;
 wire \registers[21][1] ;
 wire \registers[21][20] ;
 wire \registers[21][21] ;
 wire \registers[21][22] ;
 wire \registers[21][23] ;
 wire \registers[21][24] ;
 wire \registers[21][25] ;
 wire \registers[21][26] ;
 wire \registers[21][27] ;
 wire \registers[21][28] ;
 wire \registers[21][29] ;
 wire \registers[21][2] ;
 wire \registers[21][30] ;
 wire \registers[21][31] ;
 wire \registers[21][3] ;
 wire \registers[21][4] ;
 wire \registers[21][5] ;
 wire \registers[21][6] ;
 wire \registers[21][7] ;
 wire \registers[21][8] ;
 wire \registers[21][9] ;
 wire \registers[22][0] ;
 wire \registers[22][10] ;
 wire \registers[22][11] ;
 wire \registers[22][12] ;
 wire \registers[22][13] ;
 wire \registers[22][14] ;
 wire \registers[22][15] ;
 wire \registers[22][16] ;
 wire \registers[22][17] ;
 wire \registers[22][18] ;
 wire \registers[22][19] ;
 wire \registers[22][1] ;
 wire \registers[22][20] ;
 wire \registers[22][21] ;
 wire \registers[22][22] ;
 wire \registers[22][23] ;
 wire \registers[22][24] ;
 wire \registers[22][25] ;
 wire \registers[22][26] ;
 wire \registers[22][27] ;
 wire \registers[22][28] ;
 wire \registers[22][29] ;
 wire \registers[22][2] ;
 wire \registers[22][30] ;
 wire \registers[22][31] ;
 wire \registers[22][3] ;
 wire \registers[22][4] ;
 wire \registers[22][5] ;
 wire \registers[22][6] ;
 wire \registers[22][7] ;
 wire \registers[22][8] ;
 wire \registers[22][9] ;
 wire \registers[23][0] ;
 wire \registers[23][10] ;
 wire \registers[23][11] ;
 wire \registers[23][12] ;
 wire \registers[23][13] ;
 wire \registers[23][14] ;
 wire \registers[23][15] ;
 wire \registers[23][16] ;
 wire \registers[23][17] ;
 wire \registers[23][18] ;
 wire \registers[23][19] ;
 wire \registers[23][1] ;
 wire \registers[23][20] ;
 wire \registers[23][21] ;
 wire \registers[23][22] ;
 wire \registers[23][23] ;
 wire \registers[23][24] ;
 wire \registers[23][25] ;
 wire \registers[23][26] ;
 wire \registers[23][27] ;
 wire \registers[23][28] ;
 wire \registers[23][29] ;
 wire \registers[23][2] ;
 wire \registers[23][30] ;
 wire \registers[23][31] ;
 wire \registers[23][3] ;
 wire \registers[23][4] ;
 wire \registers[23][5] ;
 wire \registers[23][6] ;
 wire \registers[23][7] ;
 wire \registers[23][8] ;
 wire \registers[23][9] ;
 wire \registers[24][0] ;
 wire \registers[24][10] ;
 wire \registers[24][11] ;
 wire \registers[24][12] ;
 wire \registers[24][13] ;
 wire \registers[24][14] ;
 wire \registers[24][15] ;
 wire \registers[24][16] ;
 wire \registers[24][17] ;
 wire \registers[24][18] ;
 wire \registers[24][19] ;
 wire \registers[24][1] ;
 wire \registers[24][20] ;
 wire \registers[24][21] ;
 wire \registers[24][22] ;
 wire \registers[24][23] ;
 wire \registers[24][24] ;
 wire \registers[24][25] ;
 wire \registers[24][26] ;
 wire \registers[24][27] ;
 wire \registers[24][28] ;
 wire \registers[24][29] ;
 wire \registers[24][2] ;
 wire \registers[24][30] ;
 wire \registers[24][31] ;
 wire \registers[24][3] ;
 wire \registers[24][4] ;
 wire \registers[24][5] ;
 wire \registers[24][6] ;
 wire \registers[24][7] ;
 wire \registers[24][8] ;
 wire \registers[24][9] ;
 wire \registers[25][0] ;
 wire \registers[25][10] ;
 wire \registers[25][11] ;
 wire \registers[25][12] ;
 wire \registers[25][13] ;
 wire \registers[25][14] ;
 wire \registers[25][15] ;
 wire \registers[25][16] ;
 wire \registers[25][17] ;
 wire \registers[25][18] ;
 wire \registers[25][19] ;
 wire \registers[25][1] ;
 wire \registers[25][20] ;
 wire \registers[25][21] ;
 wire \registers[25][22] ;
 wire \registers[25][23] ;
 wire \registers[25][24] ;
 wire \registers[25][25] ;
 wire \registers[25][26] ;
 wire \registers[25][27] ;
 wire \registers[25][28] ;
 wire \registers[25][29] ;
 wire \registers[25][2] ;
 wire \registers[25][30] ;
 wire \registers[25][31] ;
 wire \registers[25][3] ;
 wire \registers[25][4] ;
 wire \registers[25][5] ;
 wire \registers[25][6] ;
 wire \registers[25][7] ;
 wire \registers[25][8] ;
 wire \registers[25][9] ;
 wire \registers[26][0] ;
 wire \registers[26][10] ;
 wire \registers[26][11] ;
 wire \registers[26][12] ;
 wire \registers[26][13] ;
 wire \registers[26][14] ;
 wire \registers[26][15] ;
 wire \registers[26][16] ;
 wire \registers[26][17] ;
 wire \registers[26][18] ;
 wire \registers[26][19] ;
 wire \registers[26][1] ;
 wire \registers[26][20] ;
 wire \registers[26][21] ;
 wire \registers[26][22] ;
 wire \registers[26][23] ;
 wire \registers[26][24] ;
 wire \registers[26][25] ;
 wire \registers[26][26] ;
 wire \registers[26][27] ;
 wire \registers[26][28] ;
 wire \registers[26][29] ;
 wire \registers[26][2] ;
 wire \registers[26][30] ;
 wire \registers[26][31] ;
 wire \registers[26][3] ;
 wire \registers[26][4] ;
 wire \registers[26][5] ;
 wire \registers[26][6] ;
 wire \registers[26][7] ;
 wire \registers[26][8] ;
 wire \registers[26][9] ;
 wire \registers[27][0] ;
 wire \registers[27][10] ;
 wire \registers[27][11] ;
 wire \registers[27][12] ;
 wire \registers[27][13] ;
 wire \registers[27][14] ;
 wire \registers[27][15] ;
 wire \registers[27][16] ;
 wire \registers[27][17] ;
 wire \registers[27][18] ;
 wire \registers[27][19] ;
 wire \registers[27][1] ;
 wire \registers[27][20] ;
 wire \registers[27][21] ;
 wire \registers[27][22] ;
 wire \registers[27][23] ;
 wire \registers[27][24] ;
 wire \registers[27][25] ;
 wire \registers[27][26] ;
 wire \registers[27][27] ;
 wire \registers[27][28] ;
 wire \registers[27][29] ;
 wire \registers[27][2] ;
 wire \registers[27][30] ;
 wire \registers[27][31] ;
 wire \registers[27][3] ;
 wire \registers[27][4] ;
 wire \registers[27][5] ;
 wire \registers[27][6] ;
 wire \registers[27][7] ;
 wire \registers[27][8] ;
 wire \registers[27][9] ;
 wire \registers[28][0] ;
 wire \registers[28][10] ;
 wire \registers[28][11] ;
 wire \registers[28][12] ;
 wire \registers[28][13] ;
 wire \registers[28][14] ;
 wire \registers[28][15] ;
 wire \registers[28][16] ;
 wire \registers[28][17] ;
 wire \registers[28][18] ;
 wire \registers[28][19] ;
 wire \registers[28][1] ;
 wire \registers[28][20] ;
 wire \registers[28][21] ;
 wire \registers[28][22] ;
 wire \registers[28][23] ;
 wire \registers[28][24] ;
 wire \registers[28][25] ;
 wire \registers[28][26] ;
 wire \registers[28][27] ;
 wire \registers[28][28] ;
 wire \registers[28][29] ;
 wire \registers[28][2] ;
 wire \registers[28][30] ;
 wire \registers[28][31] ;
 wire \registers[28][3] ;
 wire \registers[28][4] ;
 wire \registers[28][5] ;
 wire \registers[28][6] ;
 wire \registers[28][7] ;
 wire \registers[28][8] ;
 wire \registers[28][9] ;
 wire \registers[29][0] ;
 wire \registers[29][10] ;
 wire \registers[29][11] ;
 wire \registers[29][12] ;
 wire \registers[29][13] ;
 wire \registers[29][14] ;
 wire \registers[29][15] ;
 wire \registers[29][16] ;
 wire \registers[29][17] ;
 wire \registers[29][18] ;
 wire \registers[29][19] ;
 wire \registers[29][1] ;
 wire \registers[29][20] ;
 wire \registers[29][21] ;
 wire \registers[29][22] ;
 wire \registers[29][23] ;
 wire \registers[29][24] ;
 wire \registers[29][25] ;
 wire \registers[29][26] ;
 wire \registers[29][27] ;
 wire \registers[29][28] ;
 wire \registers[29][29] ;
 wire \registers[29][2] ;
 wire \registers[29][30] ;
 wire \registers[29][31] ;
 wire \registers[29][3] ;
 wire \registers[29][4] ;
 wire \registers[29][5] ;
 wire \registers[29][6] ;
 wire \registers[29][7] ;
 wire \registers[29][8] ;
 wire \registers[29][9] ;
 wire \registers[2][0] ;
 wire \registers[2][10] ;
 wire \registers[2][11] ;
 wire \registers[2][12] ;
 wire \registers[2][13] ;
 wire \registers[2][14] ;
 wire \registers[2][15] ;
 wire \registers[2][16] ;
 wire \registers[2][17] ;
 wire \registers[2][18] ;
 wire \registers[2][19] ;
 wire \registers[2][1] ;
 wire \registers[2][20] ;
 wire \registers[2][21] ;
 wire \registers[2][22] ;
 wire \registers[2][23] ;
 wire \registers[2][24] ;
 wire \registers[2][25] ;
 wire \registers[2][26] ;
 wire \registers[2][27] ;
 wire \registers[2][28] ;
 wire \registers[2][29] ;
 wire \registers[2][2] ;
 wire \registers[2][30] ;
 wire \registers[2][31] ;
 wire \registers[2][3] ;
 wire \registers[2][4] ;
 wire \registers[2][5] ;
 wire \registers[2][6] ;
 wire \registers[2][7] ;
 wire \registers[2][8] ;
 wire \registers[2][9] ;
 wire \registers[30][0] ;
 wire \registers[30][10] ;
 wire \registers[30][11] ;
 wire \registers[30][12] ;
 wire \registers[30][13] ;
 wire \registers[30][14] ;
 wire \registers[30][15] ;
 wire \registers[30][16] ;
 wire \registers[30][17] ;
 wire \registers[30][18] ;
 wire \registers[30][19] ;
 wire \registers[30][1] ;
 wire \registers[30][20] ;
 wire \registers[30][21] ;
 wire \registers[30][22] ;
 wire \registers[30][23] ;
 wire \registers[30][24] ;
 wire \registers[30][25] ;
 wire \registers[30][26] ;
 wire \registers[30][27] ;
 wire \registers[30][28] ;
 wire \registers[30][29] ;
 wire \registers[30][2] ;
 wire \registers[30][30] ;
 wire \registers[30][31] ;
 wire \registers[30][3] ;
 wire \registers[30][4] ;
 wire \registers[30][5] ;
 wire \registers[30][6] ;
 wire \registers[30][7] ;
 wire \registers[30][8] ;
 wire \registers[30][9] ;
 wire \registers[31][0] ;
 wire \registers[31][10] ;
 wire \registers[31][11] ;
 wire \registers[31][12] ;
 wire \registers[31][13] ;
 wire \registers[31][14] ;
 wire \registers[31][15] ;
 wire \registers[31][16] ;
 wire \registers[31][17] ;
 wire \registers[31][18] ;
 wire \registers[31][19] ;
 wire \registers[31][1] ;
 wire \registers[31][20] ;
 wire \registers[31][21] ;
 wire \registers[31][22] ;
 wire \registers[31][23] ;
 wire \registers[31][24] ;
 wire \registers[31][25] ;
 wire \registers[31][26] ;
 wire \registers[31][27] ;
 wire \registers[31][28] ;
 wire \registers[31][29] ;
 wire \registers[31][2] ;
 wire \registers[31][30] ;
 wire \registers[31][31] ;
 wire \registers[31][3] ;
 wire \registers[31][4] ;
 wire \registers[31][5] ;
 wire \registers[31][6] ;
 wire \registers[31][7] ;
 wire \registers[31][8] ;
 wire \registers[31][9] ;
 wire \registers[3][0] ;
 wire \registers[3][10] ;
 wire \registers[3][11] ;
 wire \registers[3][12] ;
 wire \registers[3][13] ;
 wire \registers[3][14] ;
 wire \registers[3][15] ;
 wire \registers[3][16] ;
 wire \registers[3][17] ;
 wire \registers[3][18] ;
 wire \registers[3][19] ;
 wire \registers[3][1] ;
 wire \registers[3][20] ;
 wire \registers[3][21] ;
 wire \registers[3][22] ;
 wire \registers[3][23] ;
 wire \registers[3][24] ;
 wire \registers[3][25] ;
 wire \registers[3][26] ;
 wire \registers[3][27] ;
 wire \registers[3][28] ;
 wire \registers[3][29] ;
 wire \registers[3][2] ;
 wire \registers[3][30] ;
 wire \registers[3][31] ;
 wire \registers[3][3] ;
 wire \registers[3][4] ;
 wire \registers[3][5] ;
 wire \registers[3][6] ;
 wire \registers[3][7] ;
 wire \registers[3][8] ;
 wire \registers[3][9] ;
 wire \registers[4][0] ;
 wire \registers[4][10] ;
 wire \registers[4][11] ;
 wire \registers[4][12] ;
 wire \registers[4][13] ;
 wire \registers[4][14] ;
 wire \registers[4][15] ;
 wire \registers[4][16] ;
 wire \registers[4][17] ;
 wire \registers[4][18] ;
 wire \registers[4][19] ;
 wire \registers[4][1] ;
 wire \registers[4][20] ;
 wire \registers[4][21] ;
 wire \registers[4][22] ;
 wire \registers[4][23] ;
 wire \registers[4][24] ;
 wire \registers[4][25] ;
 wire \registers[4][26] ;
 wire \registers[4][27] ;
 wire \registers[4][28] ;
 wire \registers[4][29] ;
 wire \registers[4][2] ;
 wire \registers[4][30] ;
 wire \registers[4][31] ;
 wire \registers[4][3] ;
 wire \registers[4][4] ;
 wire \registers[4][5] ;
 wire \registers[4][6] ;
 wire \registers[4][7] ;
 wire \registers[4][8] ;
 wire \registers[4][9] ;
 wire \registers[5][0] ;
 wire \registers[5][10] ;
 wire \registers[5][11] ;
 wire \registers[5][12] ;
 wire \registers[5][13] ;
 wire \registers[5][14] ;
 wire \registers[5][15] ;
 wire \registers[5][16] ;
 wire \registers[5][17] ;
 wire \registers[5][18] ;
 wire \registers[5][19] ;
 wire \registers[5][1] ;
 wire \registers[5][20] ;
 wire \registers[5][21] ;
 wire \registers[5][22] ;
 wire \registers[5][23] ;
 wire \registers[5][24] ;
 wire \registers[5][25] ;
 wire \registers[5][26] ;
 wire \registers[5][27] ;
 wire \registers[5][28] ;
 wire \registers[5][29] ;
 wire \registers[5][2] ;
 wire \registers[5][30] ;
 wire \registers[5][31] ;
 wire \registers[5][3] ;
 wire \registers[5][4] ;
 wire \registers[5][5] ;
 wire \registers[5][6] ;
 wire \registers[5][7] ;
 wire \registers[5][8] ;
 wire \registers[5][9] ;
 wire \registers[6][0] ;
 wire \registers[6][10] ;
 wire \registers[6][11] ;
 wire \registers[6][12] ;
 wire \registers[6][13] ;
 wire \registers[6][14] ;
 wire \registers[6][15] ;
 wire \registers[6][16] ;
 wire \registers[6][17] ;
 wire \registers[6][18] ;
 wire \registers[6][19] ;
 wire \registers[6][1] ;
 wire \registers[6][20] ;
 wire \registers[6][21] ;
 wire \registers[6][22] ;
 wire \registers[6][23] ;
 wire \registers[6][24] ;
 wire \registers[6][25] ;
 wire \registers[6][26] ;
 wire \registers[6][27] ;
 wire \registers[6][28] ;
 wire \registers[6][29] ;
 wire \registers[6][2] ;
 wire \registers[6][30] ;
 wire \registers[6][31] ;
 wire \registers[6][3] ;
 wire \registers[6][4] ;
 wire \registers[6][5] ;
 wire \registers[6][6] ;
 wire \registers[6][7] ;
 wire \registers[6][8] ;
 wire \registers[6][9] ;
 wire \registers[7][0] ;
 wire \registers[7][10] ;
 wire \registers[7][11] ;
 wire \registers[7][12] ;
 wire \registers[7][13] ;
 wire \registers[7][14] ;
 wire \registers[7][15] ;
 wire \registers[7][16] ;
 wire \registers[7][17] ;
 wire \registers[7][18] ;
 wire \registers[7][19] ;
 wire \registers[7][1] ;
 wire \registers[7][20] ;
 wire \registers[7][21] ;
 wire \registers[7][22] ;
 wire \registers[7][23] ;
 wire \registers[7][24] ;
 wire \registers[7][25] ;
 wire \registers[7][26] ;
 wire \registers[7][27] ;
 wire \registers[7][28] ;
 wire \registers[7][29] ;
 wire \registers[7][2] ;
 wire \registers[7][30] ;
 wire \registers[7][31] ;
 wire \registers[7][3] ;
 wire \registers[7][4] ;
 wire \registers[7][5] ;
 wire \registers[7][6] ;
 wire \registers[7][7] ;
 wire \registers[7][8] ;
 wire \registers[7][9] ;
 wire \registers[8][0] ;
 wire \registers[8][10] ;
 wire \registers[8][11] ;
 wire \registers[8][12] ;
 wire \registers[8][13] ;
 wire \registers[8][14] ;
 wire \registers[8][15] ;
 wire \registers[8][16] ;
 wire \registers[8][17] ;
 wire \registers[8][18] ;
 wire \registers[8][19] ;
 wire \registers[8][1] ;
 wire \registers[8][20] ;
 wire \registers[8][21] ;
 wire \registers[8][22] ;
 wire \registers[8][23] ;
 wire \registers[8][24] ;
 wire \registers[8][25] ;
 wire \registers[8][26] ;
 wire \registers[8][27] ;
 wire \registers[8][28] ;
 wire \registers[8][29] ;
 wire \registers[8][2] ;
 wire \registers[8][30] ;
 wire \registers[8][31] ;
 wire \registers[8][3] ;
 wire \registers[8][4] ;
 wire \registers[8][5] ;
 wire \registers[8][6] ;
 wire \registers[8][7] ;
 wire \registers[8][8] ;
 wire \registers[8][9] ;
 wire \registers[9][0] ;
 wire \registers[9][10] ;
 wire \registers[9][11] ;
 wire \registers[9][12] ;
 wire \registers[9][13] ;
 wire \registers[9][14] ;
 wire \registers[9][15] ;
 wire \registers[9][16] ;
 wire \registers[9][17] ;
 wire \registers[9][18] ;
 wire \registers[9][19] ;
 wire \registers[9][1] ;
 wire \registers[9][20] ;
 wire \registers[9][21] ;
 wire \registers[9][22] ;
 wire \registers[9][23] ;
 wire \registers[9][24] ;
 wire \registers[9][25] ;
 wire \registers[9][26] ;
 wire \registers[9][27] ;
 wire \registers[9][28] ;
 wire \registers[9][29] ;
 wire \registers[9][2] ;
 wire \registers[9][30] ;
 wire \registers[9][31] ;
 wire \registers[9][3] ;
 wire \registers[9][4] ;
 wire \registers[9][5] ;
 wire \registers[9][6] ;
 wire \registers[9][7] ;
 wire \registers[9][8] ;
 wire \registers[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 CLKBUF_X3 _06970_ (.A(write_data[31]),
    .Z(_01088_));
 BUF_X4 _06971_ (.A(_01088_),
    .Z(_01089_));
 BUF_X4 _06972_ (.A(net3),
    .Z(_01090_));
 BUF_X4 _06973_ (.A(write_addr[4]),
    .Z(_01091_));
 BUF_X4 _06974_ (.A(write_addr[2]),
    .Z(_01092_));
 NAND3_X2 _06975_ (.A1(_01090_),
    .A2(_01091_),
    .A3(_01092_),
    .ZN(_01093_));
 BUF_X4 _06976_ (.A(write_addr[1]),
    .Z(_01094_));
 BUF_X2 _06977_ (.A(rst_n),
    .Z(_01095_));
 CLKBUF_X3 _06978_ (.A(write_addr[0]),
    .Z(_01096_));
 NAND3_X1 _06979_ (.A1(_01095_),
    .A2(_01096_),
    .A3(net4),
    .ZN(_01097_));
 OR2_X2 _06980_ (.A1(_01094_),
    .A2(_01097_),
    .ZN(_01098_));
 NOR2_X1 _06981_ (.A1(_01093_),
    .A2(_01098_),
    .ZN(_01099_));
 BUF_X4 _06982_ (.A(_01099_),
    .Z(_01100_));
 BUF_X4 _06983_ (.A(_01100_),
    .Z(_01101_));
 NAND2_X1 _06984_ (.A1(_01089_),
    .A2(_01101_),
    .ZN(_01102_));
 BUF_X4 _06985_ (.A(_01095_),
    .Z(_01103_));
 BUF_X4 _06986_ (.A(_01103_),
    .Z(_01104_));
 BUF_X4 _06987_ (.A(_01104_),
    .Z(_01105_));
 NAND2_X1 _06988_ (.A1(_01105_),
    .A2(\registers[29][31] ),
    .ZN(_01106_));
 BUF_X4 _06989_ (.A(_01100_),
    .Z(_01107_));
 OAI21_X1 _06990_ (.A(_01102_),
    .B1(_01106_),
    .B2(_01107_),
    .ZN(_00001_));
 CLKBUF_X3 _06991_ (.A(write_data[3]),
    .Z(_01108_));
 BUF_X4 _06992_ (.A(_01108_),
    .Z(_01109_));
 NAND2_X1 _06993_ (.A1(_01109_),
    .A2(_01101_),
    .ZN(_01110_));
 NAND2_X1 _06994_ (.A1(_01105_),
    .A2(\registers[29][3] ),
    .ZN(_01111_));
 OAI21_X1 _06995_ (.A(_01110_),
    .B1(_01111_),
    .B2(_01107_),
    .ZN(_00002_));
 CLKBUF_X3 _06996_ (.A(write_data[4]),
    .Z(_01112_));
 BUF_X4 _06997_ (.A(_01112_),
    .Z(_01113_));
 NAND2_X1 _06998_ (.A1(_01113_),
    .A2(_01101_),
    .ZN(_01114_));
 NAND2_X1 _06999_ (.A1(_01105_),
    .A2(\registers[29][4] ),
    .ZN(_01115_));
 OAI21_X1 _07000_ (.A(_01114_),
    .B1(_01115_),
    .B2(_01107_),
    .ZN(_00003_));
 CLKBUF_X3 _07001_ (.A(write_data[5]),
    .Z(_01116_));
 BUF_X4 _07002_ (.A(_01116_),
    .Z(_01117_));
 NAND2_X1 _07003_ (.A1(_01117_),
    .A2(_01101_),
    .ZN(_01118_));
 NAND2_X1 _07004_ (.A1(_01105_),
    .A2(\registers[29][5] ),
    .ZN(_01119_));
 OAI21_X1 _07005_ (.A(_01118_),
    .B1(_01119_),
    .B2(_01107_),
    .ZN(_00004_));
 BUF_X4 _07006_ (.A(write_data[6]),
    .Z(_01120_));
 CLKBUF_X3 _07007_ (.A(_01120_),
    .Z(_01121_));
 NAND2_X1 _07008_ (.A1(_01121_),
    .A2(_01101_),
    .ZN(_01122_));
 NAND2_X1 _07009_ (.A1(_01105_),
    .A2(\registers[29][6] ),
    .ZN(_01123_));
 OAI21_X1 _07010_ (.A(_01122_),
    .B1(_01123_),
    .B2(_01107_),
    .ZN(_00005_));
 BUF_X4 _07011_ (.A(write_data[7]),
    .Z(_01124_));
 CLKBUF_X3 _07012_ (.A(_01124_),
    .Z(_01125_));
 NAND2_X1 _07013_ (.A1(_01125_),
    .A2(_01101_),
    .ZN(_01126_));
 NAND2_X1 _07014_ (.A1(_01105_),
    .A2(\registers[29][7] ),
    .ZN(_01127_));
 OAI21_X1 _07015_ (.A(_01126_),
    .B1(_01127_),
    .B2(_01107_),
    .ZN(_00006_));
 CLKBUF_X3 _07016_ (.A(write_data[8]),
    .Z(_01128_));
 CLKBUF_X3 _07017_ (.A(_01128_),
    .Z(_01129_));
 NAND2_X1 _07018_ (.A1(_01129_),
    .A2(_01101_),
    .ZN(_01130_));
 NAND2_X1 _07019_ (.A1(_01105_),
    .A2(\registers[29][8] ),
    .ZN(_01131_));
 OAI21_X1 _07020_ (.A(_01130_),
    .B1(_01131_),
    .B2(_01107_),
    .ZN(_00007_));
 CLKBUF_X3 _07021_ (.A(write_data[9]),
    .Z(_01132_));
 BUF_X4 _07022_ (.A(_01132_),
    .Z(_01133_));
 NAND2_X1 _07023_ (.A1(_01133_),
    .A2(_01101_),
    .ZN(_01134_));
 NAND2_X1 _07024_ (.A1(_01105_),
    .A2(\registers[29][9] ),
    .ZN(_01135_));
 OAI21_X1 _07025_ (.A(_01134_),
    .B1(_01135_),
    .B2(_01107_),
    .ZN(_00008_));
 BUF_X2 _07026_ (.A(write_data[0]),
    .Z(_01136_));
 CLKBUF_X3 _07027_ (.A(_01136_),
    .Z(_01137_));
 OR3_X1 _07028_ (.A1(net3),
    .A2(_01091_),
    .A3(_01092_),
    .ZN(_01138_));
 INV_X1 _07029_ (.A(_01096_),
    .ZN(_01139_));
 AND2_X2 _07030_ (.A1(_01095_),
    .A2(net4),
    .ZN(_01140_));
 NAND3_X4 _07031_ (.A1(_01139_),
    .A2(_01094_),
    .A3(_01140_),
    .ZN(_01141_));
 NOR2_X1 _07032_ (.A1(_01138_),
    .A2(_01141_),
    .ZN(_01142_));
 CLKBUF_X3 _07033_ (.A(_01142_),
    .Z(_01143_));
 CLKBUF_X3 _07034_ (.A(_01143_),
    .Z(_01144_));
 NAND2_X1 _07035_ (.A1(_01137_),
    .A2(_01144_),
    .ZN(_01145_));
 NAND2_X1 _07036_ (.A1(_01105_),
    .A2(\registers[2][0] ),
    .ZN(_01146_));
 CLKBUF_X3 _07037_ (.A(_01143_),
    .Z(_01147_));
 OAI21_X1 _07038_ (.A(_01145_),
    .B1(_01146_),
    .B2(_01147_),
    .ZN(_00009_));
 BUF_X2 _07039_ (.A(write_data[10]),
    .Z(_01148_));
 CLKBUF_X3 _07040_ (.A(_01148_),
    .Z(_01149_));
 NAND2_X1 _07041_ (.A1(_01149_),
    .A2(_01144_),
    .ZN(_01150_));
 NAND2_X1 _07042_ (.A1(_01105_),
    .A2(\registers[2][10] ),
    .ZN(_01151_));
 OAI21_X1 _07043_ (.A(_01150_),
    .B1(_01151_),
    .B2(_01147_),
    .ZN(_00010_));
 BUF_X2 _07044_ (.A(write_data[11]),
    .Z(_01152_));
 CLKBUF_X3 _07045_ (.A(_01152_),
    .Z(_01153_));
 NAND2_X1 _07046_ (.A1(_01153_),
    .A2(_01144_),
    .ZN(_01154_));
 CLKBUF_X3 _07047_ (.A(_01104_),
    .Z(_01155_));
 NAND2_X1 _07048_ (.A1(_01155_),
    .A2(\registers[2][11] ),
    .ZN(_01156_));
 OAI21_X1 _07049_ (.A(_01154_),
    .B1(_01156_),
    .B2(_01147_),
    .ZN(_00011_));
 BUF_X2 _07050_ (.A(write_data[12]),
    .Z(_01157_));
 CLKBUF_X3 _07051_ (.A(_01157_),
    .Z(_01158_));
 NAND2_X1 _07052_ (.A1(_01158_),
    .A2(_01144_),
    .ZN(_01159_));
 NAND2_X1 _07053_ (.A1(_01155_),
    .A2(\registers[2][12] ),
    .ZN(_01160_));
 OAI21_X1 _07054_ (.A(_01159_),
    .B1(_01160_),
    .B2(_01147_),
    .ZN(_00012_));
 BUF_X2 _07055_ (.A(write_data[13]),
    .Z(_01161_));
 BUF_X4 _07056_ (.A(_01161_),
    .Z(_01162_));
 NAND2_X1 _07057_ (.A1(_01162_),
    .A2(_01144_),
    .ZN(_01163_));
 NAND2_X1 _07058_ (.A1(_01155_),
    .A2(\registers[2][13] ),
    .ZN(_01164_));
 OAI21_X1 _07059_ (.A(_01163_),
    .B1(_01164_),
    .B2(_01147_),
    .ZN(_00013_));
 BUF_X2 _07060_ (.A(write_data[14]),
    .Z(_01165_));
 BUF_X4 _07061_ (.A(_01165_),
    .Z(_01166_));
 NAND2_X1 _07062_ (.A1(_01166_),
    .A2(_01144_),
    .ZN(_01167_));
 NAND2_X1 _07063_ (.A1(_01155_),
    .A2(\registers[2][14] ),
    .ZN(_01168_));
 OAI21_X1 _07064_ (.A(_01167_),
    .B1(_01168_),
    .B2(_01147_),
    .ZN(_00014_));
 BUF_X2 _07065_ (.A(write_data[15]),
    .Z(_01169_));
 BUF_X4 _07066_ (.A(_01169_),
    .Z(_01170_));
 NAND2_X1 _07067_ (.A1(_01170_),
    .A2(_01144_),
    .ZN(_01171_));
 NAND2_X1 _07068_ (.A1(_01155_),
    .A2(\registers[2][15] ),
    .ZN(_01172_));
 OAI21_X1 _07069_ (.A(_01171_),
    .B1(_01172_),
    .B2(_01147_),
    .ZN(_00015_));
 BUF_X2 _07070_ (.A(write_data[16]),
    .Z(_01173_));
 CLKBUF_X3 _07071_ (.A(_01173_),
    .Z(_01174_));
 NAND2_X1 _07072_ (.A1(_01174_),
    .A2(_01144_),
    .ZN(_01175_));
 NAND2_X1 _07073_ (.A1(_01155_),
    .A2(\registers[2][16] ),
    .ZN(_01176_));
 OAI21_X1 _07074_ (.A(_01175_),
    .B1(_01176_),
    .B2(_01147_),
    .ZN(_00016_));
 CLKBUF_X3 _07075_ (.A(write_data[17]),
    .Z(_01177_));
 BUF_X4 _07076_ (.A(_01177_),
    .Z(_01178_));
 CLKBUF_X3 _07077_ (.A(_01143_),
    .Z(_01179_));
 NAND2_X1 _07078_ (.A1(_01178_),
    .A2(_01179_),
    .ZN(_01180_));
 NAND2_X1 _07079_ (.A1(_01155_),
    .A2(\registers[2][17] ),
    .ZN(_01181_));
 OAI21_X1 _07080_ (.A(_01180_),
    .B1(_01181_),
    .B2(_01147_),
    .ZN(_00017_));
 CLKBUF_X3 _07081_ (.A(write_data[18]),
    .Z(_01182_));
 BUF_X4 _07082_ (.A(_01182_),
    .Z(_01183_));
 NAND2_X1 _07083_ (.A1(_01183_),
    .A2(_01179_),
    .ZN(_01184_));
 NAND2_X1 _07084_ (.A1(_01155_),
    .A2(\registers[2][18] ),
    .ZN(_01185_));
 OAI21_X1 _07085_ (.A(_01184_),
    .B1(_01185_),
    .B2(_01147_),
    .ZN(_00018_));
 BUF_X2 _07086_ (.A(write_data[19]),
    .Z(_01186_));
 CLKBUF_X3 _07087_ (.A(_01186_),
    .Z(_01187_));
 NAND2_X1 _07088_ (.A1(_01187_),
    .A2(_01179_),
    .ZN(_01188_));
 NAND2_X1 _07089_ (.A1(_01155_),
    .A2(\registers[2][19] ),
    .ZN(_01189_));
 CLKBUF_X3 _07090_ (.A(_01143_),
    .Z(_01190_));
 OAI21_X1 _07091_ (.A(_01188_),
    .B1(_01189_),
    .B2(_01190_),
    .ZN(_00019_));
 BUF_X2 _07092_ (.A(write_data[1]),
    .Z(_01191_));
 CLKBUF_X3 _07093_ (.A(_01191_),
    .Z(_01192_));
 NAND2_X1 _07094_ (.A1(_01192_),
    .A2(_01179_),
    .ZN(_01193_));
 NAND2_X1 _07095_ (.A1(_01155_),
    .A2(\registers[2][1] ),
    .ZN(_01194_));
 OAI21_X1 _07096_ (.A(_01193_),
    .B1(_01194_),
    .B2(_01190_),
    .ZN(_00020_));
 BUF_X2 _07097_ (.A(write_data[20]),
    .Z(_01195_));
 CLKBUF_X3 _07098_ (.A(_01195_),
    .Z(_01196_));
 NAND2_X1 _07099_ (.A1(_01196_),
    .A2(_01179_),
    .ZN(_01197_));
 CLKBUF_X3 _07100_ (.A(_01104_),
    .Z(_01198_));
 NAND2_X1 _07101_ (.A1(_01198_),
    .A2(\registers[2][20] ),
    .ZN(_01199_));
 OAI21_X1 _07102_ (.A(_01197_),
    .B1(_01199_),
    .B2(_01190_),
    .ZN(_00021_));
 BUF_X2 _07103_ (.A(write_data[21]),
    .Z(_01200_));
 CLKBUF_X3 _07104_ (.A(_01200_),
    .Z(_01201_));
 NAND2_X1 _07105_ (.A1(_01201_),
    .A2(_01179_),
    .ZN(_01202_));
 NAND2_X1 _07106_ (.A1(_01198_),
    .A2(\registers[2][21] ),
    .ZN(_01203_));
 OAI21_X1 _07107_ (.A(_01202_),
    .B1(_01203_),
    .B2(_01190_),
    .ZN(_00022_));
 BUF_X2 _07108_ (.A(write_data[22]),
    .Z(_01204_));
 CLKBUF_X3 _07109_ (.A(_01204_),
    .Z(_01205_));
 NAND2_X1 _07110_ (.A1(_01205_),
    .A2(_01179_),
    .ZN(_01206_));
 NAND2_X1 _07111_ (.A1(_01198_),
    .A2(\registers[2][22] ),
    .ZN(_01207_));
 OAI21_X1 _07112_ (.A(_01206_),
    .B1(_01207_),
    .B2(_01190_),
    .ZN(_00023_));
 BUF_X2 _07113_ (.A(write_data[23]),
    .Z(_01208_));
 CLKBUF_X3 _07114_ (.A(_01208_),
    .Z(_01209_));
 NAND2_X1 _07115_ (.A1(_01209_),
    .A2(_01179_),
    .ZN(_01210_));
 NAND2_X1 _07116_ (.A1(_01198_),
    .A2(\registers[2][23] ),
    .ZN(_01211_));
 OAI21_X1 _07117_ (.A(_01210_),
    .B1(_01211_),
    .B2(_01190_),
    .ZN(_00024_));
 BUF_X2 _07118_ (.A(write_data[24]),
    .Z(_01212_));
 CLKBUF_X3 _07119_ (.A(_01212_),
    .Z(_01213_));
 NAND2_X1 _07120_ (.A1(_01213_),
    .A2(_01179_),
    .ZN(_01214_));
 NAND2_X1 _07121_ (.A1(_01198_),
    .A2(\registers[2][24] ),
    .ZN(_01215_));
 OAI21_X1 _07122_ (.A(_01214_),
    .B1(_01215_),
    .B2(_01190_),
    .ZN(_00025_));
 CLKBUF_X3 _07123_ (.A(write_data[25]),
    .Z(_01216_));
 BUF_X4 _07124_ (.A(_01216_),
    .Z(_01217_));
 NAND2_X1 _07125_ (.A1(_01217_),
    .A2(_01179_),
    .ZN(_01218_));
 NAND2_X1 _07126_ (.A1(_01198_),
    .A2(\registers[2][25] ),
    .ZN(_01219_));
 OAI21_X1 _07127_ (.A(_01218_),
    .B1(_01219_),
    .B2(_01190_),
    .ZN(_00026_));
 CLKBUF_X3 _07128_ (.A(write_data[26]),
    .Z(_01220_));
 CLKBUF_X3 _07129_ (.A(_01220_),
    .Z(_01221_));
 CLKBUF_X3 _07130_ (.A(_01143_),
    .Z(_01222_));
 NAND2_X1 _07131_ (.A1(_01221_),
    .A2(_01222_),
    .ZN(_01223_));
 NAND2_X1 _07132_ (.A1(_01198_),
    .A2(\registers[2][26] ),
    .ZN(_01224_));
 OAI21_X1 _07133_ (.A(_01223_),
    .B1(_01224_),
    .B2(_01190_),
    .ZN(_00027_));
 BUF_X4 _07134_ (.A(write_data[27]),
    .Z(_01225_));
 BUF_X4 _07135_ (.A(_01225_),
    .Z(_01226_));
 NAND2_X1 _07136_ (.A1(_01226_),
    .A2(_01222_),
    .ZN(_01227_));
 NAND2_X1 _07137_ (.A1(_01198_),
    .A2(\registers[2][27] ),
    .ZN(_01228_));
 OAI21_X1 _07138_ (.A(_01227_),
    .B1(_01228_),
    .B2(_01190_),
    .ZN(_00028_));
 CLKBUF_X3 _07139_ (.A(write_data[28]),
    .Z(_01229_));
 BUF_X4 _07140_ (.A(_01229_),
    .Z(_01230_));
 NAND2_X1 _07141_ (.A1(_01230_),
    .A2(_01222_),
    .ZN(_01231_));
 NAND2_X1 _07142_ (.A1(_01198_),
    .A2(\registers[2][28] ),
    .ZN(_01232_));
 CLKBUF_X3 _07143_ (.A(_01143_),
    .Z(_01233_));
 OAI21_X1 _07144_ (.A(_01231_),
    .B1(_01232_),
    .B2(_01233_),
    .ZN(_00029_));
 CLKBUF_X3 _07145_ (.A(write_data[29]),
    .Z(_01234_));
 BUF_X4 _07146_ (.A(_01234_),
    .Z(_01235_));
 NAND2_X1 _07147_ (.A1(_01235_),
    .A2(_01222_),
    .ZN(_01236_));
 NAND2_X1 _07148_ (.A1(_01198_),
    .A2(\registers[2][29] ),
    .ZN(_01237_));
 OAI21_X1 _07149_ (.A(_01236_),
    .B1(_01237_),
    .B2(_01233_),
    .ZN(_00030_));
 BUF_X4 _07150_ (.A(write_data[2]),
    .Z(_01238_));
 BUF_X4 _07151_ (.A(_01238_),
    .Z(_01239_));
 NAND2_X1 _07152_ (.A1(_01239_),
    .A2(_01222_),
    .ZN(_01240_));
 CLKBUF_X3 _07153_ (.A(_01104_),
    .Z(_01241_));
 NAND2_X1 _07154_ (.A1(_01241_),
    .A2(\registers[2][2] ),
    .ZN(_01242_));
 OAI21_X1 _07155_ (.A(_01240_),
    .B1(_01242_),
    .B2(_01233_),
    .ZN(_00031_));
 CLKBUF_X3 _07156_ (.A(write_data[30]),
    .Z(_01243_));
 BUF_X4 _07157_ (.A(_01243_),
    .Z(_01244_));
 NAND2_X1 _07158_ (.A1(_01244_),
    .A2(_01222_),
    .ZN(_01245_));
 NAND2_X1 _07159_ (.A1(_01241_),
    .A2(\registers[2][30] ),
    .ZN(_01246_));
 OAI21_X1 _07160_ (.A(_01245_),
    .B1(_01246_),
    .B2(_01233_),
    .ZN(_00032_));
 NAND2_X1 _07161_ (.A1(_01089_),
    .A2(_01222_),
    .ZN(_01247_));
 NAND2_X1 _07162_ (.A1(_01241_),
    .A2(\registers[2][31] ),
    .ZN(_01248_));
 OAI21_X1 _07163_ (.A(_01247_),
    .B1(_01248_),
    .B2(_01233_),
    .ZN(_00033_));
 NAND2_X1 _07164_ (.A1(_01109_),
    .A2(_01222_),
    .ZN(_01249_));
 NAND2_X1 _07165_ (.A1(_01241_),
    .A2(\registers[2][3] ),
    .ZN(_01250_));
 OAI21_X1 _07166_ (.A(_01249_),
    .B1(_01250_),
    .B2(_01233_),
    .ZN(_00034_));
 NAND2_X1 _07167_ (.A1(_01113_),
    .A2(_01222_),
    .ZN(_01251_));
 NAND2_X1 _07168_ (.A1(_01241_),
    .A2(\registers[2][4] ),
    .ZN(_01252_));
 OAI21_X1 _07169_ (.A(_01251_),
    .B1(_01252_),
    .B2(_01233_),
    .ZN(_00035_));
 NAND2_X1 _07170_ (.A1(_01117_),
    .A2(_01222_),
    .ZN(_01253_));
 NAND2_X1 _07171_ (.A1(_01241_),
    .A2(\registers[2][5] ),
    .ZN(_01254_));
 OAI21_X1 _07172_ (.A(_01253_),
    .B1(_01254_),
    .B2(_01233_),
    .ZN(_00036_));
 NAND2_X1 _07173_ (.A1(_01121_),
    .A2(_01143_),
    .ZN(_01255_));
 NAND2_X1 _07174_ (.A1(_01241_),
    .A2(\registers[2][6] ),
    .ZN(_01256_));
 OAI21_X1 _07175_ (.A(_01255_),
    .B1(_01256_),
    .B2(_01233_),
    .ZN(_00037_));
 NAND2_X1 _07176_ (.A1(_01125_),
    .A2(_01143_),
    .ZN(_01257_));
 NAND2_X1 _07177_ (.A1(_01241_),
    .A2(\registers[2][7] ),
    .ZN(_01258_));
 OAI21_X1 _07178_ (.A(_01257_),
    .B1(_01258_),
    .B2(_01233_),
    .ZN(_00038_));
 NAND2_X1 _07179_ (.A1(_01129_),
    .A2(_01143_),
    .ZN(_01259_));
 NAND2_X1 _07180_ (.A1(_01241_),
    .A2(\registers[2][8] ),
    .ZN(_01260_));
 OAI21_X1 _07181_ (.A(_01259_),
    .B1(_01260_),
    .B2(_01144_),
    .ZN(_00039_));
 NAND2_X1 _07182_ (.A1(_01133_),
    .A2(_01143_),
    .ZN(_01261_));
 NAND2_X1 _07183_ (.A1(_01241_),
    .A2(\registers[2][9] ),
    .ZN(_01262_));
 OAI21_X1 _07184_ (.A(_01261_),
    .B1(_01262_),
    .B2(_01144_),
    .ZN(_00040_));
 NOR2_X1 _07185_ (.A1(_01093_),
    .A2(_01141_),
    .ZN(_01263_));
 CLKBUF_X3 _07186_ (.A(_01263_),
    .Z(_01264_));
 CLKBUF_X3 _07187_ (.A(_01264_),
    .Z(_01265_));
 NAND2_X1 _07188_ (.A1(_01137_),
    .A2(_01265_),
    .ZN(_01266_));
 BUF_X4 _07189_ (.A(_01103_),
    .Z(_01267_));
 CLKBUF_X3 _07190_ (.A(_01267_),
    .Z(_01268_));
 NAND2_X1 _07191_ (.A1(_01268_),
    .A2(\registers[30][0] ),
    .ZN(_01269_));
 CLKBUF_X3 _07192_ (.A(_01264_),
    .Z(_01270_));
 OAI21_X1 _07193_ (.A(_01266_),
    .B1(_01269_),
    .B2(_01270_),
    .ZN(_00041_));
 NAND2_X1 _07194_ (.A1(_01149_),
    .A2(_01265_),
    .ZN(_01271_));
 NAND2_X1 _07195_ (.A1(_01268_),
    .A2(\registers[30][10] ),
    .ZN(_01272_));
 OAI21_X1 _07196_ (.A(_01271_),
    .B1(_01272_),
    .B2(_01270_),
    .ZN(_00042_));
 NAND2_X1 _07197_ (.A1(_01153_),
    .A2(_01265_),
    .ZN(_01273_));
 NAND2_X1 _07198_ (.A1(_01268_),
    .A2(\registers[30][11] ),
    .ZN(_01274_));
 OAI21_X1 _07199_ (.A(_01273_),
    .B1(_01274_),
    .B2(_01270_),
    .ZN(_00043_));
 NAND2_X1 _07200_ (.A1(_01158_),
    .A2(_01265_),
    .ZN(_01275_));
 NAND2_X1 _07201_ (.A1(_01268_),
    .A2(\registers[30][12] ),
    .ZN(_01276_));
 OAI21_X1 _07202_ (.A(_01275_),
    .B1(_01276_),
    .B2(_01270_),
    .ZN(_00044_));
 NAND2_X1 _07203_ (.A1(_01162_),
    .A2(_01265_),
    .ZN(_01277_));
 NAND2_X1 _07204_ (.A1(_01268_),
    .A2(\registers[30][13] ),
    .ZN(_01278_));
 OAI21_X1 _07205_ (.A(_01277_),
    .B1(_01278_),
    .B2(_01270_),
    .ZN(_00045_));
 NAND2_X1 _07206_ (.A1(_01166_),
    .A2(_01265_),
    .ZN(_01279_));
 NAND2_X1 _07207_ (.A1(_01268_),
    .A2(\registers[30][14] ),
    .ZN(_01280_));
 OAI21_X1 _07208_ (.A(_01279_),
    .B1(_01280_),
    .B2(_01270_),
    .ZN(_00046_));
 NAND2_X1 _07209_ (.A1(_01170_),
    .A2(_01265_),
    .ZN(_01281_));
 NAND2_X1 _07210_ (.A1(_01268_),
    .A2(\registers[30][15] ),
    .ZN(_01282_));
 OAI21_X1 _07211_ (.A(_01281_),
    .B1(_01282_),
    .B2(_01270_),
    .ZN(_00047_));
 NAND2_X1 _07212_ (.A1(_01174_),
    .A2(_01265_),
    .ZN(_01283_));
 NAND2_X1 _07213_ (.A1(_01268_),
    .A2(\registers[30][16] ),
    .ZN(_01284_));
 OAI21_X1 _07214_ (.A(_01283_),
    .B1(_01284_),
    .B2(_01270_),
    .ZN(_00048_));
 CLKBUF_X3 _07215_ (.A(_01264_),
    .Z(_01285_));
 NAND2_X1 _07216_ (.A1(_01178_),
    .A2(_01285_),
    .ZN(_01286_));
 NAND2_X1 _07217_ (.A1(_01268_),
    .A2(\registers[30][17] ),
    .ZN(_01287_));
 OAI21_X1 _07218_ (.A(_01286_),
    .B1(_01287_),
    .B2(_01270_),
    .ZN(_00049_));
 NAND2_X1 _07219_ (.A1(_01183_),
    .A2(_01285_),
    .ZN(_01288_));
 NAND2_X1 _07220_ (.A1(_01268_),
    .A2(\registers[30][18] ),
    .ZN(_01289_));
 OAI21_X1 _07221_ (.A(_01288_),
    .B1(_01289_),
    .B2(_01270_),
    .ZN(_00050_));
 NAND2_X1 _07222_ (.A1(_01187_),
    .A2(_01285_),
    .ZN(_01290_));
 CLKBUF_X3 _07223_ (.A(_01267_),
    .Z(_01291_));
 NAND2_X1 _07224_ (.A1(_01291_),
    .A2(\registers[30][19] ),
    .ZN(_01292_));
 CLKBUF_X3 _07225_ (.A(_01264_),
    .Z(_01293_));
 OAI21_X1 _07226_ (.A(_01290_),
    .B1(_01292_),
    .B2(_01293_),
    .ZN(_00051_));
 NAND2_X1 _07227_ (.A1(_01192_),
    .A2(_01285_),
    .ZN(_01294_));
 NAND2_X1 _07228_ (.A1(_01291_),
    .A2(\registers[30][1] ),
    .ZN(_01295_));
 OAI21_X1 _07229_ (.A(_01294_),
    .B1(_01295_),
    .B2(_01293_),
    .ZN(_00052_));
 NAND2_X1 _07230_ (.A1(_01196_),
    .A2(_01285_),
    .ZN(_01296_));
 NAND2_X1 _07231_ (.A1(_01291_),
    .A2(\registers[30][20] ),
    .ZN(_01297_));
 OAI21_X1 _07232_ (.A(_01296_),
    .B1(_01297_),
    .B2(_01293_),
    .ZN(_00053_));
 NAND2_X1 _07233_ (.A1(_01201_),
    .A2(_01285_),
    .ZN(_01298_));
 NAND2_X1 _07234_ (.A1(_01291_),
    .A2(\registers[30][21] ),
    .ZN(_01299_));
 OAI21_X1 _07235_ (.A(_01298_),
    .B1(_01299_),
    .B2(_01293_),
    .ZN(_00054_));
 NAND2_X1 _07236_ (.A1(_01205_),
    .A2(_01285_),
    .ZN(_01300_));
 NAND2_X1 _07237_ (.A1(_01291_),
    .A2(\registers[30][22] ),
    .ZN(_01301_));
 OAI21_X1 _07238_ (.A(_01300_),
    .B1(_01301_),
    .B2(_01293_),
    .ZN(_00055_));
 NAND2_X1 _07239_ (.A1(_01209_),
    .A2(_01285_),
    .ZN(_01302_));
 NAND2_X1 _07240_ (.A1(_01291_),
    .A2(\registers[30][23] ),
    .ZN(_01303_));
 OAI21_X1 _07241_ (.A(_01302_),
    .B1(_01303_),
    .B2(_01293_),
    .ZN(_00056_));
 NAND2_X1 _07242_ (.A1(_01213_),
    .A2(_01285_),
    .ZN(_01304_));
 NAND2_X1 _07243_ (.A1(_01291_),
    .A2(\registers[30][24] ),
    .ZN(_01305_));
 OAI21_X1 _07244_ (.A(_01304_),
    .B1(_01305_),
    .B2(_01293_),
    .ZN(_00057_));
 NAND2_X1 _07245_ (.A1(_01217_),
    .A2(_01285_),
    .ZN(_01306_));
 NAND2_X1 _07246_ (.A1(_01291_),
    .A2(\registers[30][25] ),
    .ZN(_01307_));
 OAI21_X1 _07247_ (.A(_01306_),
    .B1(_01307_),
    .B2(_01293_),
    .ZN(_00058_));
 CLKBUF_X3 _07248_ (.A(_01264_),
    .Z(_01308_));
 NAND2_X1 _07249_ (.A1(_01221_),
    .A2(_01308_),
    .ZN(_01309_));
 NAND2_X1 _07250_ (.A1(_01291_),
    .A2(\registers[30][26] ),
    .ZN(_01310_));
 OAI21_X1 _07251_ (.A(_01309_),
    .B1(_01310_),
    .B2(_01293_),
    .ZN(_00059_));
 NAND2_X1 _07252_ (.A1(_01226_),
    .A2(_01308_),
    .ZN(_01311_));
 NAND2_X1 _07253_ (.A1(_01291_),
    .A2(\registers[30][27] ),
    .ZN(_01312_));
 OAI21_X1 _07254_ (.A(_01311_),
    .B1(_01312_),
    .B2(_01293_),
    .ZN(_00060_));
 NAND2_X1 _07255_ (.A1(_01230_),
    .A2(_01308_),
    .ZN(_01313_));
 CLKBUF_X3 _07256_ (.A(_01267_),
    .Z(_01314_));
 NAND2_X1 _07257_ (.A1(_01314_),
    .A2(\registers[30][28] ),
    .ZN(_01315_));
 CLKBUF_X3 _07258_ (.A(_01264_),
    .Z(_01316_));
 OAI21_X1 _07259_ (.A(_01313_),
    .B1(_01315_),
    .B2(_01316_),
    .ZN(_00061_));
 NAND2_X1 _07260_ (.A1(_01235_),
    .A2(_01308_),
    .ZN(_01317_));
 NAND2_X1 _07261_ (.A1(_01314_),
    .A2(\registers[30][29] ),
    .ZN(_01318_));
 OAI21_X1 _07262_ (.A(_01317_),
    .B1(_01318_),
    .B2(_01316_),
    .ZN(_00062_));
 NAND2_X1 _07263_ (.A1(_01239_),
    .A2(_01308_),
    .ZN(_01319_));
 NAND2_X1 _07264_ (.A1(_01314_),
    .A2(\registers[30][2] ),
    .ZN(_01320_));
 OAI21_X1 _07265_ (.A(_01319_),
    .B1(_01320_),
    .B2(_01316_),
    .ZN(_00063_));
 NAND2_X1 _07266_ (.A1(_01244_),
    .A2(_01308_),
    .ZN(_01321_));
 NAND2_X1 _07267_ (.A1(_01314_),
    .A2(\registers[30][30] ),
    .ZN(_01322_));
 OAI21_X1 _07268_ (.A(_01321_),
    .B1(_01322_),
    .B2(_01316_),
    .ZN(_00064_));
 NAND2_X1 _07269_ (.A1(_01089_),
    .A2(_01308_),
    .ZN(_01323_));
 NAND2_X1 _07270_ (.A1(_01314_),
    .A2(\registers[30][31] ),
    .ZN(_01324_));
 OAI21_X1 _07271_ (.A(_01323_),
    .B1(_01324_),
    .B2(_01316_),
    .ZN(_00065_));
 NAND2_X1 _07272_ (.A1(_01109_),
    .A2(_01308_),
    .ZN(_01325_));
 NAND2_X1 _07273_ (.A1(_01314_),
    .A2(\registers[30][3] ),
    .ZN(_01326_));
 OAI21_X1 _07274_ (.A(_01325_),
    .B1(_01326_),
    .B2(_01316_),
    .ZN(_00066_));
 NAND2_X1 _07275_ (.A1(_01113_),
    .A2(_01308_),
    .ZN(_01327_));
 NAND2_X1 _07276_ (.A1(_01314_),
    .A2(\registers[30][4] ),
    .ZN(_01328_));
 OAI21_X1 _07277_ (.A(_01327_),
    .B1(_01328_),
    .B2(_01316_),
    .ZN(_00067_));
 NAND2_X1 _07278_ (.A1(_01117_),
    .A2(_01308_),
    .ZN(_01329_));
 NAND2_X1 _07279_ (.A1(_01314_),
    .A2(\registers[30][5] ),
    .ZN(_01330_));
 OAI21_X1 _07280_ (.A(_01329_),
    .B1(_01330_),
    .B2(_01316_),
    .ZN(_00068_));
 NAND2_X1 _07281_ (.A1(_01121_),
    .A2(_01264_),
    .ZN(_01331_));
 NAND2_X1 _07282_ (.A1(_01314_),
    .A2(\registers[30][6] ),
    .ZN(_01332_));
 OAI21_X1 _07283_ (.A(_01331_),
    .B1(_01332_),
    .B2(_01316_),
    .ZN(_00069_));
 NAND2_X1 _07284_ (.A1(_01125_),
    .A2(_01264_),
    .ZN(_01333_));
 NAND2_X1 _07285_ (.A1(_01314_),
    .A2(\registers[30][7] ),
    .ZN(_01334_));
 OAI21_X1 _07286_ (.A(_01333_),
    .B1(_01334_),
    .B2(_01316_),
    .ZN(_00070_));
 NAND2_X1 _07287_ (.A1(_01129_),
    .A2(_01264_),
    .ZN(_01335_));
 CLKBUF_X3 _07288_ (.A(_01267_),
    .Z(_01336_));
 NAND2_X1 _07289_ (.A1(_01336_),
    .A2(\registers[30][8] ),
    .ZN(_01337_));
 OAI21_X1 _07290_ (.A(_01335_),
    .B1(_01337_),
    .B2(_01265_),
    .ZN(_00071_));
 NAND2_X1 _07291_ (.A1(_01133_),
    .A2(_01264_),
    .ZN(_01338_));
 NAND2_X1 _07292_ (.A1(_01336_),
    .A2(\registers[30][9] ),
    .ZN(_01339_));
 OAI21_X1 _07293_ (.A(_01338_),
    .B1(_01339_),
    .B2(_01265_),
    .ZN(_00072_));
 NAND3_X4 _07294_ (.A1(_01096_),
    .A2(_01094_),
    .A3(_01140_),
    .ZN(_01340_));
 NOR2_X1 _07295_ (.A1(_01093_),
    .A2(_01340_),
    .ZN(_01341_));
 BUF_X4 _07296_ (.A(_01341_),
    .Z(_01342_));
 BUF_X4 _07297_ (.A(_01342_),
    .Z(_01343_));
 NAND2_X1 _07298_ (.A1(_01137_),
    .A2(_01343_),
    .ZN(_01344_));
 NAND2_X1 _07299_ (.A1(_01336_),
    .A2(\registers[31][0] ),
    .ZN(_01345_));
 BUF_X4 _07300_ (.A(_01342_),
    .Z(_01346_));
 OAI21_X1 _07301_ (.A(_01344_),
    .B1(_01345_),
    .B2(_01346_),
    .ZN(_00073_));
 NAND2_X1 _07302_ (.A1(_01149_),
    .A2(_01343_),
    .ZN(_01347_));
 NAND2_X1 _07303_ (.A1(_01336_),
    .A2(\registers[31][10] ),
    .ZN(_01348_));
 OAI21_X1 _07304_ (.A(_01347_),
    .B1(_01348_),
    .B2(_01346_),
    .ZN(_00074_));
 NAND2_X1 _07305_ (.A1(_01153_),
    .A2(_01343_),
    .ZN(_01349_));
 NAND2_X1 _07306_ (.A1(_01336_),
    .A2(\registers[31][11] ),
    .ZN(_01350_));
 OAI21_X1 _07307_ (.A(_01349_),
    .B1(_01350_),
    .B2(_01346_),
    .ZN(_00075_));
 NAND2_X1 _07308_ (.A1(_01158_),
    .A2(_01343_),
    .ZN(_01351_));
 NAND2_X1 _07309_ (.A1(_01336_),
    .A2(\registers[31][12] ),
    .ZN(_01352_));
 OAI21_X1 _07310_ (.A(_01351_),
    .B1(_01352_),
    .B2(_01346_),
    .ZN(_00076_));
 NAND2_X1 _07311_ (.A1(_01162_),
    .A2(_01343_),
    .ZN(_01353_));
 NAND2_X1 _07312_ (.A1(_01336_),
    .A2(\registers[31][13] ),
    .ZN(_01354_));
 OAI21_X1 _07313_ (.A(_01353_),
    .B1(_01354_),
    .B2(_01346_),
    .ZN(_00077_));
 NAND2_X1 _07314_ (.A1(_01166_),
    .A2(_01343_),
    .ZN(_01355_));
 NAND2_X1 _07315_ (.A1(_01336_),
    .A2(\registers[31][14] ),
    .ZN(_01356_));
 OAI21_X1 _07316_ (.A(_01355_),
    .B1(_01356_),
    .B2(_01346_),
    .ZN(_00078_));
 NAND2_X1 _07317_ (.A1(_01170_),
    .A2(_01343_),
    .ZN(_01357_));
 NAND2_X1 _07318_ (.A1(_01336_),
    .A2(\registers[31][15] ),
    .ZN(_01358_));
 OAI21_X1 _07319_ (.A(_01357_),
    .B1(_01358_),
    .B2(_01346_),
    .ZN(_00079_));
 NAND2_X1 _07320_ (.A1(_01174_),
    .A2(_01343_),
    .ZN(_01359_));
 NAND2_X1 _07321_ (.A1(_01336_),
    .A2(\registers[31][16] ),
    .ZN(_01360_));
 OAI21_X1 _07322_ (.A(_01359_),
    .B1(_01360_),
    .B2(_01346_),
    .ZN(_00080_));
 CLKBUF_X3 _07323_ (.A(_01342_),
    .Z(_01361_));
 NAND2_X1 _07324_ (.A1(_01178_),
    .A2(_01361_),
    .ZN(_01362_));
 CLKBUF_X3 _07325_ (.A(_01267_),
    .Z(_01363_));
 NAND2_X1 _07326_ (.A1(_01363_),
    .A2(\registers[31][17] ),
    .ZN(_01364_));
 OAI21_X1 _07327_ (.A(_01362_),
    .B1(_01364_),
    .B2(_01346_),
    .ZN(_00081_));
 NAND2_X1 _07328_ (.A1(_01183_),
    .A2(_01361_),
    .ZN(_01365_));
 NAND2_X1 _07329_ (.A1(_01363_),
    .A2(\registers[31][18] ),
    .ZN(_01366_));
 OAI21_X1 _07330_ (.A(_01365_),
    .B1(_01366_),
    .B2(_01346_),
    .ZN(_00082_));
 NAND2_X1 _07331_ (.A1(_01187_),
    .A2(_01361_),
    .ZN(_01367_));
 NAND2_X1 _07332_ (.A1(_01363_),
    .A2(\registers[31][19] ),
    .ZN(_01368_));
 CLKBUF_X3 _07333_ (.A(_01342_),
    .Z(_01369_));
 OAI21_X1 _07334_ (.A(_01367_),
    .B1(_01368_),
    .B2(_01369_),
    .ZN(_00083_));
 NAND2_X1 _07335_ (.A1(_01192_),
    .A2(_01361_),
    .ZN(_01370_));
 NAND2_X1 _07336_ (.A1(_01363_),
    .A2(\registers[31][1] ),
    .ZN(_01371_));
 OAI21_X1 _07337_ (.A(_01370_),
    .B1(_01371_),
    .B2(_01369_),
    .ZN(_00084_));
 NAND2_X1 _07338_ (.A1(_01196_),
    .A2(_01361_),
    .ZN(_01372_));
 NAND2_X1 _07339_ (.A1(_01363_),
    .A2(\registers[31][20] ),
    .ZN(_01373_));
 OAI21_X1 _07340_ (.A(_01372_),
    .B1(_01373_),
    .B2(_01369_),
    .ZN(_00085_));
 NAND2_X1 _07341_ (.A1(_01201_),
    .A2(_01361_),
    .ZN(_01374_));
 NAND2_X1 _07342_ (.A1(_01363_),
    .A2(\registers[31][21] ),
    .ZN(_01375_));
 OAI21_X1 _07343_ (.A(_01374_),
    .B1(_01375_),
    .B2(_01369_),
    .ZN(_00086_));
 NAND2_X1 _07344_ (.A1(_01205_),
    .A2(_01361_),
    .ZN(_01376_));
 NAND2_X1 _07345_ (.A1(_01363_),
    .A2(\registers[31][22] ),
    .ZN(_01377_));
 OAI21_X1 _07346_ (.A(_01376_),
    .B1(_01377_),
    .B2(_01369_),
    .ZN(_00087_));
 NAND2_X1 _07347_ (.A1(_01209_),
    .A2(_01361_),
    .ZN(_01378_));
 NAND2_X1 _07348_ (.A1(_01363_),
    .A2(\registers[31][23] ),
    .ZN(_01379_));
 OAI21_X1 _07349_ (.A(_01378_),
    .B1(_01379_),
    .B2(_01369_),
    .ZN(_00088_));
 NAND2_X1 _07350_ (.A1(_01213_),
    .A2(_01361_),
    .ZN(_01380_));
 NAND2_X1 _07351_ (.A1(_01363_),
    .A2(\registers[31][24] ),
    .ZN(_01381_));
 OAI21_X1 _07352_ (.A(_01380_),
    .B1(_01381_),
    .B2(_01369_),
    .ZN(_00089_));
 NAND2_X1 _07353_ (.A1(_01217_),
    .A2(_01361_),
    .ZN(_01382_));
 NAND2_X1 _07354_ (.A1(_01363_),
    .A2(\registers[31][25] ),
    .ZN(_01383_));
 OAI21_X1 _07355_ (.A(_01382_),
    .B1(_01383_),
    .B2(_01369_),
    .ZN(_00090_));
 CLKBUF_X3 _07356_ (.A(_01342_),
    .Z(_01384_));
 NAND2_X1 _07357_ (.A1(_01221_),
    .A2(_01384_),
    .ZN(_01385_));
 CLKBUF_X3 _07358_ (.A(_01267_),
    .Z(_01386_));
 NAND2_X1 _07359_ (.A1(_01386_),
    .A2(\registers[31][26] ),
    .ZN(_01387_));
 OAI21_X1 _07360_ (.A(_01385_),
    .B1(_01387_),
    .B2(_01369_),
    .ZN(_00091_));
 NAND2_X1 _07361_ (.A1(_01226_),
    .A2(_01384_),
    .ZN(_01388_));
 NAND2_X1 _07362_ (.A1(_01386_),
    .A2(\registers[31][27] ),
    .ZN(_01389_));
 OAI21_X1 _07363_ (.A(_01388_),
    .B1(_01389_),
    .B2(_01369_),
    .ZN(_00092_));
 NAND2_X1 _07364_ (.A1(_01230_),
    .A2(_01384_),
    .ZN(_01390_));
 NAND2_X1 _07365_ (.A1(_01386_),
    .A2(\registers[31][28] ),
    .ZN(_01391_));
 CLKBUF_X3 _07366_ (.A(_01342_),
    .Z(_01392_));
 OAI21_X1 _07367_ (.A(_01390_),
    .B1(_01391_),
    .B2(_01392_),
    .ZN(_00093_));
 NAND2_X1 _07368_ (.A1(_01235_),
    .A2(_01384_),
    .ZN(_01393_));
 NAND2_X1 _07369_ (.A1(_01386_),
    .A2(\registers[31][29] ),
    .ZN(_01394_));
 OAI21_X1 _07370_ (.A(_01393_),
    .B1(_01394_),
    .B2(_01392_),
    .ZN(_00094_));
 NAND2_X1 _07371_ (.A1(_01239_),
    .A2(_01384_),
    .ZN(_01395_));
 NAND2_X1 _07372_ (.A1(_01386_),
    .A2(\registers[31][2] ),
    .ZN(_01396_));
 OAI21_X1 _07373_ (.A(_01395_),
    .B1(_01396_),
    .B2(_01392_),
    .ZN(_00095_));
 NAND2_X1 _07374_ (.A1(_01244_),
    .A2(_01384_),
    .ZN(_01397_));
 NAND2_X1 _07375_ (.A1(_01386_),
    .A2(\registers[31][30] ),
    .ZN(_01398_));
 OAI21_X1 _07376_ (.A(_01397_),
    .B1(_01398_),
    .B2(_01392_),
    .ZN(_00096_));
 NAND2_X1 _07377_ (.A1(_01089_),
    .A2(_01384_),
    .ZN(_01399_));
 NAND2_X1 _07378_ (.A1(_01386_),
    .A2(\registers[31][31] ),
    .ZN(_01400_));
 OAI21_X1 _07379_ (.A(_01399_),
    .B1(_01400_),
    .B2(_01392_),
    .ZN(_00097_));
 NAND2_X1 _07380_ (.A1(_01109_),
    .A2(_01384_),
    .ZN(_01401_));
 NAND2_X1 _07381_ (.A1(_01386_),
    .A2(\registers[31][3] ),
    .ZN(_01402_));
 OAI21_X1 _07382_ (.A(_01401_),
    .B1(_01402_),
    .B2(_01392_),
    .ZN(_00098_));
 NAND2_X1 _07383_ (.A1(_01113_),
    .A2(_01384_),
    .ZN(_01403_));
 NAND2_X1 _07384_ (.A1(_01386_),
    .A2(\registers[31][4] ),
    .ZN(_01404_));
 OAI21_X1 _07385_ (.A(_01403_),
    .B1(_01404_),
    .B2(_01392_),
    .ZN(_00099_));
 NAND2_X1 _07386_ (.A1(_01117_),
    .A2(_01384_),
    .ZN(_01405_));
 NAND2_X1 _07387_ (.A1(_01386_),
    .A2(\registers[31][5] ),
    .ZN(_01406_));
 OAI21_X1 _07388_ (.A(_01405_),
    .B1(_01406_),
    .B2(_01392_),
    .ZN(_00100_));
 NAND2_X1 _07389_ (.A1(_01121_),
    .A2(_01342_),
    .ZN(_01407_));
 BUF_X4 _07390_ (.A(_01267_),
    .Z(_01408_));
 NAND2_X1 _07391_ (.A1(_01408_),
    .A2(\registers[31][6] ),
    .ZN(_01409_));
 OAI21_X1 _07392_ (.A(_01407_),
    .B1(_01409_),
    .B2(_01392_),
    .ZN(_00101_));
 NAND2_X1 _07393_ (.A1(_01125_),
    .A2(_01342_),
    .ZN(_01410_));
 NAND2_X1 _07394_ (.A1(_01408_),
    .A2(\registers[31][7] ),
    .ZN(_01411_));
 OAI21_X1 _07395_ (.A(_01410_),
    .B1(_01411_),
    .B2(_01392_),
    .ZN(_00102_));
 NAND2_X1 _07396_ (.A1(_01129_),
    .A2(_01342_),
    .ZN(_01412_));
 NAND2_X1 _07397_ (.A1(_01408_),
    .A2(\registers[31][8] ),
    .ZN(_01413_));
 OAI21_X1 _07398_ (.A(_01412_),
    .B1(_01413_),
    .B2(_01343_),
    .ZN(_00103_));
 NAND2_X1 _07399_ (.A1(_01133_),
    .A2(_01342_),
    .ZN(_01414_));
 NAND2_X1 _07400_ (.A1(_01408_),
    .A2(\registers[31][9] ),
    .ZN(_01415_));
 OAI21_X1 _07401_ (.A(_01414_),
    .B1(_01415_),
    .B2(_01343_),
    .ZN(_00104_));
 BUF_X4 _07402_ (.A(_01103_),
    .Z(_01416_));
 BUF_X4 _07403_ (.A(_01416_),
    .Z(_01417_));
 CLKBUF_X3 _07404_ (.A(_01417_),
    .Z(_01418_));
 OR2_X1 _07405_ (.A1(_01138_),
    .A2(_01340_),
    .ZN(_01419_));
 CLKBUF_X3 _07406_ (.A(_01419_),
    .Z(_01420_));
 CLKBUF_X3 _07407_ (.A(_01420_),
    .Z(_01421_));
 NAND3_X1 _07408_ (.A1(_01418_),
    .A2(\registers[3][0] ),
    .A3(_01421_),
    .ZN(_01422_));
 CLKBUF_X3 _07409_ (.A(_01420_),
    .Z(_01423_));
 INV_X4 _07410_ (.A(_01136_),
    .ZN(_01424_));
 OAI21_X1 _07411_ (.A(_01422_),
    .B1(_01423_),
    .B2(_01424_),
    .ZN(_00105_));
 NAND3_X1 _07412_ (.A1(_01418_),
    .A2(\registers[3][10] ),
    .A3(_01421_),
    .ZN(_01425_));
 INV_X4 _07413_ (.A(_01148_),
    .ZN(_01426_));
 OAI21_X1 _07414_ (.A(_01425_),
    .B1(_01423_),
    .B2(_01426_),
    .ZN(_00106_));
 NAND3_X1 _07415_ (.A1(_01418_),
    .A2(\registers[3][11] ),
    .A3(_01421_),
    .ZN(_01427_));
 INV_X4 _07416_ (.A(_01152_),
    .ZN(_01428_));
 OAI21_X1 _07417_ (.A(_01427_),
    .B1(_01423_),
    .B2(_01428_),
    .ZN(_00107_));
 NAND3_X1 _07418_ (.A1(_01418_),
    .A2(\registers[3][12] ),
    .A3(_01421_),
    .ZN(_01429_));
 INV_X4 _07419_ (.A(_01157_),
    .ZN(_01430_));
 OAI21_X1 _07420_ (.A(_01429_),
    .B1(_01423_),
    .B2(_01430_),
    .ZN(_00108_));
 NAND3_X1 _07421_ (.A1(_01418_),
    .A2(\registers[3][13] ),
    .A3(_01421_),
    .ZN(_01431_));
 INV_X4 _07422_ (.A(_01161_),
    .ZN(_01432_));
 OAI21_X1 _07423_ (.A(_01431_),
    .B1(_01423_),
    .B2(_01432_),
    .ZN(_00109_));
 NAND3_X1 _07424_ (.A1(_01418_),
    .A2(\registers[3][14] ),
    .A3(_01421_),
    .ZN(_01433_));
 INV_X4 _07425_ (.A(_01165_),
    .ZN(_01434_));
 OAI21_X1 _07426_ (.A(_01433_),
    .B1(_01423_),
    .B2(_01434_),
    .ZN(_00110_));
 NAND3_X1 _07427_ (.A1(_01418_),
    .A2(\registers[3][15] ),
    .A3(_01421_),
    .ZN(_01435_));
 INV_X4 _07428_ (.A(_01169_),
    .ZN(_01436_));
 OAI21_X1 _07429_ (.A(_01435_),
    .B1(_01423_),
    .B2(_01436_),
    .ZN(_00111_));
 NAND3_X1 _07430_ (.A1(_01418_),
    .A2(\registers[3][16] ),
    .A3(_01421_),
    .ZN(_01437_));
 INV_X4 _07431_ (.A(_01173_),
    .ZN(_01438_));
 OAI21_X1 _07432_ (.A(_01437_),
    .B1(_01423_),
    .B2(_01438_),
    .ZN(_00112_));
 CLKBUF_X3 _07433_ (.A(_01420_),
    .Z(_01439_));
 NAND3_X1 _07434_ (.A1(_01418_),
    .A2(\registers[3][17] ),
    .A3(_01439_),
    .ZN(_01440_));
 INV_X4 _07435_ (.A(_01177_),
    .ZN(_01441_));
 OAI21_X1 _07436_ (.A(_01440_),
    .B1(_01423_),
    .B2(_01441_),
    .ZN(_00113_));
 NAND3_X1 _07437_ (.A1(_01418_),
    .A2(\registers[3][18] ),
    .A3(_01439_),
    .ZN(_01442_));
 INV_X4 _07438_ (.A(_01182_),
    .ZN(_01443_));
 OAI21_X1 _07439_ (.A(_01442_),
    .B1(_01423_),
    .B2(_01443_),
    .ZN(_00114_));
 CLKBUF_X3 _07440_ (.A(_01417_),
    .Z(_01444_));
 NAND3_X1 _07441_ (.A1(_01444_),
    .A2(\registers[3][19] ),
    .A3(_01439_),
    .ZN(_01445_));
 CLKBUF_X3 _07442_ (.A(_01420_),
    .Z(_01446_));
 INV_X4 _07443_ (.A(_01186_),
    .ZN(_01447_));
 OAI21_X1 _07444_ (.A(_01445_),
    .B1(_01446_),
    .B2(_01447_),
    .ZN(_00115_));
 NAND3_X1 _07445_ (.A1(_01444_),
    .A2(\registers[3][1] ),
    .A3(_01439_),
    .ZN(_01448_));
 INV_X4 _07446_ (.A(_01191_),
    .ZN(_01449_));
 OAI21_X1 _07447_ (.A(_01448_),
    .B1(_01446_),
    .B2(_01449_),
    .ZN(_00116_));
 NAND3_X1 _07448_ (.A1(_01444_),
    .A2(\registers[3][20] ),
    .A3(_01439_),
    .ZN(_01450_));
 INV_X4 _07449_ (.A(_01195_),
    .ZN(_01451_));
 OAI21_X1 _07450_ (.A(_01450_),
    .B1(_01446_),
    .B2(_01451_),
    .ZN(_00117_));
 NAND3_X1 _07451_ (.A1(_01444_),
    .A2(\registers[3][21] ),
    .A3(_01439_),
    .ZN(_01452_));
 INV_X4 _07452_ (.A(_01200_),
    .ZN(_01453_));
 OAI21_X1 _07453_ (.A(_01452_),
    .B1(_01446_),
    .B2(_01453_),
    .ZN(_00118_));
 NAND3_X1 _07454_ (.A1(_01444_),
    .A2(\registers[3][22] ),
    .A3(_01439_),
    .ZN(_01454_));
 INV_X4 _07455_ (.A(_01204_),
    .ZN(_01455_));
 OAI21_X1 _07456_ (.A(_01454_),
    .B1(_01446_),
    .B2(_01455_),
    .ZN(_00119_));
 NAND3_X1 _07457_ (.A1(_01444_),
    .A2(\registers[3][23] ),
    .A3(_01439_),
    .ZN(_01456_));
 INV_X4 _07458_ (.A(_01208_),
    .ZN(_01457_));
 OAI21_X1 _07459_ (.A(_01456_),
    .B1(_01446_),
    .B2(_01457_),
    .ZN(_00120_));
 NAND3_X1 _07460_ (.A1(_01444_),
    .A2(\registers[3][24] ),
    .A3(_01439_),
    .ZN(_01458_));
 INV_X4 _07461_ (.A(_01212_),
    .ZN(_01459_));
 OAI21_X1 _07462_ (.A(_01458_),
    .B1(_01446_),
    .B2(_01459_),
    .ZN(_00121_));
 NAND3_X1 _07463_ (.A1(_01444_),
    .A2(\registers[3][25] ),
    .A3(_01439_),
    .ZN(_01460_));
 INV_X4 _07464_ (.A(_01216_),
    .ZN(_01461_));
 OAI21_X1 _07465_ (.A(_01460_),
    .B1(_01446_),
    .B2(_01461_),
    .ZN(_00122_));
 CLKBUF_X3 _07466_ (.A(_01420_),
    .Z(_01462_));
 NAND3_X1 _07467_ (.A1(_01444_),
    .A2(\registers[3][26] ),
    .A3(_01462_),
    .ZN(_01463_));
 INV_X4 _07468_ (.A(_01220_),
    .ZN(_01464_));
 OAI21_X1 _07469_ (.A(_01463_),
    .B1(_01446_),
    .B2(_01464_),
    .ZN(_00123_));
 NAND3_X1 _07470_ (.A1(_01444_),
    .A2(\registers[3][27] ),
    .A3(_01462_),
    .ZN(_01465_));
 INV_X4 _07471_ (.A(_01225_),
    .ZN(_01466_));
 OAI21_X1 _07472_ (.A(_01465_),
    .B1(_01446_),
    .B2(_01466_),
    .ZN(_00124_));
 CLKBUF_X3 _07473_ (.A(_01417_),
    .Z(_01467_));
 NAND3_X1 _07474_ (.A1(_01467_),
    .A2(\registers[3][28] ),
    .A3(_01462_),
    .ZN(_01468_));
 CLKBUF_X3 _07475_ (.A(_01420_),
    .Z(_01469_));
 INV_X4 _07476_ (.A(_01229_),
    .ZN(_01470_));
 OAI21_X1 _07477_ (.A(_01468_),
    .B1(_01469_),
    .B2(_01470_),
    .ZN(_00125_));
 NAND3_X1 _07478_ (.A1(_01467_),
    .A2(\registers[3][29] ),
    .A3(_01462_),
    .ZN(_01471_));
 INV_X4 _07479_ (.A(_01234_),
    .ZN(_01472_));
 OAI21_X1 _07480_ (.A(_01471_),
    .B1(_01469_),
    .B2(_01472_),
    .ZN(_00126_));
 NAND3_X1 _07481_ (.A1(_01467_),
    .A2(\registers[3][2] ),
    .A3(_01462_),
    .ZN(_01473_));
 INV_X4 _07482_ (.A(_01238_),
    .ZN(_01474_));
 OAI21_X1 _07483_ (.A(_01473_),
    .B1(_01469_),
    .B2(_01474_),
    .ZN(_00127_));
 NAND3_X1 _07484_ (.A1(_01467_),
    .A2(\registers[3][30] ),
    .A3(_01462_),
    .ZN(_01475_));
 INV_X4 _07485_ (.A(_01243_),
    .ZN(_01476_));
 OAI21_X1 _07486_ (.A(_01475_),
    .B1(_01469_),
    .B2(_01476_),
    .ZN(_00128_));
 NAND3_X1 _07487_ (.A1(_01467_),
    .A2(\registers[3][31] ),
    .A3(_01462_),
    .ZN(_01477_));
 INV_X4 _07488_ (.A(_01088_),
    .ZN(_01478_));
 OAI21_X1 _07489_ (.A(_01477_),
    .B1(_01469_),
    .B2(_01478_),
    .ZN(_00129_));
 NAND3_X1 _07490_ (.A1(_01467_),
    .A2(\registers[3][3] ),
    .A3(_01462_),
    .ZN(_01479_));
 INV_X4 _07491_ (.A(_01108_),
    .ZN(_01480_));
 OAI21_X1 _07492_ (.A(_01479_),
    .B1(_01469_),
    .B2(_01480_),
    .ZN(_00130_));
 NAND3_X1 _07493_ (.A1(_01467_),
    .A2(\registers[3][4] ),
    .A3(_01462_),
    .ZN(_01481_));
 INV_X4 _07494_ (.A(_01112_),
    .ZN(_01482_));
 OAI21_X1 _07495_ (.A(_01481_),
    .B1(_01469_),
    .B2(_01482_),
    .ZN(_00131_));
 NAND3_X1 _07496_ (.A1(_01467_),
    .A2(\registers[3][5] ),
    .A3(_01462_),
    .ZN(_01483_));
 INV_X4 _07497_ (.A(_01116_),
    .ZN(_01484_));
 OAI21_X1 _07498_ (.A(_01483_),
    .B1(_01469_),
    .B2(_01484_),
    .ZN(_00132_));
 NAND3_X1 _07499_ (.A1(_01467_),
    .A2(\registers[3][6] ),
    .A3(_01420_),
    .ZN(_01485_));
 INV_X4 _07500_ (.A(_01120_),
    .ZN(_01486_));
 OAI21_X1 _07501_ (.A(_01485_),
    .B1(_01469_),
    .B2(_01486_),
    .ZN(_00133_));
 NAND3_X1 _07502_ (.A1(_01467_),
    .A2(\registers[3][7] ),
    .A3(_01420_),
    .ZN(_01487_));
 INV_X4 _07503_ (.A(_01124_),
    .ZN(_01488_));
 OAI21_X1 _07504_ (.A(_01487_),
    .B1(_01469_),
    .B2(_01488_),
    .ZN(_00134_));
 CLKBUF_X3 _07505_ (.A(_01417_),
    .Z(_01489_));
 NAND3_X1 _07506_ (.A1(_01489_),
    .A2(\registers[3][8] ),
    .A3(_01420_),
    .ZN(_01490_));
 INV_X4 _07507_ (.A(_01128_),
    .ZN(_01491_));
 OAI21_X1 _07508_ (.A(_01490_),
    .B1(_01421_),
    .B2(_01491_),
    .ZN(_00135_));
 NAND3_X1 _07509_ (.A1(_01489_),
    .A2(\registers[3][9] ),
    .A3(_01420_),
    .ZN(_01492_));
 INV_X4 _07510_ (.A(_01132_),
    .ZN(_01493_));
 OAI21_X1 _07511_ (.A(_01492_),
    .B1(_01421_),
    .B2(_01493_),
    .ZN(_00136_));
 INV_X2 _07512_ (.A(_01092_),
    .ZN(_01494_));
 NOR3_X1 _07513_ (.A1(_01090_),
    .A2(_01091_),
    .A3(_01494_),
    .ZN(_01495_));
 NAND2_X1 _07514_ (.A1(_01095_),
    .A2(net4),
    .ZN(_01496_));
 NOR3_X1 _07515_ (.A1(_01096_),
    .A2(_01094_),
    .A3(_01496_),
    .ZN(_01497_));
 NAND2_X1 _07516_ (.A1(_01495_),
    .A2(_01497_),
    .ZN(_01498_));
 CLKBUF_X3 _07517_ (.A(_01498_),
    .Z(_01499_));
 CLKBUF_X3 _07518_ (.A(_01499_),
    .Z(_01500_));
 NAND3_X1 _07519_ (.A1(_01489_),
    .A2(\registers[4][0] ),
    .A3(_01500_),
    .ZN(_01501_));
 CLKBUF_X3 _07520_ (.A(_01499_),
    .Z(_01502_));
 OAI21_X1 _07521_ (.A(_01501_),
    .B1(_01502_),
    .B2(_01424_),
    .ZN(_00137_));
 NAND3_X1 _07522_ (.A1(_01489_),
    .A2(\registers[4][10] ),
    .A3(_01500_),
    .ZN(_01503_));
 OAI21_X1 _07523_ (.A(_01503_),
    .B1(_01502_),
    .B2(_01426_),
    .ZN(_00138_));
 NAND3_X1 _07524_ (.A1(_01489_),
    .A2(\registers[4][11] ),
    .A3(_01500_),
    .ZN(_01504_));
 OAI21_X1 _07525_ (.A(_01504_),
    .B1(_01502_),
    .B2(_01428_),
    .ZN(_00139_));
 NAND3_X1 _07526_ (.A1(_01489_),
    .A2(\registers[4][12] ),
    .A3(_01500_),
    .ZN(_01505_));
 OAI21_X1 _07527_ (.A(_01505_),
    .B1(_01502_),
    .B2(_01430_),
    .ZN(_00140_));
 NAND3_X1 _07528_ (.A1(_01489_),
    .A2(\registers[4][13] ),
    .A3(_01500_),
    .ZN(_01506_));
 OAI21_X1 _07529_ (.A(_01506_),
    .B1(_01502_),
    .B2(_01432_),
    .ZN(_00141_));
 NAND3_X1 _07530_ (.A1(_01489_),
    .A2(\registers[4][14] ),
    .A3(_01500_),
    .ZN(_01507_));
 OAI21_X1 _07531_ (.A(_01507_),
    .B1(_01502_),
    .B2(_01434_),
    .ZN(_00142_));
 NAND3_X1 _07532_ (.A1(_01489_),
    .A2(\registers[4][15] ),
    .A3(_01500_),
    .ZN(_01508_));
 OAI21_X1 _07533_ (.A(_01508_),
    .B1(_01502_),
    .B2(_01436_),
    .ZN(_00143_));
 NAND3_X1 _07534_ (.A1(_01489_),
    .A2(\registers[4][16] ),
    .A3(_01500_),
    .ZN(_01509_));
 OAI21_X1 _07535_ (.A(_01509_),
    .B1(_01502_),
    .B2(_01438_),
    .ZN(_00144_));
 CLKBUF_X3 _07536_ (.A(_01417_),
    .Z(_01510_));
 CLKBUF_X3 _07537_ (.A(_01499_),
    .Z(_01511_));
 NAND3_X1 _07538_ (.A1(_01510_),
    .A2(\registers[4][17] ),
    .A3(_01511_),
    .ZN(_01512_));
 OAI21_X1 _07539_ (.A(_01512_),
    .B1(_01502_),
    .B2(_01441_),
    .ZN(_00145_));
 NAND3_X1 _07540_ (.A1(_01510_),
    .A2(\registers[4][18] ),
    .A3(_01511_),
    .ZN(_01513_));
 OAI21_X1 _07541_ (.A(_01513_),
    .B1(_01502_),
    .B2(_01443_),
    .ZN(_00146_));
 NAND3_X1 _07542_ (.A1(_01510_),
    .A2(\registers[4][19] ),
    .A3(_01511_),
    .ZN(_01514_));
 CLKBUF_X3 _07543_ (.A(_01499_),
    .Z(_01515_));
 OAI21_X1 _07544_ (.A(_01514_),
    .B1(_01515_),
    .B2(_01447_),
    .ZN(_00147_));
 NAND3_X1 _07545_ (.A1(_01510_),
    .A2(\registers[4][1] ),
    .A3(_01511_),
    .ZN(_01516_));
 OAI21_X1 _07546_ (.A(_01516_),
    .B1(_01515_),
    .B2(_01449_),
    .ZN(_00148_));
 NAND3_X1 _07547_ (.A1(_01510_),
    .A2(\registers[4][20] ),
    .A3(_01511_),
    .ZN(_01517_));
 OAI21_X1 _07548_ (.A(_01517_),
    .B1(_01515_),
    .B2(_01451_),
    .ZN(_00149_));
 NAND3_X1 _07549_ (.A1(_01510_),
    .A2(\registers[4][21] ),
    .A3(_01511_),
    .ZN(_01518_));
 OAI21_X1 _07550_ (.A(_01518_),
    .B1(_01515_),
    .B2(_01453_),
    .ZN(_00150_));
 NAND3_X1 _07551_ (.A1(_01510_),
    .A2(\registers[4][22] ),
    .A3(_01511_),
    .ZN(_01519_));
 OAI21_X1 _07552_ (.A(_01519_),
    .B1(_01515_),
    .B2(_01455_),
    .ZN(_00151_));
 NAND3_X1 _07553_ (.A1(_01510_),
    .A2(\registers[4][23] ),
    .A3(_01511_),
    .ZN(_01520_));
 OAI21_X1 _07554_ (.A(_01520_),
    .B1(_01515_),
    .B2(_01457_),
    .ZN(_00152_));
 NAND3_X1 _07555_ (.A1(_01510_),
    .A2(\registers[4][24] ),
    .A3(_01511_),
    .ZN(_01521_));
 OAI21_X1 _07556_ (.A(_01521_),
    .B1(_01515_),
    .B2(_01459_),
    .ZN(_00153_));
 NAND3_X1 _07557_ (.A1(_01510_),
    .A2(\registers[4][25] ),
    .A3(_01511_),
    .ZN(_01522_));
 OAI21_X1 _07558_ (.A(_01522_),
    .B1(_01515_),
    .B2(_01461_),
    .ZN(_00154_));
 CLKBUF_X3 _07559_ (.A(_01417_),
    .Z(_01523_));
 CLKBUF_X3 _07560_ (.A(_01499_),
    .Z(_01524_));
 NAND3_X1 _07561_ (.A1(_01523_),
    .A2(\registers[4][26] ),
    .A3(_01524_),
    .ZN(_01525_));
 OAI21_X1 _07562_ (.A(_01525_),
    .B1(_01515_),
    .B2(_01464_),
    .ZN(_00155_));
 NAND3_X1 _07563_ (.A1(_01523_),
    .A2(\registers[4][27] ),
    .A3(_01524_),
    .ZN(_01526_));
 OAI21_X1 _07564_ (.A(_01526_),
    .B1(_01515_),
    .B2(_01466_),
    .ZN(_00156_));
 NAND3_X1 _07565_ (.A1(_01523_),
    .A2(\registers[4][28] ),
    .A3(_01524_),
    .ZN(_01527_));
 CLKBUF_X3 _07566_ (.A(_01499_),
    .Z(_01528_));
 OAI21_X1 _07567_ (.A(_01527_),
    .B1(_01528_),
    .B2(_01470_),
    .ZN(_00157_));
 NAND3_X1 _07568_ (.A1(_01523_),
    .A2(\registers[4][29] ),
    .A3(_01524_),
    .ZN(_01529_));
 OAI21_X1 _07569_ (.A(_01529_),
    .B1(_01528_),
    .B2(_01472_),
    .ZN(_00158_));
 NAND3_X1 _07570_ (.A1(_01523_),
    .A2(\registers[4][2] ),
    .A3(_01524_),
    .ZN(_01530_));
 OAI21_X1 _07571_ (.A(_01530_),
    .B1(_01528_),
    .B2(_01474_),
    .ZN(_00159_));
 NAND3_X1 _07572_ (.A1(_01523_),
    .A2(\registers[4][30] ),
    .A3(_01524_),
    .ZN(_01531_));
 OAI21_X1 _07573_ (.A(_01531_),
    .B1(_01528_),
    .B2(_01476_),
    .ZN(_00160_));
 NAND3_X1 _07574_ (.A1(_01523_),
    .A2(\registers[4][31] ),
    .A3(_01524_),
    .ZN(_01532_));
 OAI21_X1 _07575_ (.A(_01532_),
    .B1(_01528_),
    .B2(_01478_),
    .ZN(_00161_));
 NAND3_X1 _07576_ (.A1(_01523_),
    .A2(\registers[4][3] ),
    .A3(_01524_),
    .ZN(_01533_));
 OAI21_X1 _07577_ (.A(_01533_),
    .B1(_01528_),
    .B2(_01480_),
    .ZN(_00162_));
 NAND3_X1 _07578_ (.A1(_01523_),
    .A2(\registers[4][4] ),
    .A3(_01524_),
    .ZN(_01534_));
 OAI21_X1 _07579_ (.A(_01534_),
    .B1(_01528_),
    .B2(_01482_),
    .ZN(_00163_));
 NAND3_X1 _07580_ (.A1(_01523_),
    .A2(\registers[4][5] ),
    .A3(_01524_),
    .ZN(_01535_));
 OAI21_X1 _07581_ (.A(_01535_),
    .B1(_01528_),
    .B2(_01484_),
    .ZN(_00164_));
 BUF_X4 _07582_ (.A(_01416_),
    .Z(_01536_));
 BUF_X4 _07583_ (.A(_01536_),
    .Z(_01537_));
 NAND3_X1 _07584_ (.A1(_01537_),
    .A2(\registers[4][6] ),
    .A3(_01499_),
    .ZN(_01538_));
 OAI21_X1 _07585_ (.A(_01538_),
    .B1(_01528_),
    .B2(_01486_),
    .ZN(_00165_));
 NAND3_X1 _07586_ (.A1(_01537_),
    .A2(\registers[4][7] ),
    .A3(_01499_),
    .ZN(_01539_));
 OAI21_X1 _07587_ (.A(_01539_),
    .B1(_01528_),
    .B2(_01488_),
    .ZN(_00166_));
 NAND3_X1 _07588_ (.A1(_01537_),
    .A2(\registers[4][8] ),
    .A3(_01499_),
    .ZN(_01540_));
 OAI21_X1 _07589_ (.A(_01540_),
    .B1(_01500_),
    .B2(_01491_),
    .ZN(_00167_));
 NAND3_X1 _07590_ (.A1(_01537_),
    .A2(\registers[4][9] ),
    .A3(_01499_),
    .ZN(_01541_));
 OAI21_X1 _07591_ (.A(_01541_),
    .B1(_01500_),
    .B2(_01493_),
    .ZN(_00168_));
 NOR2_X1 _07592_ (.A1(_01094_),
    .A2(_01097_),
    .ZN(_01542_));
 NAND2_X1 _07593_ (.A1(_01542_),
    .A2(_01495_),
    .ZN(_01543_));
 CLKBUF_X3 _07594_ (.A(_01543_),
    .Z(_01544_));
 CLKBUF_X3 _07595_ (.A(_01544_),
    .Z(_01545_));
 NAND3_X1 _07596_ (.A1(_01537_),
    .A2(\registers[5][0] ),
    .A3(_01545_),
    .ZN(_01546_));
 CLKBUF_X3 _07597_ (.A(_01544_),
    .Z(_01547_));
 OAI21_X1 _07598_ (.A(_01546_),
    .B1(_01547_),
    .B2(_01424_),
    .ZN(_00169_));
 NAND3_X1 _07599_ (.A1(_01537_),
    .A2(\registers[5][10] ),
    .A3(_01545_),
    .ZN(_01548_));
 OAI21_X1 _07600_ (.A(_01548_),
    .B1(_01547_),
    .B2(_01426_),
    .ZN(_00170_));
 NAND3_X1 _07601_ (.A1(_01537_),
    .A2(\registers[5][11] ),
    .A3(_01545_),
    .ZN(_01549_));
 OAI21_X1 _07602_ (.A(_01549_),
    .B1(_01547_),
    .B2(_01428_),
    .ZN(_00171_));
 NAND3_X1 _07603_ (.A1(_01537_),
    .A2(\registers[5][12] ),
    .A3(_01545_),
    .ZN(_01550_));
 OAI21_X1 _07604_ (.A(_01550_),
    .B1(_01547_),
    .B2(_01430_),
    .ZN(_00172_));
 NAND3_X1 _07605_ (.A1(_01537_),
    .A2(\registers[5][13] ),
    .A3(_01545_),
    .ZN(_01551_));
 OAI21_X1 _07606_ (.A(_01551_),
    .B1(_01547_),
    .B2(_01432_),
    .ZN(_00173_));
 NAND3_X1 _07607_ (.A1(_01537_),
    .A2(\registers[5][14] ),
    .A3(_01545_),
    .ZN(_01552_));
 OAI21_X1 _07608_ (.A(_01552_),
    .B1(_01547_),
    .B2(_01434_),
    .ZN(_00174_));
 CLKBUF_X3 _07609_ (.A(_01536_),
    .Z(_01553_));
 NAND3_X1 _07610_ (.A1(_01553_),
    .A2(\registers[5][15] ),
    .A3(_01545_),
    .ZN(_01554_));
 OAI21_X1 _07611_ (.A(_01554_),
    .B1(_01547_),
    .B2(_01436_),
    .ZN(_00175_));
 NAND3_X1 _07612_ (.A1(_01553_),
    .A2(\registers[5][16] ),
    .A3(_01545_),
    .ZN(_01555_));
 OAI21_X1 _07613_ (.A(_01555_),
    .B1(_01547_),
    .B2(_01438_),
    .ZN(_00176_));
 CLKBUF_X3 _07614_ (.A(_01544_),
    .Z(_01556_));
 NAND3_X1 _07615_ (.A1(_01553_),
    .A2(\registers[5][17] ),
    .A3(_01556_),
    .ZN(_01557_));
 OAI21_X1 _07616_ (.A(_01557_),
    .B1(_01547_),
    .B2(_01441_),
    .ZN(_00177_));
 NAND3_X1 _07617_ (.A1(_01553_),
    .A2(\registers[5][18] ),
    .A3(_01556_),
    .ZN(_01558_));
 OAI21_X1 _07618_ (.A(_01558_),
    .B1(_01547_),
    .B2(_01443_),
    .ZN(_00178_));
 NAND3_X1 _07619_ (.A1(_01553_),
    .A2(\registers[5][19] ),
    .A3(_01556_),
    .ZN(_01559_));
 CLKBUF_X3 _07620_ (.A(_01544_),
    .Z(_01560_));
 OAI21_X1 _07621_ (.A(_01559_),
    .B1(_01560_),
    .B2(_01447_),
    .ZN(_00179_));
 NAND3_X1 _07622_ (.A1(_01553_),
    .A2(\registers[5][1] ),
    .A3(_01556_),
    .ZN(_01561_));
 OAI21_X1 _07623_ (.A(_01561_),
    .B1(_01560_),
    .B2(_01449_),
    .ZN(_00180_));
 NAND3_X1 _07624_ (.A1(_01553_),
    .A2(\registers[5][20] ),
    .A3(_01556_),
    .ZN(_01562_));
 OAI21_X1 _07625_ (.A(_01562_),
    .B1(_01560_),
    .B2(_01451_),
    .ZN(_00181_));
 NAND3_X1 _07626_ (.A1(_01553_),
    .A2(\registers[5][21] ),
    .A3(_01556_),
    .ZN(_01563_));
 OAI21_X1 _07627_ (.A(_01563_),
    .B1(_01560_),
    .B2(_01453_),
    .ZN(_00182_));
 NAND3_X1 _07628_ (.A1(_01553_),
    .A2(\registers[5][22] ),
    .A3(_01556_),
    .ZN(_01564_));
 OAI21_X1 _07629_ (.A(_01564_),
    .B1(_01560_),
    .B2(_01455_),
    .ZN(_00183_));
 NAND3_X1 _07630_ (.A1(_01553_),
    .A2(\registers[5][23] ),
    .A3(_01556_),
    .ZN(_01565_));
 OAI21_X1 _07631_ (.A(_01565_),
    .B1(_01560_),
    .B2(_01457_),
    .ZN(_00184_));
 CLKBUF_X3 _07632_ (.A(_01536_),
    .Z(_01566_));
 NAND3_X1 _07633_ (.A1(_01566_),
    .A2(\registers[5][24] ),
    .A3(_01556_),
    .ZN(_01567_));
 OAI21_X1 _07634_ (.A(_01567_),
    .B1(_01560_),
    .B2(_01459_),
    .ZN(_00185_));
 NAND3_X1 _07635_ (.A1(_01566_),
    .A2(\registers[5][25] ),
    .A3(_01556_),
    .ZN(_01568_));
 OAI21_X1 _07636_ (.A(_01568_),
    .B1(_01560_),
    .B2(_01461_),
    .ZN(_00186_));
 CLKBUF_X3 _07637_ (.A(_01544_),
    .Z(_01569_));
 NAND3_X1 _07638_ (.A1(_01566_),
    .A2(\registers[5][26] ),
    .A3(_01569_),
    .ZN(_01570_));
 OAI21_X1 _07639_ (.A(_01570_),
    .B1(_01560_),
    .B2(_01464_),
    .ZN(_00187_));
 NAND3_X1 _07640_ (.A1(_01566_),
    .A2(\registers[5][27] ),
    .A3(_01569_),
    .ZN(_01571_));
 OAI21_X1 _07641_ (.A(_01571_),
    .B1(_01560_),
    .B2(_01466_),
    .ZN(_00188_));
 NAND3_X1 _07642_ (.A1(_01566_),
    .A2(\registers[5][28] ),
    .A3(_01569_),
    .ZN(_01572_));
 CLKBUF_X3 _07643_ (.A(_01544_),
    .Z(_01573_));
 OAI21_X1 _07644_ (.A(_01572_),
    .B1(_01573_),
    .B2(_01470_),
    .ZN(_00189_));
 NAND3_X1 _07645_ (.A1(_01566_),
    .A2(\registers[5][29] ),
    .A3(_01569_),
    .ZN(_01574_));
 OAI21_X1 _07646_ (.A(_01574_),
    .B1(_01573_),
    .B2(_01472_),
    .ZN(_00190_));
 NAND3_X1 _07647_ (.A1(_01566_),
    .A2(\registers[5][2] ),
    .A3(_01569_),
    .ZN(_01575_));
 OAI21_X1 _07648_ (.A(_01575_),
    .B1(_01573_),
    .B2(_01474_),
    .ZN(_00191_));
 NAND3_X1 _07649_ (.A1(_01566_),
    .A2(\registers[5][30] ),
    .A3(_01569_),
    .ZN(_01576_));
 OAI21_X1 _07650_ (.A(_01576_),
    .B1(_01573_),
    .B2(_01476_),
    .ZN(_00192_));
 NAND3_X1 _07651_ (.A1(_01566_),
    .A2(\registers[5][31] ),
    .A3(_01569_),
    .ZN(_01577_));
 OAI21_X1 _07652_ (.A(_01577_),
    .B1(_01573_),
    .B2(_01478_),
    .ZN(_00193_));
 NAND3_X1 _07653_ (.A1(_01566_),
    .A2(\registers[5][3] ),
    .A3(_01569_),
    .ZN(_01578_));
 OAI21_X1 _07654_ (.A(_01578_),
    .B1(_01573_),
    .B2(_01480_),
    .ZN(_00194_));
 BUF_X4 _07655_ (.A(_01536_),
    .Z(_01579_));
 NAND3_X1 _07656_ (.A1(_01579_),
    .A2(\registers[5][4] ),
    .A3(_01569_),
    .ZN(_01580_));
 OAI21_X1 _07657_ (.A(_01580_),
    .B1(_01573_),
    .B2(_01482_),
    .ZN(_00195_));
 NAND3_X1 _07658_ (.A1(_01579_),
    .A2(\registers[5][5] ),
    .A3(_01569_),
    .ZN(_01581_));
 OAI21_X1 _07659_ (.A(_01581_),
    .B1(_01573_),
    .B2(_01484_),
    .ZN(_00196_));
 NAND3_X1 _07660_ (.A1(_01579_),
    .A2(\registers[5][6] ),
    .A3(_01544_),
    .ZN(_01582_));
 OAI21_X1 _07661_ (.A(_01582_),
    .B1(_01573_),
    .B2(_01486_),
    .ZN(_00197_));
 NAND3_X1 _07662_ (.A1(_01579_),
    .A2(\registers[5][7] ),
    .A3(_01544_),
    .ZN(_01583_));
 OAI21_X1 _07663_ (.A(_01583_),
    .B1(_01573_),
    .B2(_01488_),
    .ZN(_00198_));
 NAND3_X1 _07664_ (.A1(_01579_),
    .A2(\registers[5][8] ),
    .A3(_01544_),
    .ZN(_01584_));
 OAI21_X1 _07665_ (.A(_01584_),
    .B1(_01545_),
    .B2(_01491_),
    .ZN(_00199_));
 NAND3_X1 _07666_ (.A1(_01579_),
    .A2(\registers[5][9] ),
    .A3(_01544_),
    .ZN(_01585_));
 OAI21_X1 _07667_ (.A(_01585_),
    .B1(_01545_),
    .B2(_01493_),
    .ZN(_00200_));
 NOR4_X2 _07668_ (.A1(_01090_),
    .A2(_01091_),
    .A3(_01494_),
    .A4(_01141_),
    .ZN(_01586_));
 BUF_X4 _07669_ (.A(_01586_),
    .Z(_01587_));
 BUF_X4 _07670_ (.A(_01587_),
    .Z(_01588_));
 NAND2_X1 _07671_ (.A1(_01137_),
    .A2(_01588_),
    .ZN(_01589_));
 NAND2_X1 _07672_ (.A1(_01408_),
    .A2(\registers[6][0] ),
    .ZN(_01590_));
 CLKBUF_X3 _07673_ (.A(_01587_),
    .Z(_01591_));
 OAI21_X1 _07674_ (.A(_01589_),
    .B1(_01590_),
    .B2(_01591_),
    .ZN(_00201_));
 NAND2_X1 _07675_ (.A1(_01149_),
    .A2(_01588_),
    .ZN(_01592_));
 NAND2_X1 _07676_ (.A1(_01408_),
    .A2(\registers[6][10] ),
    .ZN(_01593_));
 OAI21_X1 _07677_ (.A(_01592_),
    .B1(_01593_),
    .B2(_01591_),
    .ZN(_00202_));
 NAND2_X1 _07678_ (.A1(_01153_),
    .A2(_01588_),
    .ZN(_01594_));
 NAND2_X1 _07679_ (.A1(_01408_),
    .A2(\registers[6][11] ),
    .ZN(_01595_));
 OAI21_X1 _07680_ (.A(_01594_),
    .B1(_01595_),
    .B2(_01591_),
    .ZN(_00203_));
 NAND2_X1 _07681_ (.A1(_01158_),
    .A2(_01588_),
    .ZN(_01596_));
 NAND2_X1 _07682_ (.A1(_01408_),
    .A2(\registers[6][12] ),
    .ZN(_01597_));
 OAI21_X1 _07683_ (.A(_01596_),
    .B1(_01597_),
    .B2(_01591_),
    .ZN(_00204_));
 NAND2_X1 _07684_ (.A1(_01162_),
    .A2(_01588_),
    .ZN(_01598_));
 NAND2_X1 _07685_ (.A1(_01408_),
    .A2(\registers[6][13] ),
    .ZN(_01599_));
 OAI21_X1 _07686_ (.A(_01598_),
    .B1(_01599_),
    .B2(_01591_),
    .ZN(_00205_));
 NAND2_X1 _07687_ (.A1(_01166_),
    .A2(_01588_),
    .ZN(_01600_));
 NAND2_X1 _07688_ (.A1(_01408_),
    .A2(\registers[6][14] ),
    .ZN(_01601_));
 OAI21_X1 _07689_ (.A(_01600_),
    .B1(_01601_),
    .B2(_01591_),
    .ZN(_00206_));
 NAND2_X1 _07690_ (.A1(_01170_),
    .A2(_01588_),
    .ZN(_01602_));
 CLKBUF_X3 _07691_ (.A(_01267_),
    .Z(_01603_));
 NAND2_X1 _07692_ (.A1(_01603_),
    .A2(\registers[6][15] ),
    .ZN(_01604_));
 OAI21_X1 _07693_ (.A(_01602_),
    .B1(_01604_),
    .B2(_01591_),
    .ZN(_00207_));
 NAND2_X1 _07694_ (.A1(_01174_),
    .A2(_01588_),
    .ZN(_01605_));
 NAND2_X1 _07695_ (.A1(_01603_),
    .A2(\registers[6][16] ),
    .ZN(_01606_));
 OAI21_X1 _07696_ (.A(_01605_),
    .B1(_01606_),
    .B2(_01591_),
    .ZN(_00208_));
 BUF_X4 _07697_ (.A(_01587_),
    .Z(_01607_));
 NAND2_X1 _07698_ (.A1(_01178_),
    .A2(_01607_),
    .ZN(_01608_));
 NAND2_X1 _07699_ (.A1(_01603_),
    .A2(\registers[6][17] ),
    .ZN(_01609_));
 OAI21_X1 _07700_ (.A(_01608_),
    .B1(_01609_),
    .B2(_01591_),
    .ZN(_00209_));
 NAND2_X1 _07701_ (.A1(_01183_),
    .A2(_01607_),
    .ZN(_01610_));
 NAND2_X1 _07702_ (.A1(_01603_),
    .A2(\registers[6][18] ),
    .ZN(_01611_));
 OAI21_X1 _07703_ (.A(_01610_),
    .B1(_01611_),
    .B2(_01591_),
    .ZN(_00210_));
 NAND2_X1 _07704_ (.A1(_01187_),
    .A2(_01607_),
    .ZN(_01612_));
 NAND2_X1 _07705_ (.A1(_01603_),
    .A2(\registers[6][19] ),
    .ZN(_01613_));
 CLKBUF_X3 _07706_ (.A(_01587_),
    .Z(_01614_));
 OAI21_X1 _07707_ (.A(_01612_),
    .B1(_01613_),
    .B2(_01614_),
    .ZN(_00211_));
 NAND2_X1 _07708_ (.A1(_01192_),
    .A2(_01607_),
    .ZN(_01615_));
 NAND2_X1 _07709_ (.A1(_01603_),
    .A2(\registers[6][1] ),
    .ZN(_01616_));
 OAI21_X1 _07710_ (.A(_01615_),
    .B1(_01616_),
    .B2(_01614_),
    .ZN(_00212_));
 NAND2_X1 _07711_ (.A1(_01196_),
    .A2(_01607_),
    .ZN(_01617_));
 NAND2_X1 _07712_ (.A1(_01603_),
    .A2(\registers[6][20] ),
    .ZN(_01618_));
 OAI21_X1 _07713_ (.A(_01617_),
    .B1(_01618_),
    .B2(_01614_),
    .ZN(_00213_));
 NAND2_X1 _07714_ (.A1(_01201_),
    .A2(_01607_),
    .ZN(_01619_));
 NAND2_X1 _07715_ (.A1(_01603_),
    .A2(\registers[6][21] ),
    .ZN(_01620_));
 OAI21_X1 _07716_ (.A(_01619_),
    .B1(_01620_),
    .B2(_01614_),
    .ZN(_00214_));
 NAND2_X1 _07717_ (.A1(_01205_),
    .A2(_01607_),
    .ZN(_01621_));
 NAND2_X1 _07718_ (.A1(_01603_),
    .A2(\registers[6][22] ),
    .ZN(_01622_));
 OAI21_X1 _07719_ (.A(_01621_),
    .B1(_01622_),
    .B2(_01614_),
    .ZN(_00215_));
 NAND2_X1 _07720_ (.A1(_01209_),
    .A2(_01607_),
    .ZN(_01623_));
 NAND2_X1 _07721_ (.A1(_01603_),
    .A2(\registers[6][23] ),
    .ZN(_01624_));
 OAI21_X1 _07722_ (.A(_01623_),
    .B1(_01624_),
    .B2(_01614_),
    .ZN(_00216_));
 NAND2_X1 _07723_ (.A1(_01213_),
    .A2(_01607_),
    .ZN(_01625_));
 CLKBUF_X3 _07724_ (.A(_01267_),
    .Z(_01626_));
 NAND2_X1 _07725_ (.A1(_01626_),
    .A2(\registers[6][24] ),
    .ZN(_01627_));
 OAI21_X1 _07726_ (.A(_01625_),
    .B1(_01627_),
    .B2(_01614_),
    .ZN(_00217_));
 NAND2_X1 _07727_ (.A1(_01217_),
    .A2(_01607_),
    .ZN(_01628_));
 NAND2_X1 _07728_ (.A1(_01626_),
    .A2(\registers[6][25] ),
    .ZN(_01629_));
 OAI21_X1 _07729_ (.A(_01628_),
    .B1(_01629_),
    .B2(_01614_),
    .ZN(_00218_));
 BUF_X4 _07730_ (.A(_01587_),
    .Z(_01630_));
 NAND2_X1 _07731_ (.A1(_01221_),
    .A2(_01630_),
    .ZN(_01631_));
 NAND2_X1 _07732_ (.A1(_01626_),
    .A2(\registers[6][26] ),
    .ZN(_01632_));
 OAI21_X1 _07733_ (.A(_01631_),
    .B1(_01632_),
    .B2(_01614_),
    .ZN(_00219_));
 NAND2_X1 _07734_ (.A1(_01226_),
    .A2(_01630_),
    .ZN(_01633_));
 NAND2_X1 _07735_ (.A1(_01626_),
    .A2(\registers[6][27] ),
    .ZN(_01634_));
 OAI21_X1 _07736_ (.A(_01633_),
    .B1(_01634_),
    .B2(_01614_),
    .ZN(_00220_));
 NAND2_X1 _07737_ (.A1(_01230_),
    .A2(_01630_),
    .ZN(_01635_));
 NAND2_X1 _07738_ (.A1(_01626_),
    .A2(\registers[6][28] ),
    .ZN(_01636_));
 CLKBUF_X3 _07739_ (.A(_01587_),
    .Z(_01637_));
 OAI21_X1 _07740_ (.A(_01635_),
    .B1(_01636_),
    .B2(_01637_),
    .ZN(_00221_));
 NAND2_X1 _07741_ (.A1(_01235_),
    .A2(_01630_),
    .ZN(_01638_));
 NAND2_X1 _07742_ (.A1(_01626_),
    .A2(\registers[6][29] ),
    .ZN(_01639_));
 OAI21_X1 _07743_ (.A(_01638_),
    .B1(_01639_),
    .B2(_01637_),
    .ZN(_00222_));
 NAND2_X1 _07744_ (.A1(_01239_),
    .A2(_01630_),
    .ZN(_01640_));
 NAND2_X1 _07745_ (.A1(_01626_),
    .A2(\registers[6][2] ),
    .ZN(_01641_));
 OAI21_X1 _07746_ (.A(_01640_),
    .B1(_01641_),
    .B2(_01637_),
    .ZN(_00223_));
 NAND2_X1 _07747_ (.A1(_01244_),
    .A2(_01630_),
    .ZN(_01642_));
 NAND2_X1 _07748_ (.A1(_01626_),
    .A2(\registers[6][30] ),
    .ZN(_01643_));
 OAI21_X1 _07749_ (.A(_01642_),
    .B1(_01643_),
    .B2(_01637_),
    .ZN(_00224_));
 NAND2_X1 _07750_ (.A1(_01089_),
    .A2(_01630_),
    .ZN(_01644_));
 NAND2_X1 _07751_ (.A1(_01626_),
    .A2(\registers[6][31] ),
    .ZN(_01645_));
 OAI21_X1 _07752_ (.A(_01644_),
    .B1(_01645_),
    .B2(_01637_),
    .ZN(_00225_));
 NAND2_X1 _07753_ (.A1(_01109_),
    .A2(_01630_),
    .ZN(_01646_));
 NAND2_X1 _07754_ (.A1(_01626_),
    .A2(\registers[6][3] ),
    .ZN(_01647_));
 OAI21_X1 _07755_ (.A(_01646_),
    .B1(_01647_),
    .B2(_01637_),
    .ZN(_00226_));
 NAND2_X1 _07756_ (.A1(_01113_),
    .A2(_01630_),
    .ZN(_01648_));
 BUF_X4 _07757_ (.A(_01267_),
    .Z(_01649_));
 NAND2_X1 _07758_ (.A1(_01649_),
    .A2(\registers[6][4] ),
    .ZN(_01650_));
 OAI21_X1 _07759_ (.A(_01648_),
    .B1(_01650_),
    .B2(_01637_),
    .ZN(_00227_));
 NAND2_X1 _07760_ (.A1(_01117_),
    .A2(_01630_),
    .ZN(_01651_));
 NAND2_X1 _07761_ (.A1(_01649_),
    .A2(\registers[6][5] ),
    .ZN(_01652_));
 OAI21_X1 _07762_ (.A(_01651_),
    .B1(_01652_),
    .B2(_01637_),
    .ZN(_00228_));
 NAND2_X1 _07763_ (.A1(_01121_),
    .A2(_01587_),
    .ZN(_01653_));
 NAND2_X1 _07764_ (.A1(_01649_),
    .A2(\registers[6][6] ),
    .ZN(_01654_));
 OAI21_X1 _07765_ (.A(_01653_),
    .B1(_01654_),
    .B2(_01637_),
    .ZN(_00229_));
 NAND2_X1 _07766_ (.A1(_01125_),
    .A2(_01587_),
    .ZN(_01655_));
 NAND2_X1 _07767_ (.A1(_01649_),
    .A2(\registers[6][7] ),
    .ZN(_01656_));
 OAI21_X1 _07768_ (.A(_01655_),
    .B1(_01656_),
    .B2(_01637_),
    .ZN(_00230_));
 NAND2_X1 _07769_ (.A1(_01129_),
    .A2(_01587_),
    .ZN(_01657_));
 NAND2_X1 _07770_ (.A1(_01649_),
    .A2(\registers[6][8] ),
    .ZN(_01658_));
 OAI21_X1 _07771_ (.A(_01657_),
    .B1(_01658_),
    .B2(_01588_),
    .ZN(_00231_));
 NAND2_X1 _07772_ (.A1(_01133_),
    .A2(_01587_),
    .ZN(_01659_));
 NAND2_X1 _07773_ (.A1(_01649_),
    .A2(\registers[6][9] ),
    .ZN(_01660_));
 OAI21_X1 _07774_ (.A(_01659_),
    .B1(_01660_),
    .B2(_01588_),
    .ZN(_00232_));
 NOR4_X2 _07775_ (.A1(_01090_),
    .A2(_01091_),
    .A3(_01494_),
    .A4(_01340_),
    .ZN(_01661_));
 BUF_X4 _07776_ (.A(_01661_),
    .Z(_01662_));
 BUF_X4 _07777_ (.A(_01662_),
    .Z(_01663_));
 NAND2_X1 _07778_ (.A1(_01137_),
    .A2(_01663_),
    .ZN(_01664_));
 NAND2_X1 _07779_ (.A1(_01649_),
    .A2(\registers[7][0] ),
    .ZN(_01665_));
 CLKBUF_X3 _07780_ (.A(_01662_),
    .Z(_01666_));
 OAI21_X1 _07781_ (.A(_01664_),
    .B1(_01665_),
    .B2(_01666_),
    .ZN(_00233_));
 NAND2_X1 _07782_ (.A1(_01149_),
    .A2(_01663_),
    .ZN(_01667_));
 NAND2_X1 _07783_ (.A1(_01649_),
    .A2(\registers[7][10] ),
    .ZN(_01668_));
 OAI21_X1 _07784_ (.A(_01667_),
    .B1(_01668_),
    .B2(_01666_),
    .ZN(_00234_));
 NAND2_X1 _07785_ (.A1(_01153_),
    .A2(_01663_),
    .ZN(_01669_));
 NAND2_X1 _07786_ (.A1(_01649_),
    .A2(\registers[7][11] ),
    .ZN(_01670_));
 OAI21_X1 _07787_ (.A(_01669_),
    .B1(_01670_),
    .B2(_01666_),
    .ZN(_00235_));
 NAND2_X1 _07788_ (.A1(_01158_),
    .A2(_01663_),
    .ZN(_01671_));
 NAND2_X1 _07789_ (.A1(_01649_),
    .A2(\registers[7][12] ),
    .ZN(_01672_));
 OAI21_X1 _07790_ (.A(_01671_),
    .B1(_01672_),
    .B2(_01666_),
    .ZN(_00236_));
 NAND2_X1 _07791_ (.A1(_01162_),
    .A2(_01663_),
    .ZN(_01673_));
 BUF_X4 _07792_ (.A(_01103_),
    .Z(_01674_));
 CLKBUF_X3 _07793_ (.A(_01674_),
    .Z(_01675_));
 NAND2_X1 _07794_ (.A1(_01675_),
    .A2(\registers[7][13] ),
    .ZN(_01676_));
 OAI21_X1 _07795_ (.A(_01673_),
    .B1(_01676_),
    .B2(_01666_),
    .ZN(_00237_));
 NAND2_X1 _07796_ (.A1(_01166_),
    .A2(_01663_),
    .ZN(_01677_));
 NAND2_X1 _07797_ (.A1(_01675_),
    .A2(\registers[7][14] ),
    .ZN(_01678_));
 OAI21_X1 _07798_ (.A(_01677_),
    .B1(_01678_),
    .B2(_01666_),
    .ZN(_00238_));
 NAND2_X1 _07799_ (.A1(_01170_),
    .A2(_01663_),
    .ZN(_01679_));
 NAND2_X1 _07800_ (.A1(_01675_),
    .A2(\registers[7][15] ),
    .ZN(_01680_));
 OAI21_X1 _07801_ (.A(_01679_),
    .B1(_01680_),
    .B2(_01666_),
    .ZN(_00239_));
 NAND2_X1 _07802_ (.A1(_01174_),
    .A2(_01663_),
    .ZN(_01681_));
 NAND2_X1 _07803_ (.A1(_01675_),
    .A2(\registers[7][16] ),
    .ZN(_01682_));
 OAI21_X1 _07804_ (.A(_01681_),
    .B1(_01682_),
    .B2(_01666_),
    .ZN(_00240_));
 BUF_X4 _07805_ (.A(_01662_),
    .Z(_01683_));
 NAND2_X1 _07806_ (.A1(_01178_),
    .A2(_01683_),
    .ZN(_01684_));
 NAND2_X1 _07807_ (.A1(_01675_),
    .A2(\registers[7][17] ),
    .ZN(_01685_));
 OAI21_X1 _07808_ (.A(_01684_),
    .B1(_01685_),
    .B2(_01666_),
    .ZN(_00241_));
 NAND2_X1 _07809_ (.A1(_01183_),
    .A2(_01683_),
    .ZN(_01686_));
 NAND2_X1 _07810_ (.A1(_01675_),
    .A2(\registers[7][18] ),
    .ZN(_01687_));
 OAI21_X1 _07811_ (.A(_01686_),
    .B1(_01687_),
    .B2(_01666_),
    .ZN(_00242_));
 NAND2_X1 _07812_ (.A1(_01187_),
    .A2(_01683_),
    .ZN(_01688_));
 NAND2_X1 _07813_ (.A1(_01675_),
    .A2(\registers[7][19] ),
    .ZN(_01689_));
 CLKBUF_X3 _07814_ (.A(_01662_),
    .Z(_01690_));
 OAI21_X1 _07815_ (.A(_01688_),
    .B1(_01689_),
    .B2(_01690_),
    .ZN(_00243_));
 NAND2_X1 _07816_ (.A1(_01192_),
    .A2(_01683_),
    .ZN(_01691_));
 NAND2_X1 _07817_ (.A1(_01675_),
    .A2(\registers[7][1] ),
    .ZN(_01692_));
 OAI21_X1 _07818_ (.A(_01691_),
    .B1(_01692_),
    .B2(_01690_),
    .ZN(_00244_));
 NAND2_X1 _07819_ (.A1(_01196_),
    .A2(_01683_),
    .ZN(_01693_));
 NAND2_X1 _07820_ (.A1(_01675_),
    .A2(\registers[7][20] ),
    .ZN(_01694_));
 OAI21_X1 _07821_ (.A(_01693_),
    .B1(_01694_),
    .B2(_01690_),
    .ZN(_00245_));
 NAND2_X1 _07822_ (.A1(_01201_),
    .A2(_01683_),
    .ZN(_01695_));
 NAND2_X1 _07823_ (.A1(_01675_),
    .A2(\registers[7][21] ),
    .ZN(_01696_));
 OAI21_X1 _07824_ (.A(_01695_),
    .B1(_01696_),
    .B2(_01690_),
    .ZN(_00246_));
 NAND2_X1 _07825_ (.A1(_01205_),
    .A2(_01683_),
    .ZN(_01697_));
 CLKBUF_X3 _07826_ (.A(_01674_),
    .Z(_01698_));
 NAND2_X1 _07827_ (.A1(_01698_),
    .A2(\registers[7][22] ),
    .ZN(_01699_));
 OAI21_X1 _07828_ (.A(_01697_),
    .B1(_01699_),
    .B2(_01690_),
    .ZN(_00247_));
 NAND2_X1 _07829_ (.A1(_01209_),
    .A2(_01683_),
    .ZN(_01700_));
 NAND2_X1 _07830_ (.A1(_01698_),
    .A2(\registers[7][23] ),
    .ZN(_01701_));
 OAI21_X1 _07831_ (.A(_01700_),
    .B1(_01701_),
    .B2(_01690_),
    .ZN(_00248_));
 NAND2_X1 _07832_ (.A1(_01213_),
    .A2(_01683_),
    .ZN(_01702_));
 NAND2_X1 _07833_ (.A1(_01698_),
    .A2(\registers[7][24] ),
    .ZN(_01703_));
 OAI21_X1 _07834_ (.A(_01702_),
    .B1(_01703_),
    .B2(_01690_),
    .ZN(_00249_));
 NAND2_X1 _07835_ (.A1(_01217_),
    .A2(_01683_),
    .ZN(_01704_));
 NAND2_X1 _07836_ (.A1(_01698_),
    .A2(\registers[7][25] ),
    .ZN(_01705_));
 OAI21_X1 _07837_ (.A(_01704_),
    .B1(_01705_),
    .B2(_01690_),
    .ZN(_00250_));
 BUF_X4 _07838_ (.A(_01662_),
    .Z(_01706_));
 NAND2_X1 _07839_ (.A1(_01221_),
    .A2(_01706_),
    .ZN(_01707_));
 NAND2_X1 _07840_ (.A1(_01698_),
    .A2(\registers[7][26] ),
    .ZN(_01708_));
 OAI21_X1 _07841_ (.A(_01707_),
    .B1(_01708_),
    .B2(_01690_),
    .ZN(_00251_));
 NAND2_X1 _07842_ (.A1(_01226_),
    .A2(_01706_),
    .ZN(_01709_));
 NAND2_X1 _07843_ (.A1(_01698_),
    .A2(\registers[7][27] ),
    .ZN(_01710_));
 OAI21_X1 _07844_ (.A(_01709_),
    .B1(_01710_),
    .B2(_01690_),
    .ZN(_00252_));
 NAND2_X1 _07845_ (.A1(_01230_),
    .A2(_01706_),
    .ZN(_01711_));
 NAND2_X1 _07846_ (.A1(_01698_),
    .A2(\registers[7][28] ),
    .ZN(_01712_));
 CLKBUF_X3 _07847_ (.A(_01662_),
    .Z(_01713_));
 OAI21_X1 _07848_ (.A(_01711_),
    .B1(_01712_),
    .B2(_01713_),
    .ZN(_00253_));
 NAND2_X1 _07849_ (.A1(_01235_),
    .A2(_01706_),
    .ZN(_01714_));
 NAND2_X1 _07850_ (.A1(_01698_),
    .A2(\registers[7][29] ),
    .ZN(_01715_));
 OAI21_X1 _07851_ (.A(_01714_),
    .B1(_01715_),
    .B2(_01713_),
    .ZN(_00254_));
 NAND2_X1 _07852_ (.A1(_01239_),
    .A2(_01706_),
    .ZN(_01716_));
 NAND2_X1 _07853_ (.A1(_01698_),
    .A2(\registers[7][2] ),
    .ZN(_01717_));
 OAI21_X1 _07854_ (.A(_01716_),
    .B1(_01717_),
    .B2(_01713_),
    .ZN(_00255_));
 NAND2_X1 _07855_ (.A1(_01244_),
    .A2(_01706_),
    .ZN(_01718_));
 NAND2_X1 _07856_ (.A1(_01698_),
    .A2(\registers[7][30] ),
    .ZN(_01719_));
 OAI21_X1 _07857_ (.A(_01718_),
    .B1(_01719_),
    .B2(_01713_),
    .ZN(_00256_));
 NAND2_X1 _07858_ (.A1(_01089_),
    .A2(_01706_),
    .ZN(_01720_));
 BUF_X4 _07859_ (.A(_01674_),
    .Z(_01721_));
 NAND2_X1 _07860_ (.A1(_01721_),
    .A2(\registers[7][31] ),
    .ZN(_01722_));
 OAI21_X1 _07861_ (.A(_01720_),
    .B1(_01722_),
    .B2(_01713_),
    .ZN(_00257_));
 NAND2_X1 _07862_ (.A1(_01109_),
    .A2(_01706_),
    .ZN(_01723_));
 NAND2_X1 _07863_ (.A1(_01721_),
    .A2(\registers[7][3] ),
    .ZN(_01724_));
 OAI21_X1 _07864_ (.A(_01723_),
    .B1(_01724_),
    .B2(_01713_),
    .ZN(_00258_));
 NAND2_X1 _07865_ (.A1(_01113_),
    .A2(_01706_),
    .ZN(_01725_));
 NAND2_X1 _07866_ (.A1(_01721_),
    .A2(\registers[7][4] ),
    .ZN(_01726_));
 OAI21_X1 _07867_ (.A(_01725_),
    .B1(_01726_),
    .B2(_01713_),
    .ZN(_00259_));
 NAND2_X1 _07868_ (.A1(_01117_),
    .A2(_01706_),
    .ZN(_01727_));
 NAND2_X1 _07869_ (.A1(_01721_),
    .A2(\registers[7][5] ),
    .ZN(_01728_));
 OAI21_X1 _07870_ (.A(_01727_),
    .B1(_01728_),
    .B2(_01713_),
    .ZN(_00260_));
 NAND2_X1 _07871_ (.A1(_01121_),
    .A2(_01662_),
    .ZN(_01729_));
 NAND2_X1 _07872_ (.A1(_01721_),
    .A2(\registers[7][6] ),
    .ZN(_01730_));
 OAI21_X1 _07873_ (.A(_01729_),
    .B1(_01730_),
    .B2(_01713_),
    .ZN(_00261_));
 NAND2_X1 _07874_ (.A1(_01125_),
    .A2(_01662_),
    .ZN(_01731_));
 NAND2_X1 _07875_ (.A1(_01721_),
    .A2(\registers[7][7] ),
    .ZN(_01732_));
 OAI21_X1 _07876_ (.A(_01731_),
    .B1(_01732_),
    .B2(_01713_),
    .ZN(_00262_));
 NAND2_X1 _07877_ (.A1(_01129_),
    .A2(_01662_),
    .ZN(_01733_));
 NAND2_X1 _07878_ (.A1(_01721_),
    .A2(\registers[7][8] ),
    .ZN(_01734_));
 OAI21_X1 _07879_ (.A(_01733_),
    .B1(_01734_),
    .B2(_01663_),
    .ZN(_00263_));
 NAND2_X1 _07880_ (.A1(_01133_),
    .A2(_01662_),
    .ZN(_01735_));
 NAND2_X1 _07881_ (.A1(_01721_),
    .A2(\registers[7][9] ),
    .ZN(_01736_));
 OAI21_X1 _07882_ (.A(_01735_),
    .B1(_01736_),
    .B2(_01663_),
    .ZN(_00264_));
 OR3_X2 _07883_ (.A1(_01096_),
    .A2(_01094_),
    .A3(_01496_),
    .ZN(_01737_));
 INV_X4 _07884_ (.A(_01091_),
    .ZN(_01738_));
 NAND3_X2 _07885_ (.A1(_01090_),
    .A2(_01738_),
    .A3(_01494_),
    .ZN(_01739_));
 OR2_X1 _07886_ (.A1(_01737_),
    .A2(_01739_),
    .ZN(_01740_));
 CLKBUF_X3 _07887_ (.A(_01740_),
    .Z(_01741_));
 CLKBUF_X3 _07888_ (.A(_01741_),
    .Z(_01742_));
 NAND3_X1 _07889_ (.A1(_01579_),
    .A2(\registers[8][0] ),
    .A3(_01742_),
    .ZN(_01743_));
 CLKBUF_X3 _07890_ (.A(_01741_),
    .Z(_01744_));
 OAI21_X1 _07891_ (.A(_01743_),
    .B1(_01744_),
    .B2(_01424_),
    .ZN(_00265_));
 NAND3_X1 _07892_ (.A1(_01579_),
    .A2(\registers[8][10] ),
    .A3(_01742_),
    .ZN(_01745_));
 OAI21_X1 _07893_ (.A(_01745_),
    .B1(_01744_),
    .B2(_01426_),
    .ZN(_00266_));
 NAND3_X1 _07894_ (.A1(_01579_),
    .A2(\registers[8][11] ),
    .A3(_01742_),
    .ZN(_01746_));
 OAI21_X1 _07895_ (.A(_01746_),
    .B1(_01744_),
    .B2(_01428_),
    .ZN(_00267_));
 NAND3_X1 _07896_ (.A1(_01579_),
    .A2(\registers[8][12] ),
    .A3(_01742_),
    .ZN(_01747_));
 OAI21_X1 _07897_ (.A(_01747_),
    .B1(_01744_),
    .B2(_01430_),
    .ZN(_00268_));
 CLKBUF_X3 _07898_ (.A(_01536_),
    .Z(_01748_));
 NAND3_X1 _07899_ (.A1(_01748_),
    .A2(\registers[8][13] ),
    .A3(_01742_),
    .ZN(_01749_));
 OAI21_X1 _07900_ (.A(_01749_),
    .B1(_01744_),
    .B2(_01432_),
    .ZN(_00269_));
 NAND3_X1 _07901_ (.A1(_01748_),
    .A2(\registers[8][14] ),
    .A3(_01742_),
    .ZN(_01750_));
 OAI21_X1 _07902_ (.A(_01750_),
    .B1(_01744_),
    .B2(_01434_),
    .ZN(_00270_));
 NAND3_X1 _07903_ (.A1(_01748_),
    .A2(\registers[8][15] ),
    .A3(_01742_),
    .ZN(_01751_));
 OAI21_X1 _07904_ (.A(_01751_),
    .B1(_01744_),
    .B2(_01436_),
    .ZN(_00271_));
 NAND3_X1 _07905_ (.A1(_01748_),
    .A2(\registers[8][16] ),
    .A3(_01742_),
    .ZN(_01752_));
 OAI21_X1 _07906_ (.A(_01752_),
    .B1(_01744_),
    .B2(_01438_),
    .ZN(_00272_));
 CLKBUF_X3 _07907_ (.A(_01741_),
    .Z(_01753_));
 NAND3_X1 _07908_ (.A1(_01748_),
    .A2(\registers[8][17] ),
    .A3(_01753_),
    .ZN(_01754_));
 OAI21_X1 _07909_ (.A(_01754_),
    .B1(_01744_),
    .B2(_01441_),
    .ZN(_00273_));
 NAND3_X1 _07910_ (.A1(_01748_),
    .A2(\registers[8][18] ),
    .A3(_01753_),
    .ZN(_01755_));
 OAI21_X1 _07911_ (.A(_01755_),
    .B1(_01744_),
    .B2(_01443_),
    .ZN(_00274_));
 NAND3_X1 _07912_ (.A1(_01748_),
    .A2(\registers[8][19] ),
    .A3(_01753_),
    .ZN(_01756_));
 CLKBUF_X3 _07913_ (.A(_01741_),
    .Z(_01757_));
 OAI21_X1 _07914_ (.A(_01756_),
    .B1(_01757_),
    .B2(_01447_),
    .ZN(_00275_));
 NAND3_X1 _07915_ (.A1(_01748_),
    .A2(\registers[8][1] ),
    .A3(_01753_),
    .ZN(_01758_));
 OAI21_X1 _07916_ (.A(_01758_),
    .B1(_01757_),
    .B2(_01449_),
    .ZN(_00276_));
 NAND3_X1 _07917_ (.A1(_01748_),
    .A2(\registers[8][20] ),
    .A3(_01753_),
    .ZN(_01759_));
 OAI21_X1 _07918_ (.A(_01759_),
    .B1(_01757_),
    .B2(_01451_),
    .ZN(_00277_));
 NAND3_X1 _07919_ (.A1(_01748_),
    .A2(\registers[8][21] ),
    .A3(_01753_),
    .ZN(_01760_));
 OAI21_X1 _07920_ (.A(_01760_),
    .B1(_01757_),
    .B2(_01453_),
    .ZN(_00278_));
 CLKBUF_X3 _07921_ (.A(_01536_),
    .Z(_01761_));
 NAND3_X1 _07922_ (.A1(_01761_),
    .A2(\registers[8][22] ),
    .A3(_01753_),
    .ZN(_01762_));
 OAI21_X1 _07923_ (.A(_01762_),
    .B1(_01757_),
    .B2(_01455_),
    .ZN(_00279_));
 NAND3_X1 _07924_ (.A1(_01761_),
    .A2(\registers[8][23] ),
    .A3(_01753_),
    .ZN(_01763_));
 OAI21_X1 _07925_ (.A(_01763_),
    .B1(_01757_),
    .B2(_01457_),
    .ZN(_00280_));
 NAND3_X1 _07926_ (.A1(_01761_),
    .A2(\registers[8][24] ),
    .A3(_01753_),
    .ZN(_01764_));
 OAI21_X1 _07927_ (.A(_01764_),
    .B1(_01757_),
    .B2(_01459_),
    .ZN(_00281_));
 NAND3_X1 _07928_ (.A1(_01761_),
    .A2(\registers[8][25] ),
    .A3(_01753_),
    .ZN(_01765_));
 OAI21_X1 _07929_ (.A(_01765_),
    .B1(_01757_),
    .B2(_01461_),
    .ZN(_00282_));
 CLKBUF_X3 _07930_ (.A(_01741_),
    .Z(_01766_));
 NAND3_X1 _07931_ (.A1(_01761_),
    .A2(\registers[8][26] ),
    .A3(_01766_),
    .ZN(_01767_));
 OAI21_X1 _07932_ (.A(_01767_),
    .B1(_01757_),
    .B2(_01464_),
    .ZN(_00283_));
 NAND3_X1 _07933_ (.A1(_01761_),
    .A2(\registers[8][27] ),
    .A3(_01766_),
    .ZN(_01768_));
 OAI21_X1 _07934_ (.A(_01768_),
    .B1(_01757_),
    .B2(_01466_),
    .ZN(_00284_));
 NAND3_X1 _07935_ (.A1(_01761_),
    .A2(\registers[8][28] ),
    .A3(_01766_),
    .ZN(_01769_));
 CLKBUF_X3 _07936_ (.A(_01741_),
    .Z(_01770_));
 OAI21_X1 _07937_ (.A(_01769_),
    .B1(_01770_),
    .B2(_01470_),
    .ZN(_00285_));
 NAND3_X1 _07938_ (.A1(_01761_),
    .A2(\registers[8][29] ),
    .A3(_01766_),
    .ZN(_01771_));
 OAI21_X1 _07939_ (.A(_01771_),
    .B1(_01770_),
    .B2(_01472_),
    .ZN(_00286_));
 NAND3_X1 _07940_ (.A1(_01761_),
    .A2(\registers[8][2] ),
    .A3(_01766_),
    .ZN(_01772_));
 OAI21_X1 _07941_ (.A(_01772_),
    .B1(_01770_),
    .B2(_01474_),
    .ZN(_00287_));
 NAND3_X1 _07942_ (.A1(_01761_),
    .A2(\registers[8][30] ),
    .A3(_01766_),
    .ZN(_01773_));
 OAI21_X1 _07943_ (.A(_01773_),
    .B1(_01770_),
    .B2(_01476_),
    .ZN(_00288_));
 BUF_X4 _07944_ (.A(_01536_),
    .Z(_01774_));
 NAND3_X1 _07945_ (.A1(_01774_),
    .A2(\registers[8][31] ),
    .A3(_01766_),
    .ZN(_01775_));
 OAI21_X1 _07946_ (.A(_01775_),
    .B1(_01770_),
    .B2(_01478_),
    .ZN(_00289_));
 NAND3_X1 _07947_ (.A1(_01774_),
    .A2(\registers[8][3] ),
    .A3(_01766_),
    .ZN(_01776_));
 OAI21_X1 _07948_ (.A(_01776_),
    .B1(_01770_),
    .B2(_01480_),
    .ZN(_00290_));
 NAND3_X1 _07949_ (.A1(_01774_),
    .A2(\registers[8][4] ),
    .A3(_01766_),
    .ZN(_01777_));
 OAI21_X1 _07950_ (.A(_01777_),
    .B1(_01770_),
    .B2(_01482_),
    .ZN(_00291_));
 NAND3_X1 _07951_ (.A1(_01774_),
    .A2(\registers[8][5] ),
    .A3(_01766_),
    .ZN(_01778_));
 OAI21_X1 _07952_ (.A(_01778_),
    .B1(_01770_),
    .B2(_01484_),
    .ZN(_00292_));
 NAND3_X1 _07953_ (.A1(_01774_),
    .A2(\registers[8][6] ),
    .A3(_01741_),
    .ZN(_01779_));
 OAI21_X1 _07954_ (.A(_01779_),
    .B1(_01770_),
    .B2(_01486_),
    .ZN(_00293_));
 NAND3_X1 _07955_ (.A1(_01774_),
    .A2(\registers[8][7] ),
    .A3(_01741_),
    .ZN(_01780_));
 OAI21_X1 _07956_ (.A(_01780_),
    .B1(_01770_),
    .B2(_01488_),
    .ZN(_00294_));
 NAND3_X1 _07957_ (.A1(_01774_),
    .A2(\registers[8][8] ),
    .A3(_01741_),
    .ZN(_01781_));
 OAI21_X1 _07958_ (.A(_01781_),
    .B1(_01742_),
    .B2(_01491_),
    .ZN(_00295_));
 NAND3_X1 _07959_ (.A1(_01774_),
    .A2(\registers[8][9] ),
    .A3(_01741_),
    .ZN(_01782_));
 OAI21_X1 _07960_ (.A(_01782_),
    .B1(_01742_),
    .B2(_01493_),
    .ZN(_00296_));
 NOR2_X1 _07961_ (.A1(_01098_),
    .A2(_01739_),
    .ZN(_01783_));
 BUF_X4 _07962_ (.A(_01783_),
    .Z(_01784_));
 CLKBUF_X3 _07963_ (.A(_01784_),
    .Z(_01785_));
 NAND2_X1 _07964_ (.A1(_01137_),
    .A2(_01785_),
    .ZN(_01786_));
 NAND2_X1 _07965_ (.A1(_01721_),
    .A2(\registers[9][0] ),
    .ZN(_01787_));
 CLKBUF_X3 _07966_ (.A(_01784_),
    .Z(_01788_));
 OAI21_X1 _07967_ (.A(_01786_),
    .B1(_01787_),
    .B2(_01788_),
    .ZN(_00297_));
 NAND2_X1 _07968_ (.A1(_01149_),
    .A2(_01785_),
    .ZN(_01789_));
 NAND2_X1 _07969_ (.A1(_01721_),
    .A2(\registers[9][10] ),
    .ZN(_01790_));
 OAI21_X1 _07970_ (.A(_01789_),
    .B1(_01790_),
    .B2(_01788_),
    .ZN(_00298_));
 NAND2_X1 _07971_ (.A1(_01153_),
    .A2(_01785_),
    .ZN(_01791_));
 CLKBUF_X3 _07972_ (.A(_01674_),
    .Z(_01792_));
 NAND2_X1 _07973_ (.A1(_01792_),
    .A2(\registers[9][11] ),
    .ZN(_01793_));
 OAI21_X1 _07974_ (.A(_01791_),
    .B1(_01793_),
    .B2(_01788_),
    .ZN(_00299_));
 NAND2_X1 _07975_ (.A1(_01158_),
    .A2(_01785_),
    .ZN(_01794_));
 NAND2_X1 _07976_ (.A1(_01792_),
    .A2(\registers[9][12] ),
    .ZN(_01795_));
 OAI21_X1 _07977_ (.A(_01794_),
    .B1(_01795_),
    .B2(_01788_),
    .ZN(_00300_));
 NAND2_X1 _07978_ (.A1(_01162_),
    .A2(_01785_),
    .ZN(_01796_));
 NAND2_X1 _07979_ (.A1(_01792_),
    .A2(\registers[9][13] ),
    .ZN(_01797_));
 OAI21_X1 _07980_ (.A(_01796_),
    .B1(_01797_),
    .B2(_01788_),
    .ZN(_00301_));
 NAND2_X1 _07981_ (.A1(_01166_),
    .A2(_01785_),
    .ZN(_01798_));
 NAND2_X1 _07982_ (.A1(_01792_),
    .A2(\registers[9][14] ),
    .ZN(_01799_));
 OAI21_X1 _07983_ (.A(_01798_),
    .B1(_01799_),
    .B2(_01788_),
    .ZN(_00302_));
 NAND2_X1 _07984_ (.A1(_01170_),
    .A2(_01785_),
    .ZN(_01800_));
 NAND2_X1 _07985_ (.A1(_01792_),
    .A2(\registers[9][15] ),
    .ZN(_01801_));
 OAI21_X1 _07986_ (.A(_01800_),
    .B1(_01801_),
    .B2(_01788_),
    .ZN(_00303_));
 NAND2_X1 _07987_ (.A1(_01174_),
    .A2(_01785_),
    .ZN(_01802_));
 NAND2_X1 _07988_ (.A1(_01792_),
    .A2(\registers[9][16] ),
    .ZN(_01803_));
 OAI21_X1 _07989_ (.A(_01802_),
    .B1(_01803_),
    .B2(_01788_),
    .ZN(_00304_));
 CLKBUF_X3 _07990_ (.A(_01784_),
    .Z(_01804_));
 NAND2_X1 _07991_ (.A1(_01178_),
    .A2(_01804_),
    .ZN(_01805_));
 NAND2_X1 _07992_ (.A1(_01792_),
    .A2(\registers[9][17] ),
    .ZN(_01806_));
 OAI21_X1 _07993_ (.A(_01805_),
    .B1(_01806_),
    .B2(_01788_),
    .ZN(_00305_));
 NAND2_X1 _07994_ (.A1(_01183_),
    .A2(_01804_),
    .ZN(_01807_));
 NAND2_X1 _07995_ (.A1(_01792_),
    .A2(\registers[9][18] ),
    .ZN(_01808_));
 OAI21_X1 _07996_ (.A(_01807_),
    .B1(_01808_),
    .B2(_01788_),
    .ZN(_00306_));
 NAND2_X1 _07997_ (.A1(_01187_),
    .A2(_01804_),
    .ZN(_01809_));
 NAND2_X1 _07998_ (.A1(_01792_),
    .A2(\registers[9][19] ),
    .ZN(_01810_));
 CLKBUF_X3 _07999_ (.A(_01784_),
    .Z(_01811_));
 OAI21_X1 _08000_ (.A(_01809_),
    .B1(_01810_),
    .B2(_01811_),
    .ZN(_00307_));
 NAND2_X1 _08001_ (.A1(_01192_),
    .A2(_01804_),
    .ZN(_01812_));
 NAND2_X1 _08002_ (.A1(_01792_),
    .A2(\registers[9][1] ),
    .ZN(_01813_));
 OAI21_X1 _08003_ (.A(_01812_),
    .B1(_01813_),
    .B2(_01811_),
    .ZN(_00308_));
 NAND2_X1 _08004_ (.A1(_01196_),
    .A2(_01804_),
    .ZN(_01814_));
 CLKBUF_X3 _08005_ (.A(_01674_),
    .Z(_01815_));
 NAND2_X1 _08006_ (.A1(_01815_),
    .A2(\registers[9][20] ),
    .ZN(_01816_));
 OAI21_X1 _08007_ (.A(_01814_),
    .B1(_01816_),
    .B2(_01811_),
    .ZN(_00309_));
 NAND2_X1 _08008_ (.A1(_01201_),
    .A2(_01804_),
    .ZN(_01817_));
 NAND2_X1 _08009_ (.A1(_01815_),
    .A2(\registers[9][21] ),
    .ZN(_01818_));
 OAI21_X1 _08010_ (.A(_01817_),
    .B1(_01818_),
    .B2(_01811_),
    .ZN(_00310_));
 NAND2_X1 _08011_ (.A1(_01205_),
    .A2(_01804_),
    .ZN(_01819_));
 NAND2_X1 _08012_ (.A1(_01815_),
    .A2(\registers[9][22] ),
    .ZN(_01820_));
 OAI21_X1 _08013_ (.A(_01819_),
    .B1(_01820_),
    .B2(_01811_),
    .ZN(_00311_));
 NAND2_X1 _08014_ (.A1(_01209_),
    .A2(_01804_),
    .ZN(_01821_));
 NAND2_X1 _08015_ (.A1(_01815_),
    .A2(\registers[9][23] ),
    .ZN(_01822_));
 OAI21_X1 _08016_ (.A(_01821_),
    .B1(_01822_),
    .B2(_01811_),
    .ZN(_00312_));
 NAND2_X1 _08017_ (.A1(_01213_),
    .A2(_01804_),
    .ZN(_01823_));
 NAND2_X1 _08018_ (.A1(_01815_),
    .A2(\registers[9][24] ),
    .ZN(_01824_));
 OAI21_X1 _08019_ (.A(_01823_),
    .B1(_01824_),
    .B2(_01811_),
    .ZN(_00313_));
 NAND2_X1 _08020_ (.A1(_01217_),
    .A2(_01804_),
    .ZN(_01825_));
 NAND2_X1 _08021_ (.A1(_01815_),
    .A2(\registers[9][25] ),
    .ZN(_01826_));
 OAI21_X1 _08022_ (.A(_01825_),
    .B1(_01826_),
    .B2(_01811_),
    .ZN(_00314_));
 CLKBUF_X3 _08023_ (.A(_01784_),
    .Z(_01827_));
 NAND2_X1 _08024_ (.A1(_01221_),
    .A2(_01827_),
    .ZN(_01828_));
 NAND2_X1 _08025_ (.A1(_01815_),
    .A2(\registers[9][26] ),
    .ZN(_01829_));
 OAI21_X1 _08026_ (.A(_01828_),
    .B1(_01829_),
    .B2(_01811_),
    .ZN(_00315_));
 NAND2_X1 _08027_ (.A1(_01226_),
    .A2(_01827_),
    .ZN(_01830_));
 NAND2_X1 _08028_ (.A1(_01815_),
    .A2(\registers[9][27] ),
    .ZN(_01831_));
 OAI21_X1 _08029_ (.A(_01830_),
    .B1(_01831_),
    .B2(_01811_),
    .ZN(_00316_));
 NAND2_X1 _08030_ (.A1(_01230_),
    .A2(_01827_),
    .ZN(_01832_));
 NAND2_X1 _08031_ (.A1(_01815_),
    .A2(\registers[9][28] ),
    .ZN(_01833_));
 CLKBUF_X3 _08032_ (.A(_01784_),
    .Z(_01834_));
 OAI21_X1 _08033_ (.A(_01832_),
    .B1(_01833_),
    .B2(_01834_),
    .ZN(_00317_));
 NAND2_X1 _08034_ (.A1(_01235_),
    .A2(_01827_),
    .ZN(_01835_));
 NAND2_X1 _08035_ (.A1(_01815_),
    .A2(\registers[9][29] ),
    .ZN(_01836_));
 OAI21_X1 _08036_ (.A(_01835_),
    .B1(_01836_),
    .B2(_01834_),
    .ZN(_00318_));
 NAND2_X1 _08037_ (.A1(_01239_),
    .A2(_01827_),
    .ZN(_01837_));
 BUF_X4 _08038_ (.A(_01674_),
    .Z(_01838_));
 NAND2_X1 _08039_ (.A1(_01838_),
    .A2(\registers[9][2] ),
    .ZN(_01839_));
 OAI21_X1 _08040_ (.A(_01837_),
    .B1(_01839_),
    .B2(_01834_),
    .ZN(_00319_));
 NAND2_X1 _08041_ (.A1(_01244_),
    .A2(_01827_),
    .ZN(_01840_));
 NAND2_X1 _08042_ (.A1(_01838_),
    .A2(\registers[9][30] ),
    .ZN(_01841_));
 OAI21_X1 _08043_ (.A(_01840_),
    .B1(_01841_),
    .B2(_01834_),
    .ZN(_00320_));
 NAND2_X1 _08044_ (.A1(_01089_),
    .A2(_01827_),
    .ZN(_01842_));
 NAND2_X1 _08045_ (.A1(_01838_),
    .A2(\registers[9][31] ),
    .ZN(_01843_));
 OAI21_X1 _08046_ (.A(_01842_),
    .B1(_01843_),
    .B2(_01834_),
    .ZN(_00321_));
 NAND2_X1 _08047_ (.A1(_01109_),
    .A2(_01827_),
    .ZN(_01844_));
 NAND2_X1 _08048_ (.A1(_01838_),
    .A2(\registers[9][3] ),
    .ZN(_01845_));
 OAI21_X1 _08049_ (.A(_01844_),
    .B1(_01845_),
    .B2(_01834_),
    .ZN(_00322_));
 NAND2_X1 _08050_ (.A1(_01113_),
    .A2(_01827_),
    .ZN(_01846_));
 NAND2_X1 _08051_ (.A1(_01838_),
    .A2(\registers[9][4] ),
    .ZN(_01847_));
 OAI21_X1 _08052_ (.A(_01846_),
    .B1(_01847_),
    .B2(_01834_),
    .ZN(_00323_));
 NAND2_X1 _08053_ (.A1(_01117_),
    .A2(_01827_),
    .ZN(_01848_));
 NAND2_X1 _08054_ (.A1(_01838_),
    .A2(\registers[9][5] ),
    .ZN(_01849_));
 OAI21_X1 _08055_ (.A(_01848_),
    .B1(_01849_),
    .B2(_01834_),
    .ZN(_00324_));
 NAND2_X1 _08056_ (.A1(_01121_),
    .A2(_01784_),
    .ZN(_01850_));
 NAND2_X1 _08057_ (.A1(_01838_),
    .A2(\registers[9][6] ),
    .ZN(_01851_));
 OAI21_X1 _08058_ (.A(_01850_),
    .B1(_01851_),
    .B2(_01834_),
    .ZN(_00325_));
 NAND2_X1 _08059_ (.A1(_01125_),
    .A2(_01784_),
    .ZN(_01852_));
 NAND2_X1 _08060_ (.A1(_01838_),
    .A2(\registers[9][7] ),
    .ZN(_01853_));
 OAI21_X1 _08061_ (.A(_01852_),
    .B1(_01853_),
    .B2(_01834_),
    .ZN(_00326_));
 NAND2_X1 _08062_ (.A1(_01129_),
    .A2(_01784_),
    .ZN(_01854_));
 NAND2_X1 _08063_ (.A1(_01838_),
    .A2(\registers[9][8] ),
    .ZN(_01855_));
 OAI21_X1 _08064_ (.A(_01854_),
    .B1(_01855_),
    .B2(_01785_),
    .ZN(_00327_));
 NAND2_X1 _08065_ (.A1(_01133_),
    .A2(_01784_),
    .ZN(_01856_));
 NAND2_X1 _08066_ (.A1(_01838_),
    .A2(\registers[9][9] ),
    .ZN(_01857_));
 OAI21_X1 _08067_ (.A(_01856_),
    .B1(_01857_),
    .B2(_01785_),
    .ZN(_00328_));
 BUF_X2 _08068_ (.A(read_addr1[4]),
    .Z(_01858_));
 INV_X1 _08069_ (.A(_01858_),
    .ZN(_01859_));
 BUF_X4 _08070_ (.A(_01859_),
    .Z(_01860_));
 BUF_X4 _08071_ (.A(read_addr1[1]),
    .Z(_01861_));
 BUF_X16 _08072_ (.A(_01861_),
    .Z(_01862_));
 BUF_X8 _08073_ (.A(read_addr1[2]),
    .Z(_01863_));
 OR2_X1 _08074_ (.A1(_01862_),
    .A2(_01863_),
    .ZN(_01864_));
 BUF_X4 _08075_ (.A(_01864_),
    .Z(_01865_));
 BUF_X4 _08076_ (.A(_01865_),
    .Z(_01866_));
 BUF_X4 _08077_ (.A(read_addr1[0]),
    .Z(_01867_));
 BUF_X8 _08078_ (.A(_01867_),
    .Z(_01868_));
 BUF_X4 _08079_ (.A(_01868_),
    .Z(_01869_));
 MUX2_X1 _08080_ (.A(\registers[16][0] ),
    .B(\registers[17][0] ),
    .S(_01869_),
    .Z(_01870_));
 BUF_X8 _08081_ (.A(_01861_),
    .Z(_01871_));
 NAND2_X4 _08082_ (.A1(_01871_),
    .A2(_01863_),
    .ZN(_01872_));
 BUF_X4 _08083_ (.A(_01872_),
    .Z(_01873_));
 BUF_X4 _08084_ (.A(_01868_),
    .Z(_01874_));
 MUX2_X1 _08085_ (.A(\registers[22][0] ),
    .B(\registers[23][0] ),
    .S(_01874_),
    .Z(_01875_));
 OAI22_X1 _08086_ (.A1(_01866_),
    .A2(_01870_),
    .B1(_01873_),
    .B2(_01875_),
    .ZN(_01876_));
 BUF_X8 _08087_ (.A(_01867_),
    .Z(_01877_));
 BUF_X4 _08088_ (.A(_01877_),
    .Z(_01878_));
 MUX2_X1 _08089_ (.A(\registers[18][0] ),
    .B(\registers[19][0] ),
    .S(_01878_),
    .Z(_01879_));
 INV_X1 _08090_ (.A(_01879_),
    .ZN(_01880_));
 BUF_X16 _08091_ (.A(_01862_),
    .Z(_01881_));
 INV_X4 _08092_ (.A(_01881_),
    .ZN(_01882_));
 NOR2_X4 _08093_ (.A1(_01882_),
    .A2(_01863_),
    .ZN(_01883_));
 BUF_X4 _08094_ (.A(_01883_),
    .Z(_01884_));
 AOI21_X2 _08095_ (.A(_01876_),
    .B1(_01880_),
    .B2(_01884_),
    .ZN(_01885_));
 CLKBUF_X2 _08096_ (.A(read_addr1[3]),
    .Z(_01886_));
 BUF_X4 _08097_ (.A(_01886_),
    .Z(_01887_));
 BUF_X16 _08098_ (.A(_01881_),
    .Z(_01888_));
 INV_X4 _08099_ (.A(_01863_),
    .ZN(_01889_));
 NOR2_X2 _08100_ (.A1(_01888_),
    .A2(_01889_),
    .ZN(_01890_));
 CLKBUF_X3 _08101_ (.A(_01890_),
    .Z(_01891_));
 BUF_X4 _08102_ (.A(_01868_),
    .Z(_01892_));
 MUX2_X1 _08103_ (.A(\registers[20][0] ),
    .B(\registers[21][0] ),
    .S(_01892_),
    .Z(_01893_));
 INV_X1 _08104_ (.A(_01893_),
    .ZN(_01894_));
 AOI21_X1 _08105_ (.A(_01887_),
    .B1(_01891_),
    .B2(_01894_),
    .ZN(_01895_));
 MUX2_X1 _08106_ (.A(\registers[28][0] ),
    .B(\registers[30][0] ),
    .S(_01881_),
    .Z(_01896_));
 MUX2_X1 _08107_ (.A(\registers[29][0] ),
    .B(\registers[31][0] ),
    .S(_01881_),
    .Z(_01897_));
 BUF_X4 _08108_ (.A(_01867_),
    .Z(_01898_));
 BUF_X4 _08109_ (.A(_01898_),
    .Z(_01899_));
 MUX2_X1 _08110_ (.A(_01896_),
    .B(_01897_),
    .S(_01899_),
    .Z(_01900_));
 MUX2_X1 _08111_ (.A(\registers[24][0] ),
    .B(\registers[26][0] ),
    .S(_01881_),
    .Z(_01901_));
 MUX2_X1 _08112_ (.A(\registers[25][0] ),
    .B(\registers[27][0] ),
    .S(_01881_),
    .Z(_01902_));
 MUX2_X1 _08113_ (.A(_01901_),
    .B(_01902_),
    .S(_01899_),
    .Z(_01903_));
 BUF_X4 _08114_ (.A(_01889_),
    .Z(_01904_));
 MUX2_X1 _08115_ (.A(_01900_),
    .B(_01903_),
    .S(_01904_),
    .Z(_01905_));
 BUF_X4 _08116_ (.A(_01887_),
    .Z(_01906_));
 AOI221_X2 _08117_ (.A(_01860_),
    .B1(_01885_),
    .B2(_01895_),
    .C1(_01905_),
    .C2(_01906_),
    .ZN(_01907_));
 AND2_X1 _08118_ (.A1(net1),
    .A2(_01095_),
    .ZN(_01908_));
 CLKBUF_X2 _08119_ (.A(_01908_),
    .Z(_01909_));
 CLKBUF_X3 _08120_ (.A(_01909_),
    .Z(_01910_));
 OR2_X1 _08121_ (.A1(_01886_),
    .A2(_01858_),
    .ZN(_01911_));
 BUF_X4 _08122_ (.A(_01911_),
    .Z(_01912_));
 BUF_X4 _08123_ (.A(_01866_),
    .Z(_01913_));
 BUF_X4 _08124_ (.A(_01869_),
    .Z(_01914_));
 MUX2_X1 _08125_ (.A(\registers[0][0] ),
    .B(\registers[1][0] ),
    .S(_01914_),
    .Z(_01915_));
 NOR2_X1 _08126_ (.A1(_01913_),
    .A2(_01915_),
    .ZN(_01916_));
 BUF_X4 _08127_ (.A(_01882_),
    .Z(_01917_));
 BUF_X4 _08128_ (.A(_01863_),
    .Z(_01918_));
 MUX2_X1 _08129_ (.A(\registers[2][0] ),
    .B(\registers[3][0] ),
    .S(_01878_),
    .Z(_01919_));
 NOR3_X1 _08130_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_01919_),
    .ZN(_01920_));
 BUF_X4 _08131_ (.A(_01888_),
    .Z(_01921_));
 MUX2_X1 _08132_ (.A(\registers[4][0] ),
    .B(\registers[5][0] ),
    .S(_01892_),
    .Z(_01922_));
 NOR3_X1 _08133_ (.A1(_01921_),
    .A2(_01904_),
    .A3(_01922_),
    .ZN(_01923_));
 BUF_X4 _08134_ (.A(_01873_),
    .Z(_01924_));
 BUF_X4 _08135_ (.A(_01898_),
    .Z(_01925_));
 MUX2_X1 _08136_ (.A(\registers[6][0] ),
    .B(\registers[7][0] ),
    .S(_01925_),
    .Z(_01926_));
 NOR2_X1 _08137_ (.A1(_01924_),
    .A2(_01926_),
    .ZN(_01927_));
 NOR4_X1 _08138_ (.A1(_01916_),
    .A2(_01920_),
    .A3(_01923_),
    .A4(_01927_),
    .ZN(_01928_));
 MUX2_X1 _08139_ (.A(\registers[12][0] ),
    .B(\registers[14][0] ),
    .S(_01888_),
    .Z(_01929_));
 MUX2_X1 _08140_ (.A(\registers[13][0] ),
    .B(\registers[15][0] ),
    .S(_01888_),
    .Z(_01930_));
 BUF_X4 _08141_ (.A(_01878_),
    .Z(_01931_));
 MUX2_X1 _08142_ (.A(_01929_),
    .B(_01930_),
    .S(_01931_),
    .Z(_01932_));
 MUX2_X1 _08143_ (.A(\registers[8][0] ),
    .B(\registers[10][0] ),
    .S(_01888_),
    .Z(_01933_));
 MUX2_X1 _08144_ (.A(\registers[9][0] ),
    .B(\registers[11][0] ),
    .S(_01888_),
    .Z(_01934_));
 MUX2_X1 _08145_ (.A(_01933_),
    .B(_01934_),
    .S(_01931_),
    .Z(_01935_));
 BUF_X4 _08146_ (.A(_01904_),
    .Z(_01936_));
 MUX2_X1 _08147_ (.A(_01932_),
    .B(_01935_),
    .S(_01936_),
    .Z(_01937_));
 NAND2_X1 _08148_ (.A1(_01887_),
    .A2(_01859_),
    .ZN(_01938_));
 CLKBUF_X3 _08149_ (.A(_01938_),
    .Z(_01939_));
 OAI221_X1 _08150_ (.A(_01910_),
    .B1(_01912_),
    .B2(_01928_),
    .C1(_01937_),
    .C2(_01939_),
    .ZN(_01940_));
 INV_X1 _08151_ (.A(net1),
    .ZN(_01941_));
 NAND2_X2 _08152_ (.A1(_01941_),
    .A2(_01416_),
    .ZN(_01942_));
 INV_X1 _08153_ (.A(net5),
    .ZN(_01943_));
 OAI22_X1 _08154_ (.A1(_01907_),
    .A2(_01940_),
    .B1(_01942_),
    .B2(_01943_),
    .ZN(_00329_));
 INV_X1 _08155_ (.A(net6),
    .ZN(_01944_));
 CLKBUF_X3 _08156_ (.A(_01942_),
    .Z(_01945_));
 BUF_X4 _08157_ (.A(_01858_),
    .Z(_01946_));
 BUF_X4 _08158_ (.A(_01867_),
    .Z(_01947_));
 MUX2_X1 _08159_ (.A(\registers[0][10] ),
    .B(\registers[1][10] ),
    .S(_01947_),
    .Z(_01948_));
 MUX2_X1 _08160_ (.A(\registers[6][10] ),
    .B(\registers[7][10] ),
    .S(_01874_),
    .Z(_01949_));
 OAI22_X2 _08161_ (.A1(_01866_),
    .A2(_01948_),
    .B1(_01949_),
    .B2(_01873_),
    .ZN(_01950_));
 BUF_X4 _08162_ (.A(_01877_),
    .Z(_01951_));
 MUX2_X1 _08163_ (.A(\registers[2][10] ),
    .B(\registers[3][10] ),
    .S(_01951_),
    .Z(_01952_));
 INV_X1 _08164_ (.A(_01952_),
    .ZN(_01953_));
 AOI21_X2 _08165_ (.A(_01950_),
    .B1(_01953_),
    .B2(_01884_),
    .ZN(_01954_));
 BUF_X4 _08166_ (.A(_01868_),
    .Z(_01955_));
 MUX2_X1 _08167_ (.A(\registers[4][10] ),
    .B(\registers[5][10] ),
    .S(_01955_),
    .Z(_01956_));
 INV_X1 _08168_ (.A(_01956_),
    .ZN(_01957_));
 AOI21_X1 _08169_ (.A(_01887_),
    .B1(_01891_),
    .B2(_01957_),
    .ZN(_01958_));
 BUF_X8 _08170_ (.A(_01861_),
    .Z(_01959_));
 BUF_X4 _08171_ (.A(_01959_),
    .Z(_01960_));
 MUX2_X1 _08172_ (.A(\registers[12][10] ),
    .B(\registers[14][10] ),
    .S(_01960_),
    .Z(_01961_));
 BUF_X4 _08173_ (.A(_01959_),
    .Z(_01962_));
 MUX2_X1 _08174_ (.A(\registers[13][10] ),
    .B(\registers[15][10] ),
    .S(_01962_),
    .Z(_01963_));
 BUF_X4 _08175_ (.A(_01877_),
    .Z(_01964_));
 MUX2_X1 _08176_ (.A(_01961_),
    .B(_01963_),
    .S(_01964_),
    .Z(_01965_));
 BUF_X4 _08177_ (.A(_01959_),
    .Z(_01966_));
 MUX2_X1 _08178_ (.A(\registers[8][10] ),
    .B(\registers[10][10] ),
    .S(_01966_),
    .Z(_01967_));
 BUF_X4 _08179_ (.A(_01861_),
    .Z(_01968_));
 MUX2_X1 _08180_ (.A(\registers[9][10] ),
    .B(\registers[11][10] ),
    .S(_01968_),
    .Z(_01969_));
 MUX2_X1 _08181_ (.A(_01967_),
    .B(_01969_),
    .S(_01878_),
    .Z(_01970_));
 MUX2_X1 _08182_ (.A(_01965_),
    .B(_01970_),
    .S(_01904_),
    .Z(_01971_));
 AOI221_X2 _08183_ (.A(_01946_),
    .B1(_01954_),
    .B2(_01958_),
    .C1(_01971_),
    .C2(_01906_),
    .ZN(_01972_));
 NAND2_X1 _08184_ (.A1(_01887_),
    .A2(_01858_),
    .ZN(_01973_));
 CLKBUF_X3 _08185_ (.A(_01973_),
    .Z(_01974_));
 BUF_X8 _08186_ (.A(_01862_),
    .Z(_01975_));
 MUX2_X1 _08187_ (.A(\registers[28][10] ),
    .B(\registers[30][10] ),
    .S(_01975_),
    .Z(_01976_));
 BUF_X8 _08188_ (.A(_01862_),
    .Z(_01977_));
 MUX2_X1 _08189_ (.A(\registers[29][10] ),
    .B(\registers[31][10] ),
    .S(_01977_),
    .Z(_01978_));
 BUF_X4 _08190_ (.A(_01869_),
    .Z(_01979_));
 MUX2_X1 _08191_ (.A(_01976_),
    .B(_01978_),
    .S(_01979_),
    .Z(_01980_));
 BUF_X8 _08192_ (.A(_01862_),
    .Z(_01981_));
 MUX2_X1 _08193_ (.A(\registers[24][10] ),
    .B(\registers[26][10] ),
    .S(_01981_),
    .Z(_01982_));
 BUF_X4 _08194_ (.A(_01871_),
    .Z(_01983_));
 MUX2_X1 _08195_ (.A(\registers[25][10] ),
    .B(\registers[27][10] ),
    .S(_01983_),
    .Z(_01984_));
 MUX2_X1 _08196_ (.A(_01982_),
    .B(_01984_),
    .S(_01914_),
    .Z(_01985_));
 BUF_X4 _08197_ (.A(_01889_),
    .Z(_01986_));
 BUF_X4 _08198_ (.A(_01986_),
    .Z(_01987_));
 MUX2_X1 _08199_ (.A(_01980_),
    .B(_01985_),
    .S(_01987_),
    .Z(_01988_));
 OR2_X1 _08200_ (.A1(_01887_),
    .A2(_01859_),
    .ZN(_01989_));
 CLKBUF_X3 _08201_ (.A(_01989_),
    .Z(_01990_));
 MUX2_X1 _08202_ (.A(\registers[16][10] ),
    .B(\registers[17][10] ),
    .S(_01914_),
    .Z(_01991_));
 NOR2_X1 _08203_ (.A1(_01913_),
    .A2(_01991_),
    .ZN(_01992_));
 MUX2_X1 _08204_ (.A(\registers[18][10] ),
    .B(\registers[19][10] ),
    .S(_01899_),
    .Z(_01993_));
 NOR3_X1 _08205_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_01993_),
    .ZN(_01994_));
 BUF_X4 _08206_ (.A(_01877_),
    .Z(_01995_));
 MUX2_X1 _08207_ (.A(\registers[20][10] ),
    .B(\registers[21][10] ),
    .S(_01995_),
    .Z(_01996_));
 NOR3_X1 _08208_ (.A1(_01921_),
    .A2(_01904_),
    .A3(_01996_),
    .ZN(_01997_));
 MUX2_X1 _08209_ (.A(\registers[22][10] ),
    .B(\registers[23][10] ),
    .S(_01899_),
    .Z(_01998_));
 NOR2_X1 _08210_ (.A1(_01924_),
    .A2(_01998_),
    .ZN(_01999_));
 NOR4_X1 _08211_ (.A1(_01992_),
    .A2(_01994_),
    .A3(_01997_),
    .A4(_01999_),
    .ZN(_02000_));
 OAI221_X1 _08212_ (.A(_01910_),
    .B1(_01974_),
    .B2(_01988_),
    .C1(_01990_),
    .C2(_02000_),
    .ZN(_02001_));
 OAI22_X1 _08213_ (.A1(_01944_),
    .A2(_01945_),
    .B1(_01972_),
    .B2(_02001_),
    .ZN(_00330_));
 INV_X1 _08214_ (.A(net7),
    .ZN(_02002_));
 MUX2_X1 _08215_ (.A(\registers[0][11] ),
    .B(\registers[1][11] ),
    .S(_01947_),
    .Z(_02003_));
 MUX2_X1 _08216_ (.A(\registers[6][11] ),
    .B(\registers[7][11] ),
    .S(_01874_),
    .Z(_02004_));
 OAI22_X1 _08217_ (.A1(_01866_),
    .A2(_02003_),
    .B1(_02004_),
    .B2(_01873_),
    .ZN(_02005_));
 MUX2_X1 _08218_ (.A(\registers[2][11] ),
    .B(\registers[3][11] ),
    .S(_01951_),
    .Z(_02006_));
 INV_X1 _08219_ (.A(_02006_),
    .ZN(_02007_));
 AOI21_X1 _08220_ (.A(_02005_),
    .B1(_02007_),
    .B2(_01884_),
    .ZN(_02008_));
 CLKBUF_X3 _08221_ (.A(_01886_),
    .Z(_02009_));
 MUX2_X1 _08222_ (.A(\registers[4][11] ),
    .B(\registers[5][11] ),
    .S(_01955_),
    .Z(_02010_));
 INV_X1 _08223_ (.A(_02010_),
    .ZN(_02011_));
 AOI21_X1 _08224_ (.A(_02009_),
    .B1(_01891_),
    .B2(_02011_),
    .ZN(_02012_));
 MUX2_X1 _08225_ (.A(\registers[12][11] ),
    .B(\registers[14][11] ),
    .S(_01960_),
    .Z(_02013_));
 MUX2_X1 _08226_ (.A(\registers[13][11] ),
    .B(\registers[15][11] ),
    .S(_01962_),
    .Z(_02014_));
 MUX2_X1 _08227_ (.A(_02013_),
    .B(_02014_),
    .S(_01964_),
    .Z(_02015_));
 MUX2_X1 _08228_ (.A(\registers[8][11] ),
    .B(\registers[10][11] ),
    .S(_01966_),
    .Z(_02016_));
 MUX2_X1 _08229_ (.A(\registers[9][11] ),
    .B(\registers[11][11] ),
    .S(_01968_),
    .Z(_02017_));
 MUX2_X1 _08230_ (.A(_02016_),
    .B(_02017_),
    .S(_01878_),
    .Z(_02018_));
 MUX2_X2 _08231_ (.A(_02015_),
    .B(_02018_),
    .S(_01904_),
    .Z(_02019_));
 AOI221_X2 _08232_ (.A(_01946_),
    .B1(_02008_),
    .B2(_02012_),
    .C1(_02019_),
    .C2(_01906_),
    .ZN(_02020_));
 MUX2_X1 _08233_ (.A(\registers[28][11] ),
    .B(\registers[30][11] ),
    .S(_01975_),
    .Z(_02021_));
 MUX2_X1 _08234_ (.A(\registers[29][11] ),
    .B(\registers[31][11] ),
    .S(_01977_),
    .Z(_02022_));
 MUX2_X1 _08235_ (.A(_02021_),
    .B(_02022_),
    .S(_01979_),
    .Z(_02023_));
 MUX2_X1 _08236_ (.A(\registers[24][11] ),
    .B(\registers[26][11] ),
    .S(_01981_),
    .Z(_02024_));
 MUX2_X1 _08237_ (.A(\registers[25][11] ),
    .B(\registers[27][11] ),
    .S(_01983_),
    .Z(_02025_));
 MUX2_X1 _08238_ (.A(_02024_),
    .B(_02025_),
    .S(_01914_),
    .Z(_02026_));
 MUX2_X1 _08239_ (.A(_02023_),
    .B(_02026_),
    .S(_01987_),
    .Z(_02027_));
 BUF_X4 _08240_ (.A(_01866_),
    .Z(_02028_));
 BUF_X4 _08241_ (.A(_01868_),
    .Z(_02029_));
 BUF_X4 _08242_ (.A(_02029_),
    .Z(_02030_));
 MUX2_X1 _08243_ (.A(\registers[16][11] ),
    .B(\registers[17][11] ),
    .S(_02030_),
    .Z(_02031_));
 NOR2_X1 _08244_ (.A1(_02028_),
    .A2(_02031_),
    .ZN(_02032_));
 CLKBUF_X3 _08245_ (.A(_01882_),
    .Z(_02033_));
 CLKBUF_X3 _08246_ (.A(_01863_),
    .Z(_02034_));
 BUF_X4 _08247_ (.A(_01947_),
    .Z(_02035_));
 MUX2_X1 _08248_ (.A(\registers[18][11] ),
    .B(\registers[19][11] ),
    .S(_02035_),
    .Z(_02036_));
 NOR3_X1 _08249_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02036_),
    .ZN(_02037_));
 CLKBUF_X3 _08250_ (.A(_01888_),
    .Z(_02038_));
 BUF_X4 _08251_ (.A(_01889_),
    .Z(_02039_));
 MUX2_X1 _08252_ (.A(\registers[20][11] ),
    .B(\registers[21][11] ),
    .S(_01925_),
    .Z(_02040_));
 NOR3_X1 _08253_ (.A1(_02038_),
    .A2(_02039_),
    .A3(_02040_),
    .ZN(_02041_));
 BUF_X4 _08254_ (.A(_01873_),
    .Z(_02042_));
 BUF_X4 _08255_ (.A(_01947_),
    .Z(_02043_));
 MUX2_X1 _08256_ (.A(\registers[22][11] ),
    .B(\registers[23][11] ),
    .S(_02043_),
    .Z(_02044_));
 NOR2_X1 _08257_ (.A1(_02042_),
    .A2(_02044_),
    .ZN(_02045_));
 NOR4_X2 _08258_ (.A1(_02032_),
    .A2(_02037_),
    .A3(_02041_),
    .A4(_02045_),
    .ZN(_02046_));
 OAI221_X1 _08259_ (.A(_01910_),
    .B1(_01974_),
    .B2(_02027_),
    .C1(_02046_),
    .C2(_01990_),
    .ZN(_02047_));
 OAI22_X1 _08260_ (.A1(_02002_),
    .A2(_01945_),
    .B1(_02020_),
    .B2(_02047_),
    .ZN(_00331_));
 INV_X1 _08261_ (.A(net8),
    .ZN(_02048_));
 MUX2_X1 _08262_ (.A(\registers[0][12] ),
    .B(\registers[1][12] ),
    .S(_01947_),
    .Z(_02049_));
 MUX2_X1 _08263_ (.A(\registers[6][12] ),
    .B(\registers[7][12] ),
    .S(_01874_),
    .Z(_02050_));
 OAI22_X1 _08264_ (.A1(_01866_),
    .A2(_02049_),
    .B1(_02050_),
    .B2(_01873_),
    .ZN(_02051_));
 BUF_X4 _08265_ (.A(_01877_),
    .Z(_02052_));
 MUX2_X1 _08266_ (.A(\registers[2][12] ),
    .B(\registers[3][12] ),
    .S(_02052_),
    .Z(_02053_));
 INV_X1 _08267_ (.A(_02053_),
    .ZN(_02054_));
 AOI21_X1 _08268_ (.A(_02051_),
    .B1(_02054_),
    .B2(_01884_),
    .ZN(_02055_));
 MUX2_X1 _08269_ (.A(\registers[4][12] ),
    .B(\registers[5][12] ),
    .S(_01955_),
    .Z(_02056_));
 INV_X1 _08270_ (.A(_02056_),
    .ZN(_02057_));
 AOI21_X1 _08271_ (.A(_02009_),
    .B1(_01891_),
    .B2(_02057_),
    .ZN(_02058_));
 MUX2_X1 _08272_ (.A(\registers[12][12] ),
    .B(\registers[14][12] ),
    .S(_01960_),
    .Z(_02059_));
 MUX2_X1 _08273_ (.A(\registers[13][12] ),
    .B(\registers[15][12] ),
    .S(_01962_),
    .Z(_02060_));
 MUX2_X1 _08274_ (.A(_02059_),
    .B(_02060_),
    .S(_01964_),
    .Z(_02061_));
 MUX2_X1 _08275_ (.A(\registers[8][12] ),
    .B(\registers[10][12] ),
    .S(_01966_),
    .Z(_02062_));
 MUX2_X1 _08276_ (.A(\registers[9][12] ),
    .B(\registers[11][12] ),
    .S(_01968_),
    .Z(_02063_));
 MUX2_X1 _08277_ (.A(_02062_),
    .B(_02063_),
    .S(_01878_),
    .Z(_02064_));
 MUX2_X1 _08278_ (.A(_02061_),
    .B(_02064_),
    .S(_01904_),
    .Z(_02065_));
 AOI221_X2 _08279_ (.A(_01946_),
    .B1(_02055_),
    .B2(_02058_),
    .C1(_02065_),
    .C2(_01906_),
    .ZN(_02066_));
 MUX2_X1 _08280_ (.A(\registers[28][12] ),
    .B(\registers[30][12] ),
    .S(_01975_),
    .Z(_02067_));
 MUX2_X1 _08281_ (.A(\registers[29][12] ),
    .B(\registers[31][12] ),
    .S(_01977_),
    .Z(_02068_));
 MUX2_X1 _08282_ (.A(_02067_),
    .B(_02068_),
    .S(_01979_),
    .Z(_02069_));
 MUX2_X1 _08283_ (.A(\registers[24][12] ),
    .B(\registers[26][12] ),
    .S(_01981_),
    .Z(_02070_));
 MUX2_X1 _08284_ (.A(\registers[25][12] ),
    .B(\registers[27][12] ),
    .S(_01983_),
    .Z(_02071_));
 MUX2_X1 _08285_ (.A(_02070_),
    .B(_02071_),
    .S(_01914_),
    .Z(_02072_));
 MUX2_X1 _08286_ (.A(_02069_),
    .B(_02072_),
    .S(_01987_),
    .Z(_02073_));
 MUX2_X1 _08287_ (.A(\registers[16][12] ),
    .B(\registers[17][12] ),
    .S(_02030_),
    .Z(_02074_));
 NOR2_X1 _08288_ (.A1(_02028_),
    .A2(_02074_),
    .ZN(_02075_));
 MUX2_X1 _08289_ (.A(\registers[18][12] ),
    .B(\registers[19][12] ),
    .S(_02035_),
    .Z(_02076_));
 NOR3_X1 _08290_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02076_),
    .ZN(_02077_));
 MUX2_X1 _08291_ (.A(\registers[20][12] ),
    .B(\registers[21][12] ),
    .S(_01925_),
    .Z(_02078_));
 NOR3_X1 _08292_ (.A1(_02038_),
    .A2(_02039_),
    .A3(_02078_),
    .ZN(_02079_));
 MUX2_X1 _08293_ (.A(\registers[22][12] ),
    .B(\registers[23][12] ),
    .S(_02043_),
    .Z(_02080_));
 NOR2_X1 _08294_ (.A1(_02042_),
    .A2(_02080_),
    .ZN(_02081_));
 NOR4_X2 _08295_ (.A1(_02075_),
    .A2(_02077_),
    .A3(_02079_),
    .A4(_02081_),
    .ZN(_02082_));
 OAI221_X1 _08296_ (.A(_01910_),
    .B1(_01974_),
    .B2(_02073_),
    .C1(_02082_),
    .C2(_01990_),
    .ZN(_02083_));
 OAI22_X1 _08297_ (.A1(_02048_),
    .A2(_01945_),
    .B1(_02066_),
    .B2(_02083_),
    .ZN(_00332_));
 INV_X1 _08298_ (.A(net9),
    .ZN(_02084_));
 MUX2_X1 _08299_ (.A(\registers[0][13] ),
    .B(\registers[1][13] ),
    .S(_01947_),
    .Z(_02085_));
 MUX2_X1 _08300_ (.A(\registers[6][13] ),
    .B(\registers[7][13] ),
    .S(_01874_),
    .Z(_02086_));
 OAI22_X1 _08301_ (.A1(_01866_),
    .A2(_02085_),
    .B1(_02086_),
    .B2(_01873_),
    .ZN(_02087_));
 MUX2_X1 _08302_ (.A(\registers[2][13] ),
    .B(\registers[3][13] ),
    .S(_02052_),
    .Z(_02088_));
 INV_X1 _08303_ (.A(_02088_),
    .ZN(_02089_));
 AOI21_X1 _08304_ (.A(_02087_),
    .B1(_02089_),
    .B2(_01884_),
    .ZN(_02090_));
 MUX2_X1 _08305_ (.A(\registers[4][13] ),
    .B(\registers[5][13] ),
    .S(_01955_),
    .Z(_02091_));
 INV_X1 _08306_ (.A(_02091_),
    .ZN(_02092_));
 AOI21_X1 _08307_ (.A(_02009_),
    .B1(_01891_),
    .B2(_02092_),
    .ZN(_02093_));
 BUF_X4 _08308_ (.A(_01959_),
    .Z(_02094_));
 MUX2_X1 _08309_ (.A(\registers[12][13] ),
    .B(\registers[14][13] ),
    .S(_02094_),
    .Z(_02095_));
 MUX2_X1 _08310_ (.A(\registers[13][13] ),
    .B(\registers[15][13] ),
    .S(_01962_),
    .Z(_02096_));
 MUX2_X1 _08311_ (.A(_02095_),
    .B(_02096_),
    .S(_01964_),
    .Z(_02097_));
 MUX2_X1 _08312_ (.A(\registers[8][13] ),
    .B(\registers[10][13] ),
    .S(_01966_),
    .Z(_02098_));
 MUX2_X1 _08313_ (.A(\registers[9][13] ),
    .B(\registers[11][13] ),
    .S(_01968_),
    .Z(_02099_));
 MUX2_X1 _08314_ (.A(_02098_),
    .B(_02099_),
    .S(_01878_),
    .Z(_02100_));
 MUX2_X1 _08315_ (.A(_02097_),
    .B(_02100_),
    .S(_01904_),
    .Z(_02101_));
 AOI221_X1 _08316_ (.A(_01946_),
    .B1(_02090_),
    .B2(_02093_),
    .C1(_02101_),
    .C2(_01906_),
    .ZN(_02102_));
 MUX2_X1 _08317_ (.A(\registers[28][13] ),
    .B(\registers[30][13] ),
    .S(_01975_),
    .Z(_02103_));
 MUX2_X1 _08318_ (.A(\registers[29][13] ),
    .B(\registers[31][13] ),
    .S(_01977_),
    .Z(_02104_));
 MUX2_X1 _08319_ (.A(_02103_),
    .B(_02104_),
    .S(_01979_),
    .Z(_02105_));
 MUX2_X1 _08320_ (.A(\registers[24][13] ),
    .B(\registers[26][13] ),
    .S(_01981_),
    .Z(_02106_));
 MUX2_X1 _08321_ (.A(\registers[25][13] ),
    .B(\registers[27][13] ),
    .S(_01983_),
    .Z(_02107_));
 MUX2_X1 _08322_ (.A(_02106_),
    .B(_02107_),
    .S(_01914_),
    .Z(_02108_));
 MUX2_X1 _08323_ (.A(_02105_),
    .B(_02108_),
    .S(_01987_),
    .Z(_02109_));
 MUX2_X1 _08324_ (.A(\registers[16][13] ),
    .B(\registers[17][13] ),
    .S(_02030_),
    .Z(_02110_));
 NOR2_X1 _08325_ (.A1(_02028_),
    .A2(_02110_),
    .ZN(_02111_));
 MUX2_X1 _08326_ (.A(\registers[18][13] ),
    .B(\registers[19][13] ),
    .S(_02035_),
    .Z(_02112_));
 NOR3_X1 _08327_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02112_),
    .ZN(_02113_));
 MUX2_X1 _08328_ (.A(\registers[20][13] ),
    .B(\registers[21][13] ),
    .S(_01925_),
    .Z(_02114_));
 NOR3_X1 _08329_ (.A1(_02038_),
    .A2(_02039_),
    .A3(_02114_),
    .ZN(_02115_));
 MUX2_X1 _08330_ (.A(\registers[22][13] ),
    .B(\registers[23][13] ),
    .S(_02043_),
    .Z(_02116_));
 NOR2_X1 _08331_ (.A1(_02042_),
    .A2(_02116_),
    .ZN(_02117_));
 NOR4_X2 _08332_ (.A1(_02111_),
    .A2(_02113_),
    .A3(_02115_),
    .A4(_02117_),
    .ZN(_02118_));
 OAI221_X1 _08333_ (.A(_01910_),
    .B1(_01974_),
    .B2(_02109_),
    .C1(_02118_),
    .C2(_01990_),
    .ZN(_02119_));
 OAI22_X1 _08334_ (.A1(_02084_),
    .A2(_01945_),
    .B1(_02102_),
    .B2(_02119_),
    .ZN(_00333_));
 INV_X1 _08335_ (.A(net10),
    .ZN(_02120_));
 BUF_X4 _08336_ (.A(_01865_),
    .Z(_02121_));
 MUX2_X1 _08337_ (.A(\registers[16][14] ),
    .B(\registers[17][14] ),
    .S(_01947_),
    .Z(_02122_));
 BUF_X4 _08338_ (.A(_01867_),
    .Z(_02123_));
 MUX2_X1 _08339_ (.A(\registers[22][14] ),
    .B(\registers[23][14] ),
    .S(_02123_),
    .Z(_02124_));
 BUF_X4 _08340_ (.A(_01872_),
    .Z(_02125_));
 OAI22_X1 _08341_ (.A1(_02121_),
    .A2(_02122_),
    .B1(_02124_),
    .B2(_02125_),
    .ZN(_02126_));
 MUX2_X1 _08342_ (.A(\registers[18][14] ),
    .B(\registers[19][14] ),
    .S(_02052_),
    .Z(_02127_));
 INV_X1 _08343_ (.A(_02127_),
    .ZN(_02128_));
 AOI21_X2 _08344_ (.A(_02126_),
    .B1(_02128_),
    .B2(_01884_),
    .ZN(_02129_));
 MUX2_X1 _08345_ (.A(\registers[20][14] ),
    .B(\registers[21][14] ),
    .S(_01955_),
    .Z(_02130_));
 INV_X1 _08346_ (.A(_02130_),
    .ZN(_02131_));
 AOI21_X1 _08347_ (.A(_02009_),
    .B1(_01891_),
    .B2(_02131_),
    .ZN(_02132_));
 MUX2_X1 _08348_ (.A(\registers[28][14] ),
    .B(\registers[30][14] ),
    .S(_02094_),
    .Z(_02133_));
 BUF_X4 _08349_ (.A(_01959_),
    .Z(_02134_));
 MUX2_X1 _08350_ (.A(\registers[29][14] ),
    .B(\registers[31][14] ),
    .S(_02134_),
    .Z(_02135_));
 BUF_X4 _08351_ (.A(_01877_),
    .Z(_02136_));
 MUX2_X1 _08352_ (.A(_02133_),
    .B(_02135_),
    .S(_02136_),
    .Z(_02137_));
 MUX2_X1 _08353_ (.A(\registers[24][14] ),
    .B(\registers[26][14] ),
    .S(_01966_),
    .Z(_02138_));
 MUX2_X1 _08354_ (.A(\registers[25][14] ),
    .B(\registers[27][14] ),
    .S(_01968_),
    .Z(_02139_));
 MUX2_X1 _08355_ (.A(_02138_),
    .B(_02139_),
    .S(_01878_),
    .Z(_02140_));
 BUF_X4 _08356_ (.A(_01889_),
    .Z(_02141_));
 MUX2_X1 _08357_ (.A(_02137_),
    .B(_02140_),
    .S(_02141_),
    .Z(_02142_));
 AOI221_X2 _08358_ (.A(_01860_),
    .B1(_02129_),
    .B2(_02132_),
    .C1(_02142_),
    .C2(_01906_),
    .ZN(_02143_));
 BUF_X4 _08359_ (.A(_01869_),
    .Z(_02144_));
 MUX2_X1 _08360_ (.A(\registers[0][14] ),
    .B(\registers[1][14] ),
    .S(_02144_),
    .Z(_02145_));
 NOR2_X1 _08361_ (.A1(_01913_),
    .A2(_02145_),
    .ZN(_02146_));
 MUX2_X1 _08362_ (.A(\registers[2][14] ),
    .B(\registers[3][14] ),
    .S(_01892_),
    .Z(_02147_));
 NOR3_X1 _08363_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_02147_),
    .ZN(_02148_));
 BUF_X4 _08364_ (.A(_01889_),
    .Z(_02149_));
 BUF_X4 _08365_ (.A(_01868_),
    .Z(_02150_));
 MUX2_X1 _08366_ (.A(\registers[4][14] ),
    .B(\registers[5][14] ),
    .S(_02150_),
    .Z(_02151_));
 NOR3_X1 _08367_ (.A1(_01921_),
    .A2(_02149_),
    .A3(_02151_),
    .ZN(_02152_));
 MUX2_X1 _08368_ (.A(\registers[6][14] ),
    .B(\registers[7][14] ),
    .S(_01995_),
    .Z(_02153_));
 NOR2_X1 _08369_ (.A1(_01924_),
    .A2(_02153_),
    .ZN(_02154_));
 NOR4_X1 _08370_ (.A1(_02146_),
    .A2(_02148_),
    .A3(_02152_),
    .A4(_02154_),
    .ZN(_02155_));
 BUF_X4 _08371_ (.A(_01968_),
    .Z(_02156_));
 MUX2_X1 _08372_ (.A(\registers[12][14] ),
    .B(\registers[14][14] ),
    .S(_02156_),
    .Z(_02157_));
 BUF_X4 _08373_ (.A(_01968_),
    .Z(_02158_));
 MUX2_X1 _08374_ (.A(\registers[13][14] ),
    .B(\registers[15][14] ),
    .S(_02158_),
    .Z(_02159_));
 BUF_X4 _08375_ (.A(_01878_),
    .Z(_02160_));
 MUX2_X1 _08376_ (.A(_02157_),
    .B(_02159_),
    .S(_02160_),
    .Z(_02161_));
 BUF_X4 _08377_ (.A(_01968_),
    .Z(_02162_));
 MUX2_X1 _08378_ (.A(\registers[8][14] ),
    .B(\registers[10][14] ),
    .S(_02162_),
    .Z(_02163_));
 BUF_X4 _08379_ (.A(_01968_),
    .Z(_02164_));
 MUX2_X1 _08380_ (.A(\registers[9][14] ),
    .B(\registers[11][14] ),
    .S(_02164_),
    .Z(_02165_));
 MUX2_X1 _08381_ (.A(_02163_),
    .B(_02165_),
    .S(_01931_),
    .Z(_02166_));
 MUX2_X1 _08382_ (.A(_02161_),
    .B(_02166_),
    .S(_01936_),
    .Z(_02167_));
 OAI221_X1 _08383_ (.A(_01910_),
    .B1(_01912_),
    .B2(_02155_),
    .C1(_02167_),
    .C2(_01939_),
    .ZN(_02168_));
 OAI22_X1 _08384_ (.A1(_02120_),
    .A2(_01945_),
    .B1(_02143_),
    .B2(_02168_),
    .ZN(_00334_));
 INV_X1 _08385_ (.A(net11),
    .ZN(_02169_));
 MUX2_X1 _08386_ (.A(\registers[0][15] ),
    .B(\registers[1][15] ),
    .S(_01947_),
    .Z(_02170_));
 MUX2_X1 _08387_ (.A(\registers[6][15] ),
    .B(\registers[7][15] ),
    .S(_02123_),
    .Z(_02171_));
 OAI22_X1 _08388_ (.A1(_02121_),
    .A2(_02170_),
    .B1(_02171_),
    .B2(_02125_),
    .ZN(_02172_));
 MUX2_X1 _08389_ (.A(\registers[2][15] ),
    .B(\registers[3][15] ),
    .S(_02052_),
    .Z(_02173_));
 INV_X1 _08390_ (.A(_02173_),
    .ZN(_02174_));
 AOI21_X1 _08391_ (.A(_02172_),
    .B1(_02174_),
    .B2(_01884_),
    .ZN(_02175_));
 MUX2_X1 _08392_ (.A(\registers[4][15] ),
    .B(\registers[5][15] ),
    .S(_01955_),
    .Z(_02176_));
 INV_X1 _08393_ (.A(_02176_),
    .ZN(_02177_));
 AOI21_X1 _08394_ (.A(_02009_),
    .B1(_01891_),
    .B2(_02177_),
    .ZN(_02178_));
 MUX2_X1 _08395_ (.A(\registers[12][15] ),
    .B(\registers[14][15] ),
    .S(_02094_),
    .Z(_02179_));
 MUX2_X1 _08396_ (.A(\registers[13][15] ),
    .B(\registers[15][15] ),
    .S(_02134_),
    .Z(_02180_));
 MUX2_X1 _08397_ (.A(_02179_),
    .B(_02180_),
    .S(_02136_),
    .Z(_02181_));
 BUF_X4 _08398_ (.A(_01959_),
    .Z(_02182_));
 MUX2_X1 _08399_ (.A(\registers[8][15] ),
    .B(\registers[10][15] ),
    .S(_02182_),
    .Z(_02183_));
 MUX2_X1 _08400_ (.A(\registers[9][15] ),
    .B(\registers[11][15] ),
    .S(_01968_),
    .Z(_02184_));
 BUF_X4 _08401_ (.A(_01877_),
    .Z(_02185_));
 MUX2_X1 _08402_ (.A(_02183_),
    .B(_02184_),
    .S(_02185_),
    .Z(_02186_));
 MUX2_X2 _08403_ (.A(_02181_),
    .B(_02186_),
    .S(_02141_),
    .Z(_02187_));
 AOI221_X2 _08404_ (.A(_01946_),
    .B1(_02175_),
    .B2(_02178_),
    .C1(_02187_),
    .C2(_01906_),
    .ZN(_02188_));
 MUX2_X1 _08405_ (.A(\registers[28][15] ),
    .B(\registers[30][15] ),
    .S(_01975_),
    .Z(_02189_));
 MUX2_X1 _08406_ (.A(\registers[29][15] ),
    .B(\registers[31][15] ),
    .S(_01977_),
    .Z(_02190_));
 MUX2_X1 _08407_ (.A(_02189_),
    .B(_02190_),
    .S(_01979_),
    .Z(_02191_));
 MUX2_X1 _08408_ (.A(\registers[24][15] ),
    .B(\registers[26][15] ),
    .S(_01981_),
    .Z(_02192_));
 MUX2_X1 _08409_ (.A(\registers[25][15] ),
    .B(\registers[27][15] ),
    .S(_01983_),
    .Z(_02193_));
 MUX2_X1 _08410_ (.A(_02192_),
    .B(_02193_),
    .S(_01914_),
    .Z(_02194_));
 MUX2_X1 _08411_ (.A(_02191_),
    .B(_02194_),
    .S(_01987_),
    .Z(_02195_));
 MUX2_X1 _08412_ (.A(\registers[16][15] ),
    .B(\registers[17][15] ),
    .S(_02030_),
    .Z(_02196_));
 NOR2_X1 _08413_ (.A1(_02028_),
    .A2(_02196_),
    .ZN(_02197_));
 MUX2_X1 _08414_ (.A(\registers[18][15] ),
    .B(\registers[19][15] ),
    .S(_02035_),
    .Z(_02198_));
 NOR3_X1 _08415_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02198_),
    .ZN(_02199_));
 MUX2_X1 _08416_ (.A(\registers[20][15] ),
    .B(\registers[21][15] ),
    .S(_01925_),
    .Z(_02200_));
 NOR3_X1 _08417_ (.A1(_02038_),
    .A2(_02039_),
    .A3(_02200_),
    .ZN(_02201_));
 MUX2_X1 _08418_ (.A(\registers[22][15] ),
    .B(\registers[23][15] ),
    .S(_02043_),
    .Z(_02202_));
 NOR2_X1 _08419_ (.A1(_02042_),
    .A2(_02202_),
    .ZN(_02203_));
 NOR4_X2 _08420_ (.A1(_02197_),
    .A2(_02199_),
    .A3(_02201_),
    .A4(_02203_),
    .ZN(_02204_));
 OAI221_X1 _08421_ (.A(_01910_),
    .B1(_01974_),
    .B2(_02195_),
    .C1(_02204_),
    .C2(_01990_),
    .ZN(_02205_));
 OAI22_X1 _08422_ (.A1(_02169_),
    .A2(_01945_),
    .B1(_02188_),
    .B2(_02205_),
    .ZN(_00335_));
 INV_X1 _08423_ (.A(net12),
    .ZN(_02206_));
 BUF_X4 _08424_ (.A(_01868_),
    .Z(_02207_));
 MUX2_X1 _08425_ (.A(\registers[16][16] ),
    .B(\registers[17][16] ),
    .S(_02207_),
    .Z(_02208_));
 MUX2_X1 _08426_ (.A(\registers[22][16] ),
    .B(\registers[23][16] ),
    .S(_02123_),
    .Z(_02209_));
 OAI22_X1 _08427_ (.A1(_02121_),
    .A2(_02208_),
    .B1(_02209_),
    .B2(_02125_),
    .ZN(_02210_));
 MUX2_X1 _08428_ (.A(\registers[18][16] ),
    .B(\registers[19][16] ),
    .S(_02052_),
    .Z(_02211_));
 INV_X1 _08429_ (.A(_02211_),
    .ZN(_02212_));
 AOI21_X1 _08430_ (.A(_02210_),
    .B1(_02212_),
    .B2(_01884_),
    .ZN(_02213_));
 MUX2_X1 _08431_ (.A(\registers[20][16] ),
    .B(\registers[21][16] ),
    .S(_01955_),
    .Z(_02214_));
 INV_X1 _08432_ (.A(_02214_),
    .ZN(_02215_));
 AOI21_X1 _08433_ (.A(_02009_),
    .B1(_01891_),
    .B2(_02215_),
    .ZN(_02216_));
 MUX2_X1 _08434_ (.A(\registers[28][16] ),
    .B(\registers[30][16] ),
    .S(_02094_),
    .Z(_02217_));
 MUX2_X1 _08435_ (.A(\registers[29][16] ),
    .B(\registers[31][16] ),
    .S(_02134_),
    .Z(_02218_));
 MUX2_X1 _08436_ (.A(_02217_),
    .B(_02218_),
    .S(_02136_),
    .Z(_02219_));
 MUX2_X1 _08437_ (.A(\registers[24][16] ),
    .B(\registers[26][16] ),
    .S(_02182_),
    .Z(_02220_));
 BUF_X4 _08438_ (.A(_01862_),
    .Z(_02221_));
 MUX2_X1 _08439_ (.A(\registers[25][16] ),
    .B(\registers[27][16] ),
    .S(_02221_),
    .Z(_02222_));
 MUX2_X1 _08440_ (.A(_02220_),
    .B(_02222_),
    .S(_02185_),
    .Z(_02223_));
 MUX2_X1 _08441_ (.A(_02219_),
    .B(_02223_),
    .S(_02141_),
    .Z(_02224_));
 AOI221_X1 _08442_ (.A(_01860_),
    .B1(_02213_),
    .B2(_02216_),
    .C1(_02224_),
    .C2(_01906_),
    .ZN(_02225_));
 MUX2_X1 _08443_ (.A(\registers[0][16] ),
    .B(\registers[1][16] ),
    .S(_02144_),
    .Z(_02226_));
 NOR2_X1 _08444_ (.A1(_01913_),
    .A2(_02226_),
    .ZN(_02227_));
 MUX2_X1 _08445_ (.A(\registers[2][16] ),
    .B(\registers[3][16] ),
    .S(_01892_),
    .Z(_02228_));
 NOR3_X1 _08446_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_02228_),
    .ZN(_02229_));
 MUX2_X1 _08447_ (.A(\registers[4][16] ),
    .B(\registers[5][16] ),
    .S(_02150_),
    .Z(_02230_));
 NOR3_X1 _08448_ (.A1(_01921_),
    .A2(_02149_),
    .A3(_02230_),
    .ZN(_02231_));
 MUX2_X1 _08449_ (.A(\registers[6][16] ),
    .B(\registers[7][16] ),
    .S(_01995_),
    .Z(_02232_));
 NOR2_X1 _08450_ (.A1(_01924_),
    .A2(_02232_),
    .ZN(_02233_));
 NOR4_X1 _08451_ (.A1(_02227_),
    .A2(_02229_),
    .A3(_02231_),
    .A4(_02233_),
    .ZN(_02234_));
 MUX2_X1 _08452_ (.A(\registers[12][16] ),
    .B(\registers[14][16] ),
    .S(_02156_),
    .Z(_02235_));
 MUX2_X1 _08453_ (.A(\registers[13][16] ),
    .B(\registers[15][16] ),
    .S(_02158_),
    .Z(_02236_));
 MUX2_X1 _08454_ (.A(_02235_),
    .B(_02236_),
    .S(_02160_),
    .Z(_02237_));
 MUX2_X1 _08455_ (.A(\registers[8][16] ),
    .B(\registers[10][16] ),
    .S(_02162_),
    .Z(_02238_));
 MUX2_X1 _08456_ (.A(\registers[9][16] ),
    .B(\registers[11][16] ),
    .S(_02164_),
    .Z(_02239_));
 MUX2_X1 _08457_ (.A(_02238_),
    .B(_02239_),
    .S(_01931_),
    .Z(_02240_));
 MUX2_X1 _08458_ (.A(_02237_),
    .B(_02240_),
    .S(_01936_),
    .Z(_02241_));
 OAI221_X1 _08459_ (.A(_01910_),
    .B1(_01912_),
    .B2(_02234_),
    .C1(_02241_),
    .C2(_01939_),
    .ZN(_02242_));
 OAI22_X1 _08460_ (.A1(_02206_),
    .A2(_01945_),
    .B1(_02225_),
    .B2(_02242_),
    .ZN(_00336_));
 INV_X1 _08461_ (.A(net13),
    .ZN(_02243_));
 MUX2_X1 _08462_ (.A(\registers[16][17] ),
    .B(\registers[17][17] ),
    .S(_02207_),
    .Z(_02244_));
 MUX2_X1 _08463_ (.A(\registers[22][17] ),
    .B(\registers[23][17] ),
    .S(_02123_),
    .Z(_02245_));
 OAI22_X1 _08464_ (.A1(_02121_),
    .A2(_02244_),
    .B1(_02245_),
    .B2(_02125_),
    .ZN(_02246_));
 MUX2_X1 _08465_ (.A(\registers[18][17] ),
    .B(\registers[19][17] ),
    .S(_02052_),
    .Z(_02247_));
 INV_X1 _08466_ (.A(_02247_),
    .ZN(_02248_));
 AOI21_X2 _08467_ (.A(_02246_),
    .B1(_02248_),
    .B2(_01884_),
    .ZN(_02249_));
 BUF_X4 _08468_ (.A(_01868_),
    .Z(_02250_));
 MUX2_X1 _08469_ (.A(\registers[20][17] ),
    .B(\registers[21][17] ),
    .S(_02250_),
    .Z(_02251_));
 INV_X1 _08470_ (.A(_02251_),
    .ZN(_02252_));
 AOI21_X1 _08471_ (.A(_02009_),
    .B1(_01891_),
    .B2(_02252_),
    .ZN(_02253_));
 MUX2_X1 _08472_ (.A(\registers[28][17] ),
    .B(\registers[30][17] ),
    .S(_02094_),
    .Z(_02254_));
 MUX2_X1 _08473_ (.A(\registers[29][17] ),
    .B(\registers[31][17] ),
    .S(_02134_),
    .Z(_02255_));
 MUX2_X1 _08474_ (.A(_02254_),
    .B(_02255_),
    .S(_02136_),
    .Z(_02256_));
 MUX2_X1 _08475_ (.A(\registers[24][17] ),
    .B(\registers[26][17] ),
    .S(_02182_),
    .Z(_02257_));
 MUX2_X1 _08476_ (.A(\registers[25][17] ),
    .B(\registers[27][17] ),
    .S(_02221_),
    .Z(_02258_));
 MUX2_X1 _08477_ (.A(_02257_),
    .B(_02258_),
    .S(_02185_),
    .Z(_02259_));
 MUX2_X1 _08478_ (.A(_02256_),
    .B(_02259_),
    .S(_02141_),
    .Z(_02260_));
 AOI221_X2 _08479_ (.A(_01860_),
    .B1(_02249_),
    .B2(_02253_),
    .C1(_02260_),
    .C2(_01906_),
    .ZN(_02261_));
 MUX2_X1 _08480_ (.A(\registers[0][17] ),
    .B(\registers[1][17] ),
    .S(_02144_),
    .Z(_02262_));
 NOR2_X1 _08481_ (.A1(_01913_),
    .A2(_02262_),
    .ZN(_02263_));
 MUX2_X1 _08482_ (.A(\registers[2][17] ),
    .B(\registers[3][17] ),
    .S(_01892_),
    .Z(_02264_));
 NOR3_X1 _08483_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_02264_),
    .ZN(_02265_));
 MUX2_X1 _08484_ (.A(\registers[4][17] ),
    .B(\registers[5][17] ),
    .S(_02150_),
    .Z(_02266_));
 NOR3_X1 _08485_ (.A1(_01921_),
    .A2(_02149_),
    .A3(_02266_),
    .ZN(_02267_));
 MUX2_X1 _08486_ (.A(\registers[6][17] ),
    .B(\registers[7][17] ),
    .S(_01951_),
    .Z(_02268_));
 NOR2_X1 _08487_ (.A1(_01924_),
    .A2(_02268_),
    .ZN(_02269_));
 NOR4_X1 _08488_ (.A1(_02263_),
    .A2(_02265_),
    .A3(_02267_),
    .A4(_02269_),
    .ZN(_02270_));
 MUX2_X1 _08489_ (.A(\registers[12][17] ),
    .B(\registers[14][17] ),
    .S(_02156_),
    .Z(_02271_));
 MUX2_X1 _08490_ (.A(\registers[13][17] ),
    .B(\registers[15][17] ),
    .S(_02158_),
    .Z(_02272_));
 MUX2_X1 _08491_ (.A(_02271_),
    .B(_02272_),
    .S(_02160_),
    .Z(_02273_));
 MUX2_X1 _08492_ (.A(\registers[8][17] ),
    .B(\registers[10][17] ),
    .S(_02162_),
    .Z(_02274_));
 MUX2_X1 _08493_ (.A(\registers[9][17] ),
    .B(\registers[11][17] ),
    .S(_02164_),
    .Z(_02275_));
 MUX2_X1 _08494_ (.A(_02274_),
    .B(_02275_),
    .S(_01931_),
    .Z(_02276_));
 MUX2_X1 _08495_ (.A(_02273_),
    .B(_02276_),
    .S(_01936_),
    .Z(_02277_));
 OAI221_X1 _08496_ (.A(_01910_),
    .B1(_01912_),
    .B2(_02270_),
    .C1(_02277_),
    .C2(_01939_),
    .ZN(_02278_));
 OAI22_X1 _08497_ (.A1(_02243_),
    .A2(_01945_),
    .B1(_02261_),
    .B2(_02278_),
    .ZN(_00337_));
 INV_X1 _08498_ (.A(net14),
    .ZN(_02279_));
 MUX2_X1 _08499_ (.A(\registers[0][18] ),
    .B(\registers[1][18] ),
    .S(_02207_),
    .Z(_02280_));
 MUX2_X1 _08500_ (.A(\registers[6][18] ),
    .B(\registers[7][18] ),
    .S(_02123_),
    .Z(_02281_));
 OAI22_X1 _08501_ (.A1(_02121_),
    .A2(_02280_),
    .B1(_02281_),
    .B2(_02125_),
    .ZN(_02282_));
 MUX2_X1 _08502_ (.A(\registers[2][18] ),
    .B(\registers[3][18] ),
    .S(_02052_),
    .Z(_02283_));
 INV_X1 _08503_ (.A(_02283_),
    .ZN(_02284_));
 AOI21_X1 _08504_ (.A(_02282_),
    .B1(_02284_),
    .B2(_01884_),
    .ZN(_02285_));
 MUX2_X1 _08505_ (.A(\registers[4][18] ),
    .B(\registers[5][18] ),
    .S(_02250_),
    .Z(_02286_));
 INV_X1 _08506_ (.A(_02286_),
    .ZN(_02287_));
 AOI21_X1 _08507_ (.A(_02009_),
    .B1(_01891_),
    .B2(_02287_),
    .ZN(_02288_));
 MUX2_X1 _08508_ (.A(\registers[12][18] ),
    .B(\registers[14][18] ),
    .S(_02094_),
    .Z(_02289_));
 MUX2_X1 _08509_ (.A(\registers[13][18] ),
    .B(\registers[15][18] ),
    .S(_02134_),
    .Z(_02290_));
 MUX2_X1 _08510_ (.A(_02289_),
    .B(_02290_),
    .S(_02136_),
    .Z(_02291_));
 MUX2_X1 _08511_ (.A(\registers[8][18] ),
    .B(\registers[10][18] ),
    .S(_02182_),
    .Z(_02292_));
 MUX2_X1 _08512_ (.A(\registers[9][18] ),
    .B(\registers[11][18] ),
    .S(_02221_),
    .Z(_02293_));
 MUX2_X1 _08513_ (.A(_02292_),
    .B(_02293_),
    .S(_02185_),
    .Z(_02294_));
 MUX2_X2 _08514_ (.A(_02291_),
    .B(_02294_),
    .S(_02141_),
    .Z(_02295_));
 AOI221_X2 _08515_ (.A(_01946_),
    .B1(_02285_),
    .B2(_02288_),
    .C1(_02295_),
    .C2(_01906_),
    .ZN(_02296_));
 MUX2_X1 _08516_ (.A(\registers[28][18] ),
    .B(\registers[30][18] ),
    .S(_01975_),
    .Z(_02297_));
 MUX2_X1 _08517_ (.A(\registers[29][18] ),
    .B(\registers[31][18] ),
    .S(_01977_),
    .Z(_02298_));
 BUF_X4 _08518_ (.A(_01869_),
    .Z(_02299_));
 MUX2_X1 _08519_ (.A(_02297_),
    .B(_02298_),
    .S(_02299_),
    .Z(_02300_));
 MUX2_X1 _08520_ (.A(\registers[24][18] ),
    .B(\registers[26][18] ),
    .S(_01981_),
    .Z(_02301_));
 MUX2_X1 _08521_ (.A(\registers[25][18] ),
    .B(\registers[27][18] ),
    .S(_01983_),
    .Z(_02302_));
 MUX2_X1 _08522_ (.A(_02301_),
    .B(_02302_),
    .S(_01914_),
    .Z(_02303_));
 MUX2_X1 _08523_ (.A(_02300_),
    .B(_02303_),
    .S(_01987_),
    .Z(_02304_));
 MUX2_X1 _08524_ (.A(\registers[16][18] ),
    .B(\registers[17][18] ),
    .S(_02030_),
    .Z(_02305_));
 NOR2_X1 _08525_ (.A1(_02028_),
    .A2(_02305_),
    .ZN(_02306_));
 BUF_X4 _08526_ (.A(_01947_),
    .Z(_02307_));
 MUX2_X1 _08527_ (.A(\registers[18][18] ),
    .B(\registers[19][18] ),
    .S(_02307_),
    .Z(_02308_));
 NOR3_X1 _08528_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02308_),
    .ZN(_02309_));
 MUX2_X1 _08529_ (.A(\registers[20][18] ),
    .B(\registers[21][18] ),
    .S(_01925_),
    .Z(_02310_));
 NOR3_X1 _08530_ (.A1(_02038_),
    .A2(_02039_),
    .A3(_02310_),
    .ZN(_02311_));
 BUF_X4 _08531_ (.A(_01947_),
    .Z(_02312_));
 MUX2_X1 _08532_ (.A(\registers[22][18] ),
    .B(\registers[23][18] ),
    .S(_02312_),
    .Z(_02313_));
 NOR2_X1 _08533_ (.A1(_02042_),
    .A2(_02313_),
    .ZN(_02314_));
 NOR4_X2 _08534_ (.A1(_02306_),
    .A2(_02309_),
    .A3(_02311_),
    .A4(_02314_),
    .ZN(_02315_));
 OAI221_X1 _08535_ (.A(_01910_),
    .B1(_01974_),
    .B2(_02304_),
    .C1(_02315_),
    .C2(_01990_),
    .ZN(_02316_));
 OAI22_X1 _08536_ (.A1(_02279_),
    .A2(_01945_),
    .B1(_02296_),
    .B2(_02316_),
    .ZN(_00338_));
 INV_X1 _08537_ (.A(net15),
    .ZN(_02317_));
 MUX2_X1 _08538_ (.A(\registers[0][19] ),
    .B(\registers[1][19] ),
    .S(_02207_),
    .Z(_02318_));
 MUX2_X1 _08539_ (.A(\registers[6][19] ),
    .B(\registers[7][19] ),
    .S(_02123_),
    .Z(_02319_));
 OAI22_X1 _08540_ (.A1(_02121_),
    .A2(_02318_),
    .B1(_02319_),
    .B2(_02125_),
    .ZN(_02320_));
 MUX2_X1 _08541_ (.A(\registers[2][19] ),
    .B(\registers[3][19] ),
    .S(_02052_),
    .Z(_02321_));
 INV_X1 _08542_ (.A(_02321_),
    .ZN(_02322_));
 CLKBUF_X3 _08543_ (.A(_01883_),
    .Z(_02323_));
 AOI21_X1 _08544_ (.A(_02320_),
    .B1(_02322_),
    .B2(_02323_),
    .ZN(_02324_));
 CLKBUF_X3 _08545_ (.A(_01890_),
    .Z(_02325_));
 MUX2_X1 _08546_ (.A(\registers[4][19] ),
    .B(\registers[5][19] ),
    .S(_02250_),
    .Z(_02326_));
 INV_X1 _08547_ (.A(_02326_),
    .ZN(_02327_));
 AOI21_X1 _08548_ (.A(_02009_),
    .B1(_02325_),
    .B2(_02327_),
    .ZN(_02328_));
 MUX2_X1 _08549_ (.A(\registers[12][19] ),
    .B(\registers[14][19] ),
    .S(_02094_),
    .Z(_02329_));
 MUX2_X1 _08550_ (.A(\registers[13][19] ),
    .B(\registers[15][19] ),
    .S(_02134_),
    .Z(_02330_));
 MUX2_X1 _08551_ (.A(_02329_),
    .B(_02330_),
    .S(_02136_),
    .Z(_02331_));
 MUX2_X1 _08552_ (.A(\registers[8][19] ),
    .B(\registers[10][19] ),
    .S(_02182_),
    .Z(_02332_));
 MUX2_X1 _08553_ (.A(\registers[9][19] ),
    .B(\registers[11][19] ),
    .S(_02221_),
    .Z(_02333_));
 MUX2_X1 _08554_ (.A(_02332_),
    .B(_02333_),
    .S(_02185_),
    .Z(_02334_));
 MUX2_X1 _08555_ (.A(_02331_),
    .B(_02334_),
    .S(_02141_),
    .Z(_02335_));
 BUF_X4 _08556_ (.A(_01887_),
    .Z(_02336_));
 AOI221_X1 _08557_ (.A(_01946_),
    .B1(_02324_),
    .B2(_02328_),
    .C1(_02335_),
    .C2(_02336_),
    .ZN(_02337_));
 CLKBUF_X3 _08558_ (.A(_01909_),
    .Z(_02338_));
 MUX2_X1 _08559_ (.A(\registers[28][19] ),
    .B(\registers[30][19] ),
    .S(_01975_),
    .Z(_02339_));
 MUX2_X1 _08560_ (.A(\registers[29][19] ),
    .B(\registers[31][19] ),
    .S(_01977_),
    .Z(_02340_));
 MUX2_X1 _08561_ (.A(_02339_),
    .B(_02340_),
    .S(_02299_),
    .Z(_02341_));
 MUX2_X1 _08562_ (.A(\registers[24][19] ),
    .B(\registers[26][19] ),
    .S(_01981_),
    .Z(_02342_));
 MUX2_X1 _08563_ (.A(\registers[25][19] ),
    .B(\registers[27][19] ),
    .S(_01983_),
    .Z(_02343_));
 BUF_X4 _08564_ (.A(_01869_),
    .Z(_02344_));
 MUX2_X1 _08565_ (.A(_02342_),
    .B(_02343_),
    .S(_02344_),
    .Z(_02345_));
 MUX2_X1 _08566_ (.A(_02341_),
    .B(_02345_),
    .S(_01987_),
    .Z(_02346_));
 MUX2_X1 _08567_ (.A(\registers[16][19] ),
    .B(\registers[17][19] ),
    .S(_02030_),
    .Z(_02347_));
 NOR2_X1 _08568_ (.A1(_02028_),
    .A2(_02347_),
    .ZN(_02348_));
 MUX2_X1 _08569_ (.A(\registers[18][19] ),
    .B(\registers[19][19] ),
    .S(_02307_),
    .Z(_02349_));
 NOR3_X1 _08570_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02349_),
    .ZN(_02350_));
 MUX2_X1 _08571_ (.A(\registers[20][19] ),
    .B(\registers[21][19] ),
    .S(_01925_),
    .Z(_02351_));
 NOR3_X1 _08572_ (.A1(_02038_),
    .A2(_02039_),
    .A3(_02351_),
    .ZN(_02352_));
 MUX2_X1 _08573_ (.A(\registers[22][19] ),
    .B(\registers[23][19] ),
    .S(_02312_),
    .Z(_02353_));
 NOR2_X1 _08574_ (.A1(_02042_),
    .A2(_02353_),
    .ZN(_02354_));
 NOR4_X2 _08575_ (.A1(_02348_),
    .A2(_02350_),
    .A3(_02352_),
    .A4(_02354_),
    .ZN(_02355_));
 OAI221_X1 _08576_ (.A(_02338_),
    .B1(_01974_),
    .B2(_02346_),
    .C1(_02355_),
    .C2(_01990_),
    .ZN(_02356_));
 OAI22_X1 _08577_ (.A1(_02317_),
    .A2(_01945_),
    .B1(_02337_),
    .B2(_02356_),
    .ZN(_00339_));
 INV_X1 _08578_ (.A(net16),
    .ZN(_02357_));
 CLKBUF_X3 _08579_ (.A(_01942_),
    .Z(_02358_));
 MUX2_X1 _08580_ (.A(\registers[0][1] ),
    .B(\registers[1][1] ),
    .S(_02207_),
    .Z(_02359_));
 MUX2_X1 _08581_ (.A(\registers[6][1] ),
    .B(\registers[7][1] ),
    .S(_02123_),
    .Z(_02360_));
 OAI22_X1 _08582_ (.A1(_02121_),
    .A2(_02359_),
    .B1(_02360_),
    .B2(_02125_),
    .ZN(_02361_));
 MUX2_X1 _08583_ (.A(\registers[2][1] ),
    .B(\registers[3][1] ),
    .S(_02052_),
    .Z(_02362_));
 INV_X1 _08584_ (.A(_02362_),
    .ZN(_02363_));
 AOI21_X1 _08585_ (.A(_02361_),
    .B1(_02363_),
    .B2(_02323_),
    .ZN(_02364_));
 MUX2_X1 _08586_ (.A(\registers[4][1] ),
    .B(\registers[5][1] ),
    .S(_02250_),
    .Z(_02365_));
 INV_X1 _08587_ (.A(_02365_),
    .ZN(_02366_));
 AOI21_X1 _08588_ (.A(_02009_),
    .B1(_02325_),
    .B2(_02366_),
    .ZN(_02367_));
 MUX2_X1 _08589_ (.A(\registers[12][1] ),
    .B(\registers[14][1] ),
    .S(_02094_),
    .Z(_02368_));
 MUX2_X1 _08590_ (.A(\registers[13][1] ),
    .B(\registers[15][1] ),
    .S(_02134_),
    .Z(_02369_));
 MUX2_X1 _08591_ (.A(_02368_),
    .B(_02369_),
    .S(_02136_),
    .Z(_02370_));
 MUX2_X1 _08592_ (.A(\registers[8][1] ),
    .B(\registers[10][1] ),
    .S(_02182_),
    .Z(_02371_));
 MUX2_X1 _08593_ (.A(\registers[9][1] ),
    .B(\registers[11][1] ),
    .S(_02221_),
    .Z(_02372_));
 MUX2_X1 _08594_ (.A(_02371_),
    .B(_02372_),
    .S(_02185_),
    .Z(_02373_));
 MUX2_X2 _08595_ (.A(_02370_),
    .B(_02373_),
    .S(_02141_),
    .Z(_02374_));
 AOI221_X2 _08596_ (.A(_01946_),
    .B1(_02364_),
    .B2(_02367_),
    .C1(_02374_),
    .C2(_02336_),
    .ZN(_02375_));
 BUF_X8 _08597_ (.A(_01862_),
    .Z(_02376_));
 MUX2_X1 _08598_ (.A(\registers[28][1] ),
    .B(\registers[30][1] ),
    .S(_02376_),
    .Z(_02377_));
 MUX2_X1 _08599_ (.A(\registers[29][1] ),
    .B(\registers[31][1] ),
    .S(_01977_),
    .Z(_02378_));
 MUX2_X1 _08600_ (.A(_02377_),
    .B(_02378_),
    .S(_02299_),
    .Z(_02379_));
 MUX2_X1 _08601_ (.A(\registers[24][1] ),
    .B(\registers[26][1] ),
    .S(_01981_),
    .Z(_02380_));
 MUX2_X1 _08602_ (.A(\registers[25][1] ),
    .B(\registers[27][1] ),
    .S(_01983_),
    .Z(_02381_));
 MUX2_X1 _08603_ (.A(_02380_),
    .B(_02381_),
    .S(_02344_),
    .Z(_02382_));
 MUX2_X1 _08604_ (.A(_02379_),
    .B(_02382_),
    .S(_01987_),
    .Z(_02383_));
 MUX2_X1 _08605_ (.A(\registers[16][1] ),
    .B(\registers[17][1] ),
    .S(_02030_),
    .Z(_02384_));
 NOR2_X1 _08606_ (.A1(_02028_),
    .A2(_02384_),
    .ZN(_02385_));
 MUX2_X1 _08607_ (.A(\registers[18][1] ),
    .B(\registers[19][1] ),
    .S(_02307_),
    .Z(_02386_));
 NOR3_X1 _08608_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02386_),
    .ZN(_02387_));
 MUX2_X1 _08609_ (.A(\registers[20][1] ),
    .B(\registers[21][1] ),
    .S(_01925_),
    .Z(_02388_));
 NOR3_X1 _08610_ (.A1(_02038_),
    .A2(_02039_),
    .A3(_02388_),
    .ZN(_02389_));
 MUX2_X1 _08611_ (.A(\registers[22][1] ),
    .B(\registers[23][1] ),
    .S(_02312_),
    .Z(_02390_));
 NOR2_X1 _08612_ (.A1(_02042_),
    .A2(_02390_),
    .ZN(_02391_));
 NOR4_X2 _08613_ (.A1(_02385_),
    .A2(_02387_),
    .A3(_02389_),
    .A4(_02391_),
    .ZN(_02392_));
 OAI221_X1 _08614_ (.A(_02338_),
    .B1(_01974_),
    .B2(_02383_),
    .C1(_02392_),
    .C2(_01990_),
    .ZN(_02393_));
 OAI22_X1 _08615_ (.A1(_02357_),
    .A2(_02358_),
    .B1(_02375_),
    .B2(_02393_),
    .ZN(_00340_));
 INV_X1 _08616_ (.A(net17),
    .ZN(_02394_));
 MUX2_X1 _08617_ (.A(\registers[0][20] ),
    .B(\registers[1][20] ),
    .S(_02207_),
    .Z(_02395_));
 MUX2_X1 _08618_ (.A(\registers[6][20] ),
    .B(\registers[7][20] ),
    .S(_02123_),
    .Z(_02396_));
 OAI22_X1 _08619_ (.A1(_02121_),
    .A2(_02395_),
    .B1(_02396_),
    .B2(_02125_),
    .ZN(_02397_));
 MUX2_X1 _08620_ (.A(\registers[2][20] ),
    .B(\registers[3][20] ),
    .S(_02052_),
    .Z(_02398_));
 INV_X1 _08621_ (.A(_02398_),
    .ZN(_02399_));
 AOI21_X1 _08622_ (.A(_02397_),
    .B1(_02399_),
    .B2(_02323_),
    .ZN(_02400_));
 CLKBUF_X3 _08623_ (.A(_01886_),
    .Z(_02401_));
 MUX2_X1 _08624_ (.A(\registers[4][20] ),
    .B(\registers[5][20] ),
    .S(_02250_),
    .Z(_02402_));
 INV_X1 _08625_ (.A(_02402_),
    .ZN(_02403_));
 AOI21_X1 _08626_ (.A(_02401_),
    .B1(_02325_),
    .B2(_02403_),
    .ZN(_02404_));
 MUX2_X1 _08627_ (.A(\registers[12][20] ),
    .B(\registers[14][20] ),
    .S(_02094_),
    .Z(_02405_));
 MUX2_X1 _08628_ (.A(\registers[13][20] ),
    .B(\registers[15][20] ),
    .S(_02134_),
    .Z(_02406_));
 MUX2_X1 _08629_ (.A(_02405_),
    .B(_02406_),
    .S(_02136_),
    .Z(_02407_));
 MUX2_X1 _08630_ (.A(\registers[8][20] ),
    .B(\registers[10][20] ),
    .S(_02182_),
    .Z(_02408_));
 MUX2_X1 _08631_ (.A(\registers[9][20] ),
    .B(\registers[11][20] ),
    .S(_02221_),
    .Z(_02409_));
 MUX2_X1 _08632_ (.A(_02408_),
    .B(_02409_),
    .S(_02185_),
    .Z(_02410_));
 MUX2_X1 _08633_ (.A(_02407_),
    .B(_02410_),
    .S(_02141_),
    .Z(_02411_));
 AOI221_X1 _08634_ (.A(_01946_),
    .B1(_02400_),
    .B2(_02404_),
    .C1(_02411_),
    .C2(_02336_),
    .ZN(_02412_));
 MUX2_X1 _08635_ (.A(\registers[28][20] ),
    .B(\registers[30][20] ),
    .S(_02376_),
    .Z(_02413_));
 BUF_X8 _08636_ (.A(_01862_),
    .Z(_02414_));
 MUX2_X1 _08637_ (.A(\registers[29][20] ),
    .B(\registers[31][20] ),
    .S(_02414_),
    .Z(_02415_));
 MUX2_X1 _08638_ (.A(_02413_),
    .B(_02415_),
    .S(_02299_),
    .Z(_02416_));
 MUX2_X1 _08639_ (.A(\registers[24][20] ),
    .B(\registers[26][20] ),
    .S(_01981_),
    .Z(_02417_));
 MUX2_X1 _08640_ (.A(\registers[25][20] ),
    .B(\registers[27][20] ),
    .S(_01983_),
    .Z(_02418_));
 MUX2_X1 _08641_ (.A(_02417_),
    .B(_02418_),
    .S(_02344_),
    .Z(_02419_));
 MUX2_X1 _08642_ (.A(_02416_),
    .B(_02419_),
    .S(_01987_),
    .Z(_02420_));
 MUX2_X1 _08643_ (.A(\registers[16][20] ),
    .B(\registers[17][20] ),
    .S(_02030_),
    .Z(_02421_));
 NOR2_X1 _08644_ (.A1(_02028_),
    .A2(_02421_),
    .ZN(_02422_));
 MUX2_X1 _08645_ (.A(\registers[18][20] ),
    .B(\registers[19][20] ),
    .S(_02307_),
    .Z(_02423_));
 NOR3_X1 _08646_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02423_),
    .ZN(_02424_));
 MUX2_X1 _08647_ (.A(\registers[20][20] ),
    .B(\registers[21][20] ),
    .S(_01925_),
    .Z(_02425_));
 NOR3_X1 _08648_ (.A1(_02038_),
    .A2(_02039_),
    .A3(_02425_),
    .ZN(_02426_));
 MUX2_X1 _08649_ (.A(\registers[22][20] ),
    .B(\registers[23][20] ),
    .S(_02312_),
    .Z(_02427_));
 NOR2_X1 _08650_ (.A1(_02042_),
    .A2(_02427_),
    .ZN(_02428_));
 NOR4_X2 _08651_ (.A1(_02422_),
    .A2(_02424_),
    .A3(_02426_),
    .A4(_02428_),
    .ZN(_02429_));
 OAI221_X1 _08652_ (.A(_02338_),
    .B1(_01974_),
    .B2(_02420_),
    .C1(_02429_),
    .C2(_01990_),
    .ZN(_02430_));
 OAI22_X1 _08653_ (.A1(_02394_),
    .A2(_02358_),
    .B1(_02412_),
    .B2(_02430_),
    .ZN(_00341_));
 INV_X1 _08654_ (.A(net18),
    .ZN(_02431_));
 MUX2_X1 _08655_ (.A(\registers[0][21] ),
    .B(\registers[1][21] ),
    .S(_02207_),
    .Z(_02432_));
 MUX2_X1 _08656_ (.A(\registers[6][21] ),
    .B(\registers[7][21] ),
    .S(_02123_),
    .Z(_02433_));
 OAI22_X1 _08657_ (.A1(_02121_),
    .A2(_02432_),
    .B1(_02433_),
    .B2(_02125_),
    .ZN(_02434_));
 BUF_X4 _08658_ (.A(_01877_),
    .Z(_02435_));
 MUX2_X1 _08659_ (.A(\registers[2][21] ),
    .B(\registers[3][21] ),
    .S(_02435_),
    .Z(_02436_));
 INV_X1 _08660_ (.A(_02436_),
    .ZN(_02437_));
 AOI21_X1 _08661_ (.A(_02434_),
    .B1(_02437_),
    .B2(_02323_),
    .ZN(_02438_));
 MUX2_X1 _08662_ (.A(\registers[4][21] ),
    .B(\registers[5][21] ),
    .S(_02250_),
    .Z(_02439_));
 INV_X1 _08663_ (.A(_02439_),
    .ZN(_02440_));
 AOI21_X1 _08664_ (.A(_02401_),
    .B1(_02325_),
    .B2(_02440_),
    .ZN(_02441_));
 MUX2_X1 _08665_ (.A(\registers[12][21] ),
    .B(\registers[14][21] ),
    .S(_02094_),
    .Z(_02442_));
 MUX2_X1 _08666_ (.A(\registers[13][21] ),
    .B(\registers[15][21] ),
    .S(_02134_),
    .Z(_02443_));
 MUX2_X1 _08667_ (.A(_02442_),
    .B(_02443_),
    .S(_02136_),
    .Z(_02444_));
 MUX2_X1 _08668_ (.A(\registers[8][21] ),
    .B(\registers[10][21] ),
    .S(_02182_),
    .Z(_02445_));
 MUX2_X1 _08669_ (.A(\registers[9][21] ),
    .B(\registers[11][21] ),
    .S(_02221_),
    .Z(_02446_));
 MUX2_X1 _08670_ (.A(_02445_),
    .B(_02446_),
    .S(_02185_),
    .Z(_02447_));
 MUX2_X2 _08671_ (.A(_02444_),
    .B(_02447_),
    .S(_02141_),
    .Z(_02448_));
 AOI221_X2 _08672_ (.A(_01946_),
    .B1(_02438_),
    .B2(_02441_),
    .C1(_02448_),
    .C2(_02336_),
    .ZN(_02449_));
 MUX2_X1 _08673_ (.A(\registers[28][21] ),
    .B(\registers[30][21] ),
    .S(_02376_),
    .Z(_02450_));
 MUX2_X1 _08674_ (.A(\registers[29][21] ),
    .B(\registers[31][21] ),
    .S(_02414_),
    .Z(_02451_));
 MUX2_X1 _08675_ (.A(_02450_),
    .B(_02451_),
    .S(_02299_),
    .Z(_02452_));
 BUF_X8 _08676_ (.A(_01862_),
    .Z(_02453_));
 MUX2_X1 _08677_ (.A(\registers[24][21] ),
    .B(\registers[26][21] ),
    .S(_02453_),
    .Z(_02454_));
 MUX2_X1 _08678_ (.A(\registers[25][21] ),
    .B(\registers[27][21] ),
    .S(_01983_),
    .Z(_02455_));
 MUX2_X1 _08679_ (.A(_02454_),
    .B(_02455_),
    .S(_02344_),
    .Z(_02456_));
 BUF_X4 _08680_ (.A(_01986_),
    .Z(_02457_));
 MUX2_X1 _08681_ (.A(_02452_),
    .B(_02456_),
    .S(_02457_),
    .Z(_02458_));
 BUF_X4 _08682_ (.A(_01892_),
    .Z(_02459_));
 MUX2_X1 _08683_ (.A(\registers[16][21] ),
    .B(\registers[17][21] ),
    .S(_02459_),
    .Z(_02460_));
 NOR2_X1 _08684_ (.A1(_02028_),
    .A2(_02460_),
    .ZN(_02461_));
 MUX2_X1 _08685_ (.A(\registers[18][21] ),
    .B(\registers[19][21] ),
    .S(_02307_),
    .Z(_02462_));
 NOR3_X1 _08686_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02462_),
    .ZN(_02463_));
 CLKBUF_X3 _08687_ (.A(_01986_),
    .Z(_02464_));
 MUX2_X1 _08688_ (.A(\registers[20][21] ),
    .B(\registers[21][21] ),
    .S(_01925_),
    .Z(_02465_));
 NOR3_X1 _08689_ (.A1(_02038_),
    .A2(_02464_),
    .A3(_02465_),
    .ZN(_02466_));
 MUX2_X1 _08690_ (.A(\registers[22][21] ),
    .B(\registers[23][21] ),
    .S(_02312_),
    .Z(_02467_));
 NOR2_X1 _08691_ (.A1(_02042_),
    .A2(_02467_),
    .ZN(_02468_));
 NOR4_X2 _08692_ (.A1(_02461_),
    .A2(_02463_),
    .A3(_02466_),
    .A4(_02468_),
    .ZN(_02469_));
 OAI221_X1 _08693_ (.A(_02338_),
    .B1(_01974_),
    .B2(_02458_),
    .C1(_02469_),
    .C2(_01990_),
    .ZN(_02470_));
 OAI22_X1 _08694_ (.A1(_02431_),
    .A2(_02358_),
    .B1(_02449_),
    .B2(_02470_),
    .ZN(_00342_));
 INV_X1 _08695_ (.A(net19),
    .ZN(_02471_));
 BUF_X4 _08696_ (.A(_01858_),
    .Z(_02472_));
 MUX2_X1 _08697_ (.A(\registers[0][22] ),
    .B(\registers[1][22] ),
    .S(_02207_),
    .Z(_02473_));
 MUX2_X1 _08698_ (.A(\registers[6][22] ),
    .B(\registers[7][22] ),
    .S(_02123_),
    .Z(_02474_));
 OAI22_X1 _08699_ (.A1(_02121_),
    .A2(_02473_),
    .B1(_02474_),
    .B2(_02125_),
    .ZN(_02475_));
 MUX2_X1 _08700_ (.A(\registers[2][22] ),
    .B(\registers[3][22] ),
    .S(_02435_),
    .Z(_02476_));
 INV_X1 _08701_ (.A(_02476_),
    .ZN(_02477_));
 AOI21_X1 _08702_ (.A(_02475_),
    .B1(_02477_),
    .B2(_02323_),
    .ZN(_02478_));
 MUX2_X1 _08703_ (.A(\registers[4][22] ),
    .B(\registers[5][22] ),
    .S(_02250_),
    .Z(_02479_));
 INV_X1 _08704_ (.A(_02479_),
    .ZN(_02480_));
 AOI21_X1 _08705_ (.A(_02401_),
    .B1(_02325_),
    .B2(_02480_),
    .ZN(_02481_));
 BUF_X4 _08706_ (.A(_01959_),
    .Z(_02482_));
 MUX2_X1 _08707_ (.A(\registers[12][22] ),
    .B(\registers[14][22] ),
    .S(_02482_),
    .Z(_02483_));
 MUX2_X1 _08708_ (.A(\registers[13][22] ),
    .B(\registers[15][22] ),
    .S(_02134_),
    .Z(_02484_));
 MUX2_X1 _08709_ (.A(_02483_),
    .B(_02484_),
    .S(_02136_),
    .Z(_02485_));
 MUX2_X1 _08710_ (.A(\registers[8][22] ),
    .B(\registers[10][22] ),
    .S(_02182_),
    .Z(_02486_));
 MUX2_X1 _08711_ (.A(\registers[9][22] ),
    .B(\registers[11][22] ),
    .S(_02221_),
    .Z(_02487_));
 MUX2_X1 _08712_ (.A(_02486_),
    .B(_02487_),
    .S(_02185_),
    .Z(_02488_));
 MUX2_X1 _08713_ (.A(_02485_),
    .B(_02488_),
    .S(_02141_),
    .Z(_02489_));
 AOI221_X1 _08714_ (.A(_02472_),
    .B1(_02478_),
    .B2(_02481_),
    .C1(_02489_),
    .C2(_02336_),
    .ZN(_02490_));
 CLKBUF_X3 _08715_ (.A(_01973_),
    .Z(_02491_));
 MUX2_X1 _08716_ (.A(\registers[28][22] ),
    .B(\registers[30][22] ),
    .S(_02376_),
    .Z(_02492_));
 MUX2_X1 _08717_ (.A(\registers[29][22] ),
    .B(\registers[31][22] ),
    .S(_02414_),
    .Z(_02493_));
 MUX2_X1 _08718_ (.A(_02492_),
    .B(_02493_),
    .S(_02299_),
    .Z(_02494_));
 MUX2_X1 _08719_ (.A(\registers[24][22] ),
    .B(\registers[26][22] ),
    .S(_02453_),
    .Z(_02495_));
 BUF_X8 _08720_ (.A(_01862_),
    .Z(_02496_));
 MUX2_X1 _08721_ (.A(\registers[25][22] ),
    .B(\registers[27][22] ),
    .S(_02496_),
    .Z(_02497_));
 MUX2_X1 _08722_ (.A(_02495_),
    .B(_02497_),
    .S(_02344_),
    .Z(_02498_));
 MUX2_X1 _08723_ (.A(_02494_),
    .B(_02498_),
    .S(_02457_),
    .Z(_02499_));
 MUX2_X1 _08724_ (.A(\registers[16][22] ),
    .B(\registers[17][22] ),
    .S(_02459_),
    .Z(_02500_));
 NOR2_X1 _08725_ (.A1(_02028_),
    .A2(_02500_),
    .ZN(_02501_));
 MUX2_X1 _08726_ (.A(\registers[18][22] ),
    .B(\registers[19][22] ),
    .S(_02307_),
    .Z(_02502_));
 NOR3_X1 _08727_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02502_),
    .ZN(_02503_));
 BUF_X4 _08728_ (.A(_01898_),
    .Z(_02504_));
 MUX2_X1 _08729_ (.A(\registers[20][22] ),
    .B(\registers[21][22] ),
    .S(_02504_),
    .Z(_02505_));
 NOR3_X1 _08730_ (.A1(_02038_),
    .A2(_02464_),
    .A3(_02505_),
    .ZN(_02506_));
 MUX2_X1 _08731_ (.A(\registers[22][22] ),
    .B(\registers[23][22] ),
    .S(_02312_),
    .Z(_02507_));
 NOR2_X1 _08732_ (.A1(_02042_),
    .A2(_02507_),
    .ZN(_02508_));
 NOR4_X2 _08733_ (.A1(_02501_),
    .A2(_02503_),
    .A3(_02506_),
    .A4(_02508_),
    .ZN(_02509_));
 CLKBUF_X3 _08734_ (.A(_01989_),
    .Z(_02510_));
 OAI221_X1 _08735_ (.A(_02338_),
    .B1(_02491_),
    .B2(_02499_),
    .C1(_02509_),
    .C2(_02510_),
    .ZN(_02511_));
 OAI22_X1 _08736_ (.A1(_02471_),
    .A2(_02358_),
    .B1(_02490_),
    .B2(_02511_),
    .ZN(_00343_));
 INV_X1 _08737_ (.A(net20),
    .ZN(_02512_));
 BUF_X4 _08738_ (.A(_01865_),
    .Z(_02513_));
 MUX2_X1 _08739_ (.A(\registers[0][23] ),
    .B(\registers[1][23] ),
    .S(_02207_),
    .Z(_02514_));
 BUF_X4 _08740_ (.A(_01867_),
    .Z(_02515_));
 MUX2_X1 _08741_ (.A(\registers[6][23] ),
    .B(\registers[7][23] ),
    .S(_02515_),
    .Z(_02516_));
 BUF_X4 _08742_ (.A(_01872_),
    .Z(_02517_));
 OAI22_X1 _08743_ (.A1(_02513_),
    .A2(_02514_),
    .B1(_02516_),
    .B2(_02517_),
    .ZN(_02518_));
 MUX2_X1 _08744_ (.A(\registers[2][23] ),
    .B(\registers[3][23] ),
    .S(_02435_),
    .Z(_02519_));
 INV_X1 _08745_ (.A(_02519_),
    .ZN(_02520_));
 AOI21_X1 _08746_ (.A(_02518_),
    .B1(_02520_),
    .B2(_02323_),
    .ZN(_02521_));
 MUX2_X1 _08747_ (.A(\registers[4][23] ),
    .B(\registers[5][23] ),
    .S(_02250_),
    .Z(_02522_));
 INV_X1 _08748_ (.A(_02522_),
    .ZN(_02523_));
 AOI21_X1 _08749_ (.A(_02401_),
    .B1(_02325_),
    .B2(_02523_),
    .ZN(_02524_));
 MUX2_X1 _08750_ (.A(\registers[12][23] ),
    .B(\registers[14][23] ),
    .S(_02482_),
    .Z(_02525_));
 BUF_X4 _08751_ (.A(_01959_),
    .Z(_02526_));
 MUX2_X1 _08752_ (.A(\registers[13][23] ),
    .B(\registers[15][23] ),
    .S(_02526_),
    .Z(_02527_));
 BUF_X4 _08753_ (.A(_01877_),
    .Z(_02528_));
 MUX2_X1 _08754_ (.A(_02525_),
    .B(_02527_),
    .S(_02528_),
    .Z(_02529_));
 MUX2_X1 _08755_ (.A(\registers[8][23] ),
    .B(\registers[10][23] ),
    .S(_02182_),
    .Z(_02530_));
 MUX2_X1 _08756_ (.A(\registers[9][23] ),
    .B(\registers[11][23] ),
    .S(_02221_),
    .Z(_02531_));
 MUX2_X1 _08757_ (.A(_02530_),
    .B(_02531_),
    .S(_02185_),
    .Z(_02532_));
 BUF_X4 _08758_ (.A(_01889_),
    .Z(_02533_));
 MUX2_X1 _08759_ (.A(_02529_),
    .B(_02532_),
    .S(_02533_),
    .Z(_02534_));
 AOI221_X1 _08760_ (.A(_02472_),
    .B1(_02521_),
    .B2(_02524_),
    .C1(_02534_),
    .C2(_02336_),
    .ZN(_02535_));
 MUX2_X1 _08761_ (.A(\registers[28][23] ),
    .B(\registers[30][23] ),
    .S(_02376_),
    .Z(_02536_));
 MUX2_X1 _08762_ (.A(\registers[29][23] ),
    .B(\registers[31][23] ),
    .S(_02414_),
    .Z(_02537_));
 MUX2_X1 _08763_ (.A(_02536_),
    .B(_02537_),
    .S(_02299_),
    .Z(_02538_));
 MUX2_X1 _08764_ (.A(\registers[24][23] ),
    .B(\registers[26][23] ),
    .S(_02453_),
    .Z(_02539_));
 MUX2_X1 _08765_ (.A(\registers[25][23] ),
    .B(\registers[27][23] ),
    .S(_02496_),
    .Z(_02540_));
 MUX2_X1 _08766_ (.A(_02539_),
    .B(_02540_),
    .S(_02344_),
    .Z(_02541_));
 MUX2_X1 _08767_ (.A(_02538_),
    .B(_02541_),
    .S(_02457_),
    .Z(_02542_));
 BUF_X4 _08768_ (.A(_01866_),
    .Z(_02543_));
 MUX2_X1 _08769_ (.A(\registers[16][23] ),
    .B(\registers[17][23] ),
    .S(_02459_),
    .Z(_02544_));
 NOR2_X1 _08770_ (.A1(_02543_),
    .A2(_02544_),
    .ZN(_02545_));
 CLKBUF_X3 _08771_ (.A(_01882_),
    .Z(_02546_));
 CLKBUF_X3 _08772_ (.A(_01863_),
    .Z(_02547_));
 MUX2_X1 _08773_ (.A(\registers[18][23] ),
    .B(\registers[19][23] ),
    .S(_02307_),
    .Z(_02548_));
 NOR3_X1 _08774_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_02548_),
    .ZN(_02549_));
 CLKBUF_X3 _08775_ (.A(_01888_),
    .Z(_02550_));
 MUX2_X1 _08776_ (.A(\registers[20][23] ),
    .B(\registers[21][23] ),
    .S(_02504_),
    .Z(_02551_));
 NOR3_X1 _08777_ (.A1(_02550_),
    .A2(_02464_),
    .A3(_02551_),
    .ZN(_02552_));
 BUF_X4 _08778_ (.A(_01873_),
    .Z(_02553_));
 MUX2_X1 _08779_ (.A(\registers[22][23] ),
    .B(\registers[23][23] ),
    .S(_02312_),
    .Z(_02554_));
 NOR2_X1 _08780_ (.A1(_02553_),
    .A2(_02554_),
    .ZN(_02555_));
 NOR4_X2 _08781_ (.A1(_02545_),
    .A2(_02549_),
    .A3(_02552_),
    .A4(_02555_),
    .ZN(_02556_));
 OAI221_X1 _08782_ (.A(_02338_),
    .B1(_02491_),
    .B2(_02542_),
    .C1(_02556_),
    .C2(_02510_),
    .ZN(_02557_));
 OAI22_X1 _08783_ (.A1(_02512_),
    .A2(_02358_),
    .B1(_02535_),
    .B2(_02557_),
    .ZN(_00344_));
 INV_X1 _08784_ (.A(net21),
    .ZN(_02558_));
 MUX2_X1 _08785_ (.A(\registers[0][24] ),
    .B(\registers[1][24] ),
    .S(_02207_),
    .Z(_02559_));
 MUX2_X1 _08786_ (.A(\registers[6][24] ),
    .B(\registers[7][24] ),
    .S(_02515_),
    .Z(_02560_));
 OAI22_X1 _08787_ (.A1(_02513_),
    .A2(_02559_),
    .B1(_02560_),
    .B2(_02517_),
    .ZN(_02561_));
 MUX2_X1 _08788_ (.A(\registers[2][24] ),
    .B(\registers[3][24] ),
    .S(_02435_),
    .Z(_02562_));
 INV_X1 _08789_ (.A(_02562_),
    .ZN(_02563_));
 AOI21_X1 _08790_ (.A(_02561_),
    .B1(_02563_),
    .B2(_02323_),
    .ZN(_02564_));
 MUX2_X1 _08791_ (.A(\registers[4][24] ),
    .B(\registers[5][24] ),
    .S(_02250_),
    .Z(_02565_));
 INV_X1 _08792_ (.A(_02565_),
    .ZN(_02566_));
 AOI21_X1 _08793_ (.A(_02401_),
    .B1(_02325_),
    .B2(_02566_),
    .ZN(_02567_));
 MUX2_X1 _08794_ (.A(\registers[12][24] ),
    .B(\registers[14][24] ),
    .S(_02482_),
    .Z(_02568_));
 MUX2_X1 _08795_ (.A(\registers[13][24] ),
    .B(\registers[15][24] ),
    .S(_02526_),
    .Z(_02569_));
 MUX2_X1 _08796_ (.A(_02568_),
    .B(_02569_),
    .S(_02528_),
    .Z(_02570_));
 BUF_X4 _08797_ (.A(_01959_),
    .Z(_02571_));
 MUX2_X1 _08798_ (.A(\registers[8][24] ),
    .B(\registers[10][24] ),
    .S(_02571_),
    .Z(_02572_));
 MUX2_X1 _08799_ (.A(\registers[9][24] ),
    .B(\registers[11][24] ),
    .S(_02221_),
    .Z(_02573_));
 BUF_X4 _08800_ (.A(_01877_),
    .Z(_02574_));
 MUX2_X1 _08801_ (.A(_02572_),
    .B(_02573_),
    .S(_02574_),
    .Z(_02575_));
 MUX2_X2 _08802_ (.A(_02570_),
    .B(_02575_),
    .S(_02533_),
    .Z(_02576_));
 AOI221_X1 _08803_ (.A(_02472_),
    .B1(_02564_),
    .B2(_02567_),
    .C1(_02576_),
    .C2(_02336_),
    .ZN(_02577_));
 MUX2_X1 _08804_ (.A(\registers[28][24] ),
    .B(\registers[30][24] ),
    .S(_02376_),
    .Z(_02578_));
 MUX2_X1 _08805_ (.A(\registers[29][24] ),
    .B(\registers[31][24] ),
    .S(_02414_),
    .Z(_02579_));
 MUX2_X1 _08806_ (.A(_02578_),
    .B(_02579_),
    .S(_02299_),
    .Z(_02580_));
 MUX2_X1 _08807_ (.A(\registers[24][24] ),
    .B(\registers[26][24] ),
    .S(_02453_),
    .Z(_02581_));
 MUX2_X1 _08808_ (.A(\registers[25][24] ),
    .B(\registers[27][24] ),
    .S(_02496_),
    .Z(_02582_));
 MUX2_X1 _08809_ (.A(_02581_),
    .B(_02582_),
    .S(_02344_),
    .Z(_02583_));
 MUX2_X1 _08810_ (.A(_02580_),
    .B(_02583_),
    .S(_02457_),
    .Z(_02584_));
 MUX2_X1 _08811_ (.A(\registers[16][24] ),
    .B(\registers[17][24] ),
    .S(_02459_),
    .Z(_02585_));
 NOR2_X1 _08812_ (.A1(_02543_),
    .A2(_02585_),
    .ZN(_02586_));
 MUX2_X1 _08813_ (.A(\registers[18][24] ),
    .B(\registers[19][24] ),
    .S(_02307_),
    .Z(_02587_));
 NOR3_X1 _08814_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_02587_),
    .ZN(_02588_));
 MUX2_X1 _08815_ (.A(\registers[20][24] ),
    .B(\registers[21][24] ),
    .S(_02504_),
    .Z(_02589_));
 NOR3_X1 _08816_ (.A1(_02550_),
    .A2(_02464_),
    .A3(_02589_),
    .ZN(_02590_));
 MUX2_X1 _08817_ (.A(\registers[22][24] ),
    .B(\registers[23][24] ),
    .S(_02312_),
    .Z(_02591_));
 NOR2_X1 _08818_ (.A1(_02553_),
    .A2(_02591_),
    .ZN(_02592_));
 NOR4_X2 _08819_ (.A1(_02586_),
    .A2(_02588_),
    .A3(_02590_),
    .A4(_02592_),
    .ZN(_02593_));
 OAI221_X1 _08820_ (.A(_02338_),
    .B1(_02491_),
    .B2(_02584_),
    .C1(_02593_),
    .C2(_02510_),
    .ZN(_02594_));
 OAI22_X1 _08821_ (.A1(_02558_),
    .A2(_02358_),
    .B1(_02577_),
    .B2(_02594_),
    .ZN(_00345_));
 INV_X1 _08822_ (.A(net22),
    .ZN(_02595_));
 BUF_X4 _08823_ (.A(_01868_),
    .Z(_02596_));
 MUX2_X1 _08824_ (.A(\registers[0][25] ),
    .B(\registers[1][25] ),
    .S(_02596_),
    .Z(_02597_));
 MUX2_X1 _08825_ (.A(\registers[6][25] ),
    .B(\registers[7][25] ),
    .S(_02515_),
    .Z(_02598_));
 OAI22_X1 _08826_ (.A1(_02513_),
    .A2(_02597_),
    .B1(_02598_),
    .B2(_02517_),
    .ZN(_02599_));
 MUX2_X1 _08827_ (.A(\registers[2][25] ),
    .B(\registers[3][25] ),
    .S(_02435_),
    .Z(_02600_));
 INV_X1 _08828_ (.A(_02600_),
    .ZN(_02601_));
 AOI21_X1 _08829_ (.A(_02599_),
    .B1(_02601_),
    .B2(_02323_),
    .ZN(_02602_));
 MUX2_X1 _08830_ (.A(\registers[4][25] ),
    .B(\registers[5][25] ),
    .S(_02250_),
    .Z(_02603_));
 INV_X1 _08831_ (.A(_02603_),
    .ZN(_02604_));
 AOI21_X1 _08832_ (.A(_02401_),
    .B1(_02325_),
    .B2(_02604_),
    .ZN(_02605_));
 MUX2_X1 _08833_ (.A(\registers[12][25] ),
    .B(\registers[14][25] ),
    .S(_02482_),
    .Z(_02606_));
 MUX2_X1 _08834_ (.A(\registers[13][25] ),
    .B(\registers[15][25] ),
    .S(_02526_),
    .Z(_02607_));
 MUX2_X1 _08835_ (.A(_02606_),
    .B(_02607_),
    .S(_02528_),
    .Z(_02608_));
 MUX2_X1 _08836_ (.A(\registers[8][25] ),
    .B(\registers[10][25] ),
    .S(_02571_),
    .Z(_02609_));
 BUF_X4 _08837_ (.A(_01959_),
    .Z(_02610_));
 MUX2_X1 _08838_ (.A(\registers[9][25] ),
    .B(\registers[11][25] ),
    .S(_02610_),
    .Z(_02611_));
 MUX2_X1 _08839_ (.A(_02609_),
    .B(_02611_),
    .S(_02574_),
    .Z(_02612_));
 MUX2_X1 _08840_ (.A(_02608_),
    .B(_02612_),
    .S(_02533_),
    .Z(_02613_));
 AOI221_X1 _08841_ (.A(_02472_),
    .B1(_02602_),
    .B2(_02605_),
    .C1(_02613_),
    .C2(_02336_),
    .ZN(_02614_));
 MUX2_X1 _08842_ (.A(\registers[28][25] ),
    .B(\registers[30][25] ),
    .S(_02376_),
    .Z(_02615_));
 MUX2_X1 _08843_ (.A(\registers[29][25] ),
    .B(\registers[31][25] ),
    .S(_02414_),
    .Z(_02616_));
 MUX2_X1 _08844_ (.A(_02615_),
    .B(_02616_),
    .S(_02299_),
    .Z(_02617_));
 MUX2_X1 _08845_ (.A(\registers[24][25] ),
    .B(\registers[26][25] ),
    .S(_02453_),
    .Z(_02618_));
 MUX2_X1 _08846_ (.A(\registers[25][25] ),
    .B(\registers[27][25] ),
    .S(_02496_),
    .Z(_02619_));
 MUX2_X1 _08847_ (.A(_02618_),
    .B(_02619_),
    .S(_02344_),
    .Z(_02620_));
 MUX2_X1 _08848_ (.A(_02617_),
    .B(_02620_),
    .S(_02457_),
    .Z(_02621_));
 MUX2_X1 _08849_ (.A(\registers[16][25] ),
    .B(\registers[17][25] ),
    .S(_02459_),
    .Z(_02622_));
 NOR2_X1 _08850_ (.A1(_02543_),
    .A2(_02622_),
    .ZN(_02623_));
 MUX2_X1 _08851_ (.A(\registers[18][25] ),
    .B(\registers[19][25] ),
    .S(_02307_),
    .Z(_02624_));
 NOR3_X1 _08852_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_02624_),
    .ZN(_02625_));
 MUX2_X1 _08853_ (.A(\registers[20][25] ),
    .B(\registers[21][25] ),
    .S(_02504_),
    .Z(_02626_));
 NOR3_X1 _08854_ (.A1(_02550_),
    .A2(_02464_),
    .A3(_02626_),
    .ZN(_02627_));
 MUX2_X1 _08855_ (.A(\registers[22][25] ),
    .B(\registers[23][25] ),
    .S(_02312_),
    .Z(_02628_));
 NOR2_X1 _08856_ (.A1(_02553_),
    .A2(_02628_),
    .ZN(_02629_));
 NOR4_X2 _08857_ (.A1(_02623_),
    .A2(_02625_),
    .A3(_02627_),
    .A4(_02629_),
    .ZN(_02630_));
 OAI221_X1 _08858_ (.A(_02338_),
    .B1(_02491_),
    .B2(_02621_),
    .C1(_02630_),
    .C2(_02510_),
    .ZN(_02631_));
 OAI22_X1 _08859_ (.A1(_02595_),
    .A2(_02358_),
    .B1(_02614_),
    .B2(_02631_),
    .ZN(_00346_));
 INV_X1 _08860_ (.A(net23),
    .ZN(_02632_));
 MUX2_X1 _08861_ (.A(\registers[16][26] ),
    .B(\registers[17][26] ),
    .S(_02596_),
    .Z(_02633_));
 MUX2_X1 _08862_ (.A(\registers[22][26] ),
    .B(\registers[23][26] ),
    .S(_02515_),
    .Z(_02634_));
 OAI22_X2 _08863_ (.A1(_02513_),
    .A2(_02633_),
    .B1(_02634_),
    .B2(_02517_),
    .ZN(_02635_));
 MUX2_X1 _08864_ (.A(\registers[18][26] ),
    .B(\registers[19][26] ),
    .S(_02435_),
    .Z(_02636_));
 INV_X1 _08865_ (.A(_02636_),
    .ZN(_02637_));
 AOI21_X1 _08866_ (.A(_02635_),
    .B1(_02637_),
    .B2(_02323_),
    .ZN(_02638_));
 BUF_X4 _08867_ (.A(_01868_),
    .Z(_02639_));
 MUX2_X1 _08868_ (.A(\registers[20][26] ),
    .B(\registers[21][26] ),
    .S(_02639_),
    .Z(_02640_));
 INV_X1 _08869_ (.A(_02640_),
    .ZN(_02641_));
 AOI21_X1 _08870_ (.A(_02401_),
    .B1(_02325_),
    .B2(_02641_),
    .ZN(_02642_));
 MUX2_X1 _08871_ (.A(\registers[28][26] ),
    .B(\registers[30][26] ),
    .S(_02482_),
    .Z(_02643_));
 MUX2_X1 _08872_ (.A(\registers[29][26] ),
    .B(\registers[31][26] ),
    .S(_02526_),
    .Z(_02644_));
 MUX2_X1 _08873_ (.A(_02643_),
    .B(_02644_),
    .S(_02528_),
    .Z(_02645_));
 MUX2_X1 _08874_ (.A(\registers[24][26] ),
    .B(\registers[26][26] ),
    .S(_02571_),
    .Z(_02646_));
 MUX2_X1 _08875_ (.A(\registers[25][26] ),
    .B(\registers[27][26] ),
    .S(_02610_),
    .Z(_02647_));
 MUX2_X1 _08876_ (.A(_02646_),
    .B(_02647_),
    .S(_02574_),
    .Z(_02648_));
 MUX2_X1 _08877_ (.A(_02645_),
    .B(_02648_),
    .S(_02533_),
    .Z(_02649_));
 AOI221_X1 _08878_ (.A(_01860_),
    .B1(_02638_),
    .B2(_02642_),
    .C1(_02649_),
    .C2(_02336_),
    .ZN(_02650_));
 MUX2_X1 _08879_ (.A(\registers[0][26] ),
    .B(\registers[1][26] ),
    .S(_02144_),
    .Z(_02651_));
 NOR2_X1 _08880_ (.A1(_01913_),
    .A2(_02651_),
    .ZN(_02652_));
 MUX2_X1 _08881_ (.A(\registers[2][26] ),
    .B(\registers[3][26] ),
    .S(_01892_),
    .Z(_02653_));
 NOR3_X1 _08882_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_02653_),
    .ZN(_02654_));
 MUX2_X1 _08883_ (.A(\registers[4][26] ),
    .B(\registers[5][26] ),
    .S(_02150_),
    .Z(_02655_));
 NOR3_X1 _08884_ (.A1(_01921_),
    .A2(_01986_),
    .A3(_02655_),
    .ZN(_02656_));
 MUX2_X1 _08885_ (.A(\registers[6][26] ),
    .B(\registers[7][26] ),
    .S(_01951_),
    .Z(_02657_));
 NOR2_X1 _08886_ (.A1(_01924_),
    .A2(_02657_),
    .ZN(_02658_));
 NOR4_X1 _08887_ (.A1(_02652_),
    .A2(_02654_),
    .A3(_02656_),
    .A4(_02658_),
    .ZN(_02659_));
 MUX2_X1 _08888_ (.A(\registers[12][26] ),
    .B(\registers[14][26] ),
    .S(_02156_),
    .Z(_02660_));
 MUX2_X1 _08889_ (.A(\registers[13][26] ),
    .B(\registers[15][26] ),
    .S(_02158_),
    .Z(_02661_));
 MUX2_X1 _08890_ (.A(_02660_),
    .B(_02661_),
    .S(_02160_),
    .Z(_02662_));
 MUX2_X1 _08891_ (.A(\registers[8][26] ),
    .B(\registers[10][26] ),
    .S(_02162_),
    .Z(_02663_));
 MUX2_X1 _08892_ (.A(\registers[9][26] ),
    .B(\registers[11][26] ),
    .S(_02164_),
    .Z(_02664_));
 MUX2_X1 _08893_ (.A(_02663_),
    .B(_02664_),
    .S(_01931_),
    .Z(_02665_));
 MUX2_X1 _08894_ (.A(_02662_),
    .B(_02665_),
    .S(_01936_),
    .Z(_02666_));
 OAI221_X1 _08895_ (.A(_02338_),
    .B1(_01912_),
    .B2(_02659_),
    .C1(_02666_),
    .C2(_01939_),
    .ZN(_02667_));
 OAI22_X1 _08896_ (.A1(_02632_),
    .A2(_02358_),
    .B1(_02650_),
    .B2(_02667_),
    .ZN(_00347_));
 INV_X1 _08897_ (.A(net24),
    .ZN(_02668_));
 MUX2_X1 _08898_ (.A(\registers[0][27] ),
    .B(\registers[1][27] ),
    .S(_02596_),
    .Z(_02669_));
 MUX2_X1 _08899_ (.A(\registers[6][27] ),
    .B(\registers[7][27] ),
    .S(_02515_),
    .Z(_02670_));
 OAI22_X1 _08900_ (.A1(_02513_),
    .A2(_02669_),
    .B1(_02670_),
    .B2(_02517_),
    .ZN(_02671_));
 MUX2_X1 _08901_ (.A(\registers[2][27] ),
    .B(\registers[3][27] ),
    .S(_02435_),
    .Z(_02672_));
 INV_X1 _08902_ (.A(_02672_),
    .ZN(_02673_));
 AOI21_X1 _08903_ (.A(_02671_),
    .B1(_02673_),
    .B2(_02323_),
    .ZN(_02674_));
 MUX2_X1 _08904_ (.A(\registers[4][27] ),
    .B(\registers[5][27] ),
    .S(_02639_),
    .Z(_02675_));
 INV_X1 _08905_ (.A(_02675_),
    .ZN(_02676_));
 AOI21_X1 _08906_ (.A(_02401_),
    .B1(_02325_),
    .B2(_02676_),
    .ZN(_02677_));
 MUX2_X1 _08907_ (.A(\registers[12][27] ),
    .B(\registers[14][27] ),
    .S(_02482_),
    .Z(_02678_));
 MUX2_X1 _08908_ (.A(\registers[13][27] ),
    .B(\registers[15][27] ),
    .S(_02526_),
    .Z(_02679_));
 MUX2_X1 _08909_ (.A(_02678_),
    .B(_02679_),
    .S(_02528_),
    .Z(_02680_));
 MUX2_X1 _08910_ (.A(\registers[8][27] ),
    .B(\registers[10][27] ),
    .S(_02571_),
    .Z(_02681_));
 MUX2_X1 _08911_ (.A(\registers[9][27] ),
    .B(\registers[11][27] ),
    .S(_02610_),
    .Z(_02682_));
 MUX2_X1 _08912_ (.A(_02681_),
    .B(_02682_),
    .S(_02574_),
    .Z(_02683_));
 MUX2_X2 _08913_ (.A(_02680_),
    .B(_02683_),
    .S(_02533_),
    .Z(_02684_));
 AOI221_X2 _08914_ (.A(_02472_),
    .B1(_02674_),
    .B2(_02677_),
    .C1(_02684_),
    .C2(_02336_),
    .ZN(_02685_));
 MUX2_X1 _08915_ (.A(\registers[28][27] ),
    .B(\registers[30][27] ),
    .S(_02376_),
    .Z(_02686_));
 MUX2_X1 _08916_ (.A(\registers[29][27] ),
    .B(\registers[31][27] ),
    .S(_02414_),
    .Z(_02687_));
 MUX2_X1 _08917_ (.A(_02686_),
    .B(_02687_),
    .S(_02299_),
    .Z(_02688_));
 MUX2_X1 _08918_ (.A(\registers[24][27] ),
    .B(\registers[26][27] ),
    .S(_02453_),
    .Z(_02689_));
 MUX2_X1 _08919_ (.A(\registers[25][27] ),
    .B(\registers[27][27] ),
    .S(_02496_),
    .Z(_02690_));
 MUX2_X1 _08920_ (.A(_02689_),
    .B(_02690_),
    .S(_02344_),
    .Z(_02691_));
 MUX2_X1 _08921_ (.A(_02688_),
    .B(_02691_),
    .S(_02457_),
    .Z(_02692_));
 MUX2_X1 _08922_ (.A(\registers[16][27] ),
    .B(\registers[17][27] ),
    .S(_02459_),
    .Z(_02693_));
 NOR2_X1 _08923_ (.A1(_02543_),
    .A2(_02693_),
    .ZN(_02694_));
 MUX2_X1 _08924_ (.A(\registers[18][27] ),
    .B(\registers[19][27] ),
    .S(_02307_),
    .Z(_02695_));
 NOR3_X1 _08925_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_02695_),
    .ZN(_02696_));
 MUX2_X1 _08926_ (.A(\registers[20][27] ),
    .B(\registers[21][27] ),
    .S(_02504_),
    .Z(_02697_));
 NOR3_X1 _08927_ (.A1(_02550_),
    .A2(_02464_),
    .A3(_02697_),
    .ZN(_02698_));
 MUX2_X1 _08928_ (.A(\registers[22][27] ),
    .B(\registers[23][27] ),
    .S(_02312_),
    .Z(_02699_));
 NOR2_X1 _08929_ (.A1(_02553_),
    .A2(_02699_),
    .ZN(_02700_));
 NOR4_X2 _08930_ (.A1(_02694_),
    .A2(_02696_),
    .A3(_02698_),
    .A4(_02700_),
    .ZN(_02701_));
 OAI221_X1 _08931_ (.A(_02338_),
    .B1(_02491_),
    .B2(_02692_),
    .C1(_02701_),
    .C2(_02510_),
    .ZN(_02702_));
 OAI22_X1 _08932_ (.A1(_02668_),
    .A2(_02358_),
    .B1(_02685_),
    .B2(_02702_),
    .ZN(_00348_));
 INV_X1 _08933_ (.A(net25),
    .ZN(_02703_));
 MUX2_X1 _08934_ (.A(\registers[0][28] ),
    .B(\registers[1][28] ),
    .S(_02596_),
    .Z(_02704_));
 MUX2_X1 _08935_ (.A(\registers[6][28] ),
    .B(\registers[7][28] ),
    .S(_02515_),
    .Z(_02705_));
 OAI22_X1 _08936_ (.A1(_02513_),
    .A2(_02704_),
    .B1(_02705_),
    .B2(_02517_),
    .ZN(_02706_));
 MUX2_X1 _08937_ (.A(\registers[2][28] ),
    .B(\registers[3][28] ),
    .S(_02435_),
    .Z(_02707_));
 INV_X1 _08938_ (.A(_02707_),
    .ZN(_02708_));
 BUF_X4 _08939_ (.A(_01883_),
    .Z(_02709_));
 AOI21_X1 _08940_ (.A(_02706_),
    .B1(_02708_),
    .B2(_02709_),
    .ZN(_02710_));
 CLKBUF_X3 _08941_ (.A(_01890_),
    .Z(_02711_));
 MUX2_X1 _08942_ (.A(\registers[4][28] ),
    .B(\registers[5][28] ),
    .S(_02639_),
    .Z(_02712_));
 INV_X1 _08943_ (.A(_02712_),
    .ZN(_02713_));
 AOI21_X1 _08944_ (.A(_02401_),
    .B1(_02711_),
    .B2(_02713_),
    .ZN(_02714_));
 MUX2_X1 _08945_ (.A(\registers[12][28] ),
    .B(\registers[14][28] ),
    .S(_02482_),
    .Z(_02715_));
 MUX2_X1 _08946_ (.A(\registers[13][28] ),
    .B(\registers[15][28] ),
    .S(_02526_),
    .Z(_02716_));
 MUX2_X1 _08947_ (.A(_02715_),
    .B(_02716_),
    .S(_02528_),
    .Z(_02717_));
 MUX2_X1 _08948_ (.A(\registers[8][28] ),
    .B(\registers[10][28] ),
    .S(_02571_),
    .Z(_02718_));
 MUX2_X1 _08949_ (.A(\registers[9][28] ),
    .B(\registers[11][28] ),
    .S(_02610_),
    .Z(_02719_));
 MUX2_X1 _08950_ (.A(_02718_),
    .B(_02719_),
    .S(_02574_),
    .Z(_02720_));
 MUX2_X1 _08951_ (.A(_02717_),
    .B(_02720_),
    .S(_02533_),
    .Z(_02721_));
 BUF_X4 _08952_ (.A(_01887_),
    .Z(_02722_));
 AOI221_X1 _08953_ (.A(_02472_),
    .B1(_02710_),
    .B2(_02714_),
    .C1(_02721_),
    .C2(_02722_),
    .ZN(_02723_));
 CLKBUF_X3 _08954_ (.A(_01909_),
    .Z(_02724_));
 MUX2_X1 _08955_ (.A(\registers[28][28] ),
    .B(\registers[30][28] ),
    .S(_02376_),
    .Z(_02725_));
 MUX2_X1 _08956_ (.A(\registers[29][28] ),
    .B(\registers[31][28] ),
    .S(_02414_),
    .Z(_02726_));
 MUX2_X1 _08957_ (.A(_02725_),
    .B(_02726_),
    .S(_02144_),
    .Z(_02727_));
 MUX2_X1 _08958_ (.A(\registers[24][28] ),
    .B(\registers[26][28] ),
    .S(_02453_),
    .Z(_02728_));
 MUX2_X1 _08959_ (.A(\registers[25][28] ),
    .B(\registers[27][28] ),
    .S(_02496_),
    .Z(_02729_));
 MUX2_X1 _08960_ (.A(_02728_),
    .B(_02729_),
    .S(_02344_),
    .Z(_02730_));
 MUX2_X1 _08961_ (.A(_02727_),
    .B(_02730_),
    .S(_02457_),
    .Z(_02731_));
 MUX2_X1 _08962_ (.A(\registers[16][28] ),
    .B(\registers[17][28] ),
    .S(_02459_),
    .Z(_02732_));
 NOR2_X1 _08963_ (.A1(_02543_),
    .A2(_02732_),
    .ZN(_02733_));
 MUX2_X1 _08964_ (.A(\registers[18][28] ),
    .B(\registers[19][28] ),
    .S(_01899_),
    .Z(_02734_));
 NOR3_X1 _08965_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_02734_),
    .ZN(_02735_));
 MUX2_X1 _08966_ (.A(\registers[20][28] ),
    .B(\registers[21][28] ),
    .S(_02504_),
    .Z(_02736_));
 NOR3_X1 _08967_ (.A1(_02550_),
    .A2(_02464_),
    .A3(_02736_),
    .ZN(_02737_));
 MUX2_X1 _08968_ (.A(\registers[22][28] ),
    .B(\registers[23][28] ),
    .S(_02035_),
    .Z(_02738_));
 NOR2_X1 _08969_ (.A1(_02553_),
    .A2(_02738_),
    .ZN(_02739_));
 NOR4_X2 _08970_ (.A1(_02733_),
    .A2(_02735_),
    .A3(_02737_),
    .A4(_02739_),
    .ZN(_02740_));
 OAI221_X1 _08971_ (.A(_02724_),
    .B1(_02491_),
    .B2(_02731_),
    .C1(_02740_),
    .C2(_02510_),
    .ZN(_02741_));
 OAI22_X1 _08972_ (.A1(_02703_),
    .A2(_02358_),
    .B1(_02723_),
    .B2(_02741_),
    .ZN(_00349_));
 INV_X1 _08973_ (.A(net26),
    .ZN(_02742_));
 CLKBUF_X3 _08974_ (.A(_01942_),
    .Z(_02743_));
 MUX2_X1 _08975_ (.A(\registers[16][29] ),
    .B(\registers[17][29] ),
    .S(_02596_),
    .Z(_02744_));
 MUX2_X1 _08976_ (.A(\registers[22][29] ),
    .B(\registers[23][29] ),
    .S(_02515_),
    .Z(_02745_));
 OAI22_X2 _08977_ (.A1(_02513_),
    .A2(_02744_),
    .B1(_02745_),
    .B2(_02517_),
    .ZN(_02746_));
 MUX2_X1 _08978_ (.A(\registers[18][29] ),
    .B(\registers[19][29] ),
    .S(_02435_),
    .Z(_02747_));
 INV_X1 _08979_ (.A(_02747_),
    .ZN(_02748_));
 AOI21_X2 _08980_ (.A(_02746_),
    .B1(_02748_),
    .B2(_02709_),
    .ZN(_02749_));
 MUX2_X1 _08981_ (.A(\registers[20][29] ),
    .B(\registers[21][29] ),
    .S(_02639_),
    .Z(_02750_));
 INV_X1 _08982_ (.A(_02750_),
    .ZN(_02751_));
 AOI21_X1 _08983_ (.A(_02401_),
    .B1(_02711_),
    .B2(_02751_),
    .ZN(_02752_));
 MUX2_X1 _08984_ (.A(\registers[28][29] ),
    .B(\registers[30][29] ),
    .S(_02482_),
    .Z(_02753_));
 MUX2_X1 _08985_ (.A(\registers[29][29] ),
    .B(\registers[31][29] ),
    .S(_02526_),
    .Z(_02754_));
 MUX2_X1 _08986_ (.A(_02753_),
    .B(_02754_),
    .S(_02528_),
    .Z(_02755_));
 MUX2_X1 _08987_ (.A(\registers[24][29] ),
    .B(\registers[26][29] ),
    .S(_02571_),
    .Z(_02756_));
 MUX2_X1 _08988_ (.A(\registers[25][29] ),
    .B(\registers[27][29] ),
    .S(_02610_),
    .Z(_02757_));
 MUX2_X1 _08989_ (.A(_02756_),
    .B(_02757_),
    .S(_02574_),
    .Z(_02758_));
 MUX2_X1 _08990_ (.A(_02755_),
    .B(_02758_),
    .S(_02533_),
    .Z(_02759_));
 AOI221_X2 _08991_ (.A(_01860_),
    .B1(_02749_),
    .B2(_02752_),
    .C1(_02759_),
    .C2(_02722_),
    .ZN(_02760_));
 MUX2_X1 _08992_ (.A(\registers[0][29] ),
    .B(\registers[1][29] ),
    .S(_02043_),
    .Z(_02761_));
 NOR2_X1 _08993_ (.A1(_01913_),
    .A2(_02761_),
    .ZN(_02762_));
 MUX2_X1 _08994_ (.A(\registers[2][29] ),
    .B(\registers[3][29] ),
    .S(_01892_),
    .Z(_02763_));
 NOR3_X1 _08995_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_02763_),
    .ZN(_02764_));
 MUX2_X1 _08996_ (.A(\registers[4][29] ),
    .B(\registers[5][29] ),
    .S(_02150_),
    .Z(_02765_));
 NOR3_X1 _08997_ (.A1(_01921_),
    .A2(_01986_),
    .A3(_02765_),
    .ZN(_02766_));
 MUX2_X1 _08998_ (.A(\registers[6][29] ),
    .B(\registers[7][29] ),
    .S(_01951_),
    .Z(_02767_));
 NOR2_X1 _08999_ (.A1(_01924_),
    .A2(_02767_),
    .ZN(_02768_));
 NOR4_X1 _09000_ (.A1(_02762_),
    .A2(_02764_),
    .A3(_02766_),
    .A4(_02768_),
    .ZN(_02769_));
 MUX2_X1 _09001_ (.A(\registers[12][29] ),
    .B(\registers[14][29] ),
    .S(_02156_),
    .Z(_02770_));
 MUX2_X1 _09002_ (.A(\registers[13][29] ),
    .B(\registers[15][29] ),
    .S(_02158_),
    .Z(_02771_));
 MUX2_X1 _09003_ (.A(_02770_),
    .B(_02771_),
    .S(_02160_),
    .Z(_02772_));
 MUX2_X1 _09004_ (.A(\registers[8][29] ),
    .B(\registers[10][29] ),
    .S(_02162_),
    .Z(_02773_));
 MUX2_X1 _09005_ (.A(\registers[9][29] ),
    .B(\registers[11][29] ),
    .S(_02164_),
    .Z(_02774_));
 MUX2_X1 _09006_ (.A(_02773_),
    .B(_02774_),
    .S(_01931_),
    .Z(_02775_));
 MUX2_X1 _09007_ (.A(_02772_),
    .B(_02775_),
    .S(_01936_),
    .Z(_02776_));
 OAI221_X1 _09008_ (.A(_02724_),
    .B1(_01912_),
    .B2(_02769_),
    .C1(_02776_),
    .C2(_01939_),
    .ZN(_02777_));
 OAI22_X1 _09009_ (.A1(_02742_),
    .A2(_02743_),
    .B1(_02760_),
    .B2(_02777_),
    .ZN(_00350_));
 INV_X1 _09010_ (.A(net27),
    .ZN(_02778_));
 MUX2_X1 _09011_ (.A(\registers[16][2] ),
    .B(\registers[17][2] ),
    .S(_02596_),
    .Z(_02779_));
 MUX2_X1 _09012_ (.A(\registers[22][2] ),
    .B(\registers[23][2] ),
    .S(_02515_),
    .Z(_02780_));
 OAI22_X2 _09013_ (.A1(_02513_),
    .A2(_02779_),
    .B1(_02780_),
    .B2(_02517_),
    .ZN(_02781_));
 MUX2_X1 _09014_ (.A(\registers[18][2] ),
    .B(\registers[19][2] ),
    .S(_02435_),
    .Z(_02782_));
 INV_X1 _09015_ (.A(_02782_),
    .ZN(_02783_));
 AOI21_X2 _09016_ (.A(_02781_),
    .B1(_02783_),
    .B2(_02709_),
    .ZN(_02784_));
 CLKBUF_X3 _09017_ (.A(_01886_),
    .Z(_02785_));
 MUX2_X1 _09018_ (.A(\registers[20][2] ),
    .B(\registers[21][2] ),
    .S(_02639_),
    .Z(_02786_));
 INV_X1 _09019_ (.A(_02786_),
    .ZN(_02787_));
 AOI21_X1 _09020_ (.A(_02785_),
    .B1(_02711_),
    .B2(_02787_),
    .ZN(_02788_));
 MUX2_X1 _09021_ (.A(\registers[28][2] ),
    .B(\registers[30][2] ),
    .S(_02482_),
    .Z(_02789_));
 MUX2_X1 _09022_ (.A(\registers[29][2] ),
    .B(\registers[31][2] ),
    .S(_02526_),
    .Z(_02790_));
 MUX2_X1 _09023_ (.A(_02789_),
    .B(_02790_),
    .S(_02528_),
    .Z(_02791_));
 MUX2_X1 _09024_ (.A(\registers[24][2] ),
    .B(\registers[26][2] ),
    .S(_02571_),
    .Z(_02792_));
 MUX2_X1 _09025_ (.A(\registers[25][2] ),
    .B(\registers[27][2] ),
    .S(_02610_),
    .Z(_02793_));
 MUX2_X1 _09026_ (.A(_02792_),
    .B(_02793_),
    .S(_02574_),
    .Z(_02794_));
 MUX2_X1 _09027_ (.A(_02791_),
    .B(_02794_),
    .S(_02533_),
    .Z(_02795_));
 AOI221_X2 _09028_ (.A(_01860_),
    .B1(_02784_),
    .B2(_02788_),
    .C1(_02795_),
    .C2(_02722_),
    .ZN(_02796_));
 MUX2_X1 _09029_ (.A(\registers[0][2] ),
    .B(\registers[1][2] ),
    .S(_02043_),
    .Z(_02797_));
 NOR2_X1 _09030_ (.A1(_01913_),
    .A2(_02797_),
    .ZN(_02798_));
 MUX2_X1 _09031_ (.A(\registers[2][2] ),
    .B(\registers[3][2] ),
    .S(_01892_),
    .Z(_02799_));
 NOR3_X1 _09032_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_02799_),
    .ZN(_02800_));
 MUX2_X1 _09033_ (.A(\registers[4][2] ),
    .B(\registers[5][2] ),
    .S(_02150_),
    .Z(_02801_));
 NOR3_X1 _09034_ (.A1(_01921_),
    .A2(_01986_),
    .A3(_02801_),
    .ZN(_02802_));
 MUX2_X1 _09035_ (.A(\registers[6][2] ),
    .B(\registers[7][2] ),
    .S(_01951_),
    .Z(_02803_));
 NOR2_X1 _09036_ (.A1(_01924_),
    .A2(_02803_),
    .ZN(_02804_));
 NOR4_X1 _09037_ (.A1(_02798_),
    .A2(_02800_),
    .A3(_02802_),
    .A4(_02804_),
    .ZN(_02805_));
 MUX2_X1 _09038_ (.A(\registers[12][2] ),
    .B(\registers[14][2] ),
    .S(_02156_),
    .Z(_02806_));
 MUX2_X1 _09039_ (.A(\registers[13][2] ),
    .B(\registers[15][2] ),
    .S(_02158_),
    .Z(_02807_));
 MUX2_X1 _09040_ (.A(_02806_),
    .B(_02807_),
    .S(_02160_),
    .Z(_02808_));
 MUX2_X1 _09041_ (.A(\registers[8][2] ),
    .B(\registers[10][2] ),
    .S(_02162_),
    .Z(_02809_));
 MUX2_X1 _09042_ (.A(\registers[9][2] ),
    .B(\registers[11][2] ),
    .S(_02164_),
    .Z(_02810_));
 MUX2_X1 _09043_ (.A(_02809_),
    .B(_02810_),
    .S(_01931_),
    .Z(_02811_));
 MUX2_X1 _09044_ (.A(_02808_),
    .B(_02811_),
    .S(_01936_),
    .Z(_02812_));
 OAI221_X1 _09045_ (.A(_02724_),
    .B1(_01912_),
    .B2(_02805_),
    .C1(_02812_),
    .C2(_01939_),
    .ZN(_02813_));
 OAI22_X1 _09046_ (.A1(_02778_),
    .A2(_02743_),
    .B1(_02796_),
    .B2(_02813_),
    .ZN(_00351_));
 INV_X1 _09047_ (.A(net28),
    .ZN(_02814_));
 MUX2_X1 _09048_ (.A(\registers[0][30] ),
    .B(\registers[1][30] ),
    .S(_02596_),
    .Z(_02815_));
 MUX2_X1 _09049_ (.A(\registers[6][30] ),
    .B(\registers[7][30] ),
    .S(_02515_),
    .Z(_02816_));
 OAI22_X1 _09050_ (.A1(_02513_),
    .A2(_02815_),
    .B1(_02816_),
    .B2(_02517_),
    .ZN(_02817_));
 MUX2_X1 _09051_ (.A(\registers[2][30] ),
    .B(\registers[3][30] ),
    .S(_02029_),
    .Z(_02818_));
 INV_X1 _09052_ (.A(_02818_),
    .ZN(_02819_));
 AOI21_X1 _09053_ (.A(_02817_),
    .B1(_02819_),
    .B2(_02709_),
    .ZN(_02820_));
 MUX2_X1 _09054_ (.A(\registers[4][30] ),
    .B(\registers[5][30] ),
    .S(_02639_),
    .Z(_02821_));
 INV_X1 _09055_ (.A(_02821_),
    .ZN(_02822_));
 AOI21_X1 _09056_ (.A(_02785_),
    .B1(_02711_),
    .B2(_02822_),
    .ZN(_02823_));
 MUX2_X1 _09057_ (.A(\registers[12][30] ),
    .B(\registers[14][30] ),
    .S(_02482_),
    .Z(_02824_));
 MUX2_X1 _09058_ (.A(\registers[13][30] ),
    .B(\registers[15][30] ),
    .S(_02526_),
    .Z(_02825_));
 MUX2_X1 _09059_ (.A(_02824_),
    .B(_02825_),
    .S(_02528_),
    .Z(_02826_));
 MUX2_X1 _09060_ (.A(\registers[8][30] ),
    .B(\registers[10][30] ),
    .S(_02571_),
    .Z(_02827_));
 MUX2_X1 _09061_ (.A(\registers[9][30] ),
    .B(\registers[11][30] ),
    .S(_02610_),
    .Z(_02828_));
 MUX2_X1 _09062_ (.A(_02827_),
    .B(_02828_),
    .S(_02574_),
    .Z(_02829_));
 MUX2_X2 _09063_ (.A(_02826_),
    .B(_02829_),
    .S(_02533_),
    .Z(_02830_));
 AOI221_X2 _09064_ (.A(_02472_),
    .B1(_02820_),
    .B2(_02823_),
    .C1(_02830_),
    .C2(_02722_),
    .ZN(_02831_));
 MUX2_X1 _09065_ (.A(\registers[28][30] ),
    .B(\registers[30][30] ),
    .S(_02376_),
    .Z(_02832_));
 MUX2_X1 _09066_ (.A(\registers[29][30] ),
    .B(\registers[31][30] ),
    .S(_02414_),
    .Z(_02833_));
 MUX2_X1 _09067_ (.A(_02832_),
    .B(_02833_),
    .S(_02144_),
    .Z(_02834_));
 MUX2_X1 _09068_ (.A(\registers[24][30] ),
    .B(\registers[26][30] ),
    .S(_02453_),
    .Z(_02835_));
 MUX2_X1 _09069_ (.A(\registers[25][30] ),
    .B(\registers[27][30] ),
    .S(_02496_),
    .Z(_02836_));
 MUX2_X1 _09070_ (.A(_02835_),
    .B(_02836_),
    .S(_01979_),
    .Z(_02837_));
 MUX2_X1 _09071_ (.A(_02834_),
    .B(_02837_),
    .S(_02457_),
    .Z(_02838_));
 MUX2_X1 _09072_ (.A(\registers[16][30] ),
    .B(\registers[17][30] ),
    .S(_02459_),
    .Z(_02839_));
 NOR2_X1 _09073_ (.A1(_02543_),
    .A2(_02839_),
    .ZN(_02840_));
 MUX2_X1 _09074_ (.A(\registers[18][30] ),
    .B(\registers[19][30] ),
    .S(_01899_),
    .Z(_02841_));
 NOR3_X1 _09075_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_02841_),
    .ZN(_02842_));
 MUX2_X1 _09076_ (.A(\registers[20][30] ),
    .B(\registers[21][30] ),
    .S(_02504_),
    .Z(_02843_));
 NOR3_X1 _09077_ (.A1(_02550_),
    .A2(_02464_),
    .A3(_02843_),
    .ZN(_02844_));
 MUX2_X1 _09078_ (.A(\registers[22][30] ),
    .B(\registers[23][30] ),
    .S(_02035_),
    .Z(_02845_));
 NOR2_X1 _09079_ (.A1(_02553_),
    .A2(_02845_),
    .ZN(_02846_));
 NOR4_X2 _09080_ (.A1(_02840_),
    .A2(_02842_),
    .A3(_02844_),
    .A4(_02846_),
    .ZN(_02847_));
 OAI221_X1 _09081_ (.A(_02724_),
    .B1(_02491_),
    .B2(_02838_),
    .C1(_02847_),
    .C2(_02510_),
    .ZN(_02848_));
 OAI22_X1 _09082_ (.A1(_02814_),
    .A2(_02743_),
    .B1(_02831_),
    .B2(_02848_),
    .ZN(_00352_));
 INV_X1 _09083_ (.A(net29),
    .ZN(_02849_));
 MUX2_X1 _09084_ (.A(\registers[0][31] ),
    .B(\registers[1][31] ),
    .S(_02596_),
    .Z(_02850_));
 MUX2_X1 _09085_ (.A(\registers[6][31] ),
    .B(\registers[7][31] ),
    .S(_02515_),
    .Z(_02851_));
 OAI22_X1 _09086_ (.A1(_02513_),
    .A2(_02850_),
    .B1(_02851_),
    .B2(_02517_),
    .ZN(_02852_));
 MUX2_X1 _09087_ (.A(\registers[2][31] ),
    .B(\registers[3][31] ),
    .S(_02029_),
    .Z(_02853_));
 INV_X1 _09088_ (.A(_02853_),
    .ZN(_02854_));
 AOI21_X1 _09089_ (.A(_02852_),
    .B1(_02854_),
    .B2(_02709_),
    .ZN(_02855_));
 MUX2_X1 _09090_ (.A(\registers[4][31] ),
    .B(\registers[5][31] ),
    .S(_02639_),
    .Z(_02856_));
 INV_X1 _09091_ (.A(_02856_),
    .ZN(_02857_));
 AOI21_X1 _09092_ (.A(_02785_),
    .B1(_02711_),
    .B2(_02857_),
    .ZN(_02858_));
 MUX2_X1 _09093_ (.A(\registers[12][31] ),
    .B(\registers[14][31] ),
    .S(_01871_),
    .Z(_02859_));
 MUX2_X1 _09094_ (.A(\registers[13][31] ),
    .B(\registers[15][31] ),
    .S(_02526_),
    .Z(_02860_));
 MUX2_X1 _09095_ (.A(_02859_),
    .B(_02860_),
    .S(_02528_),
    .Z(_02861_));
 MUX2_X1 _09096_ (.A(\registers[8][31] ),
    .B(\registers[10][31] ),
    .S(_02571_),
    .Z(_02862_));
 MUX2_X1 _09097_ (.A(\registers[9][31] ),
    .B(\registers[11][31] ),
    .S(_02610_),
    .Z(_02863_));
 MUX2_X1 _09098_ (.A(_02862_),
    .B(_02863_),
    .S(_02574_),
    .Z(_02864_));
 MUX2_X1 _09099_ (.A(_02861_),
    .B(_02864_),
    .S(_02533_),
    .Z(_02865_));
 AOI221_X1 _09100_ (.A(_02472_),
    .B1(_02855_),
    .B2(_02858_),
    .C1(_02865_),
    .C2(_02722_),
    .ZN(_02866_));
 MUX2_X1 _09101_ (.A(\registers[28][31] ),
    .B(\registers[30][31] ),
    .S(_01881_),
    .Z(_02867_));
 MUX2_X1 _09102_ (.A(\registers[29][31] ),
    .B(\registers[31][31] ),
    .S(_02414_),
    .Z(_02868_));
 MUX2_X1 _09103_ (.A(_02867_),
    .B(_02868_),
    .S(_02144_),
    .Z(_02869_));
 MUX2_X1 _09104_ (.A(\registers[24][31] ),
    .B(\registers[26][31] ),
    .S(_02453_),
    .Z(_02870_));
 MUX2_X1 _09105_ (.A(\registers[25][31] ),
    .B(\registers[27][31] ),
    .S(_02496_),
    .Z(_02871_));
 MUX2_X1 _09106_ (.A(_02870_),
    .B(_02871_),
    .S(_01979_),
    .Z(_02872_));
 MUX2_X1 _09107_ (.A(_02869_),
    .B(_02872_),
    .S(_02457_),
    .Z(_02873_));
 MUX2_X1 _09108_ (.A(\registers[16][31] ),
    .B(\registers[17][31] ),
    .S(_02459_),
    .Z(_02874_));
 NOR2_X1 _09109_ (.A1(_02543_),
    .A2(_02874_),
    .ZN(_02875_));
 MUX2_X1 _09110_ (.A(\registers[18][31] ),
    .B(\registers[19][31] ),
    .S(_01899_),
    .Z(_02876_));
 NOR3_X1 _09111_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_02876_),
    .ZN(_02877_));
 MUX2_X1 _09112_ (.A(\registers[20][31] ),
    .B(\registers[21][31] ),
    .S(_02504_),
    .Z(_02878_));
 NOR3_X1 _09113_ (.A1(_02550_),
    .A2(_02464_),
    .A3(_02878_),
    .ZN(_02879_));
 MUX2_X1 _09114_ (.A(\registers[22][31] ),
    .B(\registers[23][31] ),
    .S(_02035_),
    .Z(_02880_));
 NOR2_X1 _09115_ (.A1(_02553_),
    .A2(_02880_),
    .ZN(_02881_));
 NOR4_X2 _09116_ (.A1(_02875_),
    .A2(_02877_),
    .A3(_02879_),
    .A4(_02881_),
    .ZN(_02882_));
 OAI221_X1 _09117_ (.A(_02724_),
    .B1(_02491_),
    .B2(_02873_),
    .C1(_02882_),
    .C2(_02510_),
    .ZN(_02883_));
 OAI22_X1 _09118_ (.A1(_02849_),
    .A2(_02743_),
    .B1(_02866_),
    .B2(_02883_),
    .ZN(_00353_));
 INV_X1 _09119_ (.A(net30),
    .ZN(_02884_));
 MUX2_X1 _09120_ (.A(\registers[0][3] ),
    .B(\registers[1][3] ),
    .S(_02596_),
    .Z(_02885_));
 MUX2_X1 _09121_ (.A(\registers[6][3] ),
    .B(\registers[7][3] ),
    .S(_01898_),
    .Z(_02886_));
 OAI22_X2 _09122_ (.A1(_01865_),
    .A2(_02885_),
    .B1(_02886_),
    .B2(_01872_),
    .ZN(_02887_));
 MUX2_X1 _09123_ (.A(\registers[2][3] ),
    .B(\registers[3][3] ),
    .S(_02029_),
    .Z(_02888_));
 INV_X1 _09124_ (.A(_02888_),
    .ZN(_02889_));
 AOI21_X1 _09125_ (.A(_02887_),
    .B1(_02889_),
    .B2(_02709_),
    .ZN(_02890_));
 MUX2_X1 _09126_ (.A(\registers[4][3] ),
    .B(\registers[5][3] ),
    .S(_02639_),
    .Z(_02891_));
 INV_X1 _09127_ (.A(_02891_),
    .ZN(_02892_));
 AOI21_X1 _09128_ (.A(_02785_),
    .B1(_02711_),
    .B2(_02892_),
    .ZN(_02893_));
 MUX2_X1 _09129_ (.A(\registers[12][3] ),
    .B(\registers[14][3] ),
    .S(_01871_),
    .Z(_02894_));
 MUX2_X1 _09130_ (.A(\registers[13][3] ),
    .B(\registers[15][3] ),
    .S(_01960_),
    .Z(_02895_));
 MUX2_X1 _09131_ (.A(_02894_),
    .B(_02895_),
    .S(_01995_),
    .Z(_02896_));
 MUX2_X1 _09132_ (.A(\registers[8][3] ),
    .B(\registers[10][3] ),
    .S(_02571_),
    .Z(_02897_));
 MUX2_X1 _09133_ (.A(\registers[9][3] ),
    .B(\registers[11][3] ),
    .S(_02610_),
    .Z(_02898_));
 MUX2_X1 _09134_ (.A(_02897_),
    .B(_02898_),
    .S(_02574_),
    .Z(_02899_));
 MUX2_X2 _09135_ (.A(_02896_),
    .B(_02899_),
    .S(_02149_),
    .Z(_02900_));
 AOI221_X2 _09136_ (.A(_02472_),
    .B1(_02890_),
    .B2(_02893_),
    .C1(_02900_),
    .C2(_02722_),
    .ZN(_02901_));
 MUX2_X1 _09137_ (.A(\registers[28][3] ),
    .B(\registers[30][3] ),
    .S(_01881_),
    .Z(_02902_));
 MUX2_X1 _09138_ (.A(\registers[29][3] ),
    .B(\registers[31][3] ),
    .S(_01975_),
    .Z(_02903_));
 MUX2_X1 _09139_ (.A(_02902_),
    .B(_02903_),
    .S(_02144_),
    .Z(_02904_));
 MUX2_X1 _09140_ (.A(\registers[24][3] ),
    .B(\registers[26][3] ),
    .S(_02453_),
    .Z(_02905_));
 MUX2_X1 _09141_ (.A(\registers[25][3] ),
    .B(\registers[27][3] ),
    .S(_02496_),
    .Z(_02906_));
 MUX2_X1 _09142_ (.A(_02905_),
    .B(_02906_),
    .S(_01979_),
    .Z(_02907_));
 MUX2_X1 _09143_ (.A(_02904_),
    .B(_02907_),
    .S(_02457_),
    .Z(_02908_));
 MUX2_X1 _09144_ (.A(\registers[16][3] ),
    .B(\registers[17][3] ),
    .S(_02459_),
    .Z(_02909_));
 NOR2_X1 _09145_ (.A1(_02543_),
    .A2(_02909_),
    .ZN(_02910_));
 MUX2_X1 _09146_ (.A(\registers[18][3] ),
    .B(\registers[19][3] ),
    .S(_01899_),
    .Z(_02911_));
 NOR3_X1 _09147_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_02911_),
    .ZN(_02912_));
 MUX2_X1 _09148_ (.A(\registers[20][3] ),
    .B(\registers[21][3] ),
    .S(_02504_),
    .Z(_02913_));
 NOR3_X1 _09149_ (.A1(_02550_),
    .A2(_02464_),
    .A3(_02913_),
    .ZN(_02914_));
 MUX2_X1 _09150_ (.A(\registers[22][3] ),
    .B(\registers[23][3] ),
    .S(_02035_),
    .Z(_02915_));
 NOR2_X1 _09151_ (.A1(_02553_),
    .A2(_02915_),
    .ZN(_02916_));
 NOR4_X2 _09152_ (.A1(_02910_),
    .A2(_02912_),
    .A3(_02914_),
    .A4(_02916_),
    .ZN(_02917_));
 OAI221_X1 _09153_ (.A(_02724_),
    .B1(_02491_),
    .B2(_02908_),
    .C1(_02917_),
    .C2(_02510_),
    .ZN(_02918_));
 OAI22_X1 _09154_ (.A1(_02884_),
    .A2(_02743_),
    .B1(_02901_),
    .B2(_02918_),
    .ZN(_00354_));
 INV_X1 _09155_ (.A(net31),
    .ZN(_02919_));
 MUX2_X1 _09156_ (.A(\registers[0][4] ),
    .B(\registers[1][4] ),
    .S(_02596_),
    .Z(_02920_));
 MUX2_X1 _09157_ (.A(\registers[6][4] ),
    .B(\registers[7][4] ),
    .S(_01898_),
    .Z(_02921_));
 OAI22_X2 _09158_ (.A1(_01865_),
    .A2(_02920_),
    .B1(_02921_),
    .B2(_01872_),
    .ZN(_02922_));
 MUX2_X1 _09159_ (.A(\registers[2][4] ),
    .B(\registers[3][4] ),
    .S(_02029_),
    .Z(_02923_));
 INV_X1 _09160_ (.A(_02923_),
    .ZN(_02924_));
 AOI21_X1 _09161_ (.A(_02922_),
    .B1(_02924_),
    .B2(_02709_),
    .ZN(_02925_));
 MUX2_X1 _09162_ (.A(\registers[4][4] ),
    .B(\registers[5][4] ),
    .S(_02639_),
    .Z(_02926_));
 INV_X1 _09163_ (.A(_02926_),
    .ZN(_02927_));
 AOI21_X1 _09164_ (.A(_02785_),
    .B1(_02711_),
    .B2(_02927_),
    .ZN(_02928_));
 MUX2_X1 _09165_ (.A(\registers[12][4] ),
    .B(\registers[14][4] ),
    .S(_01871_),
    .Z(_02929_));
 MUX2_X1 _09166_ (.A(\registers[13][4] ),
    .B(\registers[15][4] ),
    .S(_01960_),
    .Z(_02930_));
 MUX2_X1 _09167_ (.A(_02929_),
    .B(_02930_),
    .S(_01995_),
    .Z(_02931_));
 MUX2_X1 _09168_ (.A(\registers[8][4] ),
    .B(\registers[10][4] ),
    .S(_01962_),
    .Z(_02932_));
 MUX2_X1 _09169_ (.A(\registers[9][4] ),
    .B(\registers[11][4] ),
    .S(_02610_),
    .Z(_02933_));
 MUX2_X1 _09170_ (.A(_02932_),
    .B(_02933_),
    .S(_01964_),
    .Z(_02934_));
 MUX2_X2 _09171_ (.A(_02931_),
    .B(_02934_),
    .S(_02149_),
    .Z(_02935_));
 AOI221_X2 _09172_ (.A(_02472_),
    .B1(_02925_),
    .B2(_02928_),
    .C1(_02935_),
    .C2(_02722_),
    .ZN(_02936_));
 MUX2_X1 _09173_ (.A(\registers[28][4] ),
    .B(\registers[30][4] ),
    .S(_01881_),
    .Z(_02937_));
 MUX2_X1 _09174_ (.A(\registers[29][4] ),
    .B(\registers[31][4] ),
    .S(_01975_),
    .Z(_02938_));
 MUX2_X1 _09175_ (.A(_02937_),
    .B(_02938_),
    .S(_02144_),
    .Z(_02939_));
 MUX2_X1 _09176_ (.A(\registers[24][4] ),
    .B(\registers[26][4] ),
    .S(_01977_),
    .Z(_02940_));
 MUX2_X1 _09177_ (.A(\registers[25][4] ),
    .B(\registers[27][4] ),
    .S(_02496_),
    .Z(_02941_));
 MUX2_X1 _09178_ (.A(_02940_),
    .B(_02941_),
    .S(_01979_),
    .Z(_02942_));
 MUX2_X1 _09179_ (.A(_02939_),
    .B(_02942_),
    .S(_02039_),
    .Z(_02943_));
 MUX2_X1 _09180_ (.A(\registers[16][4] ),
    .B(\registers[17][4] ),
    .S(_01914_),
    .Z(_02944_));
 NOR2_X1 _09181_ (.A1(_02543_),
    .A2(_02944_),
    .ZN(_02945_));
 MUX2_X1 _09182_ (.A(\registers[18][4] ),
    .B(\registers[19][4] ),
    .S(_01899_),
    .Z(_02946_));
 NOR3_X1 _09183_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_02946_),
    .ZN(_02947_));
 MUX2_X1 _09184_ (.A(\registers[20][4] ),
    .B(\registers[21][4] ),
    .S(_02504_),
    .Z(_02948_));
 NOR3_X1 _09185_ (.A1(_02550_),
    .A2(_01904_),
    .A3(_02948_),
    .ZN(_02949_));
 MUX2_X1 _09186_ (.A(\registers[22][4] ),
    .B(\registers[23][4] ),
    .S(_02035_),
    .Z(_02950_));
 NOR2_X1 _09187_ (.A1(_02553_),
    .A2(_02950_),
    .ZN(_02951_));
 NOR4_X2 _09188_ (.A1(_02945_),
    .A2(_02947_),
    .A3(_02949_),
    .A4(_02951_),
    .ZN(_02952_));
 OAI221_X1 _09189_ (.A(_02724_),
    .B1(_02491_),
    .B2(_02943_),
    .C1(_02952_),
    .C2(_02510_),
    .ZN(_02953_));
 OAI22_X1 _09190_ (.A1(_02919_),
    .A2(_02743_),
    .B1(_02936_),
    .B2(_02953_),
    .ZN(_00355_));
 INV_X1 _09191_ (.A(net32),
    .ZN(_02954_));
 MUX2_X1 _09192_ (.A(\registers[16][5] ),
    .B(\registers[17][5] ),
    .S(_01874_),
    .Z(_02955_));
 MUX2_X1 _09193_ (.A(\registers[22][5] ),
    .B(\registers[23][5] ),
    .S(_01898_),
    .Z(_02956_));
 OAI22_X1 _09194_ (.A1(_01865_),
    .A2(_02955_),
    .B1(_02956_),
    .B2(_01872_),
    .ZN(_02957_));
 MUX2_X1 _09195_ (.A(\registers[18][5] ),
    .B(\registers[19][5] ),
    .S(_02029_),
    .Z(_02958_));
 INV_X1 _09196_ (.A(_02958_),
    .ZN(_02959_));
 AOI21_X2 _09197_ (.A(_02957_),
    .B1(_02959_),
    .B2(_02709_),
    .ZN(_02960_));
 MUX2_X1 _09198_ (.A(\registers[20][5] ),
    .B(\registers[21][5] ),
    .S(_02639_),
    .Z(_02961_));
 INV_X1 _09199_ (.A(_02961_),
    .ZN(_02962_));
 AOI21_X1 _09200_ (.A(_02785_),
    .B1(_02711_),
    .B2(_02962_),
    .ZN(_02963_));
 MUX2_X1 _09201_ (.A(\registers[28][5] ),
    .B(\registers[30][5] ),
    .S(_01871_),
    .Z(_02964_));
 MUX2_X1 _09202_ (.A(\registers[29][5] ),
    .B(\registers[31][5] ),
    .S(_01960_),
    .Z(_02965_));
 MUX2_X1 _09203_ (.A(_02964_),
    .B(_02965_),
    .S(_01995_),
    .Z(_02966_));
 MUX2_X1 _09204_ (.A(\registers[24][5] ),
    .B(\registers[26][5] ),
    .S(_01962_),
    .Z(_02967_));
 MUX2_X1 _09205_ (.A(\registers[25][5] ),
    .B(\registers[27][5] ),
    .S(_01966_),
    .Z(_02968_));
 MUX2_X1 _09206_ (.A(_02967_),
    .B(_02968_),
    .S(_01964_),
    .Z(_02969_));
 MUX2_X1 _09207_ (.A(_02966_),
    .B(_02969_),
    .S(_02149_),
    .Z(_02970_));
 AOI221_X2 _09208_ (.A(_01860_),
    .B1(_02960_),
    .B2(_02963_),
    .C1(_02970_),
    .C2(_02722_),
    .ZN(_02971_));
 MUX2_X1 _09209_ (.A(\registers[0][5] ),
    .B(\registers[1][5] ),
    .S(_02043_),
    .Z(_02972_));
 NOR2_X1 _09210_ (.A1(_01913_),
    .A2(_02972_),
    .ZN(_02973_));
 MUX2_X1 _09211_ (.A(\registers[2][5] ),
    .B(\registers[3][5] ),
    .S(_01892_),
    .Z(_02974_));
 NOR3_X1 _09212_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_02974_),
    .ZN(_02975_));
 MUX2_X1 _09213_ (.A(\registers[4][5] ),
    .B(\registers[5][5] ),
    .S(_02150_),
    .Z(_02976_));
 NOR3_X1 _09214_ (.A1(_01921_),
    .A2(_01986_),
    .A3(_02976_),
    .ZN(_02977_));
 MUX2_X1 _09215_ (.A(\registers[6][5] ),
    .B(\registers[7][5] ),
    .S(_01951_),
    .Z(_02978_));
 NOR2_X1 _09216_ (.A1(_01924_),
    .A2(_02978_),
    .ZN(_02979_));
 NOR4_X1 _09217_ (.A1(_02973_),
    .A2(_02975_),
    .A3(_02977_),
    .A4(_02979_),
    .ZN(_02980_));
 MUX2_X1 _09218_ (.A(\registers[12][5] ),
    .B(\registers[14][5] ),
    .S(_02156_),
    .Z(_02981_));
 MUX2_X1 _09219_ (.A(\registers[13][5] ),
    .B(\registers[15][5] ),
    .S(_02158_),
    .Z(_02982_));
 MUX2_X1 _09220_ (.A(_02981_),
    .B(_02982_),
    .S(_02160_),
    .Z(_02983_));
 MUX2_X1 _09221_ (.A(\registers[8][5] ),
    .B(\registers[10][5] ),
    .S(_02162_),
    .Z(_02984_));
 MUX2_X1 _09222_ (.A(\registers[9][5] ),
    .B(\registers[11][5] ),
    .S(_02164_),
    .Z(_02985_));
 MUX2_X1 _09223_ (.A(_02984_),
    .B(_02985_),
    .S(_01931_),
    .Z(_02986_));
 MUX2_X1 _09224_ (.A(_02983_),
    .B(_02986_),
    .S(_01936_),
    .Z(_02987_));
 OAI221_X1 _09225_ (.A(_02724_),
    .B1(_01912_),
    .B2(_02980_),
    .C1(_02987_),
    .C2(_01939_),
    .ZN(_02988_));
 OAI22_X1 _09226_ (.A1(_02954_),
    .A2(_02743_),
    .B1(_02971_),
    .B2(_02988_),
    .ZN(_00356_));
 INV_X1 _09227_ (.A(net33),
    .ZN(_02989_));
 MUX2_X1 _09228_ (.A(\registers[16][6] ),
    .B(\registers[17][6] ),
    .S(_01874_),
    .Z(_02990_));
 MUX2_X1 _09229_ (.A(\registers[22][6] ),
    .B(\registers[23][6] ),
    .S(_01898_),
    .Z(_02991_));
 OAI22_X1 _09230_ (.A1(_01865_),
    .A2(_02990_),
    .B1(_02991_),
    .B2(_01872_),
    .ZN(_02992_));
 MUX2_X1 _09231_ (.A(\registers[18][6] ),
    .B(\registers[19][6] ),
    .S(_02029_),
    .Z(_02993_));
 INV_X1 _09232_ (.A(_02993_),
    .ZN(_02994_));
 AOI21_X2 _09233_ (.A(_02992_),
    .B1(_02994_),
    .B2(_02709_),
    .ZN(_02995_));
 MUX2_X1 _09234_ (.A(\registers[20][6] ),
    .B(\registers[21][6] ),
    .S(_01869_),
    .Z(_02996_));
 INV_X1 _09235_ (.A(_02996_),
    .ZN(_02997_));
 AOI21_X1 _09236_ (.A(_02785_),
    .B1(_02711_),
    .B2(_02997_),
    .ZN(_02998_));
 MUX2_X1 _09237_ (.A(\registers[28][6] ),
    .B(\registers[30][6] ),
    .S(_01871_),
    .Z(_02999_));
 MUX2_X1 _09238_ (.A(\registers[29][6] ),
    .B(\registers[31][6] ),
    .S(_01960_),
    .Z(_03000_));
 MUX2_X1 _09239_ (.A(_02999_),
    .B(_03000_),
    .S(_01995_),
    .Z(_03001_));
 MUX2_X1 _09240_ (.A(\registers[24][6] ),
    .B(\registers[26][6] ),
    .S(_01962_),
    .Z(_03002_));
 MUX2_X1 _09241_ (.A(\registers[25][6] ),
    .B(\registers[27][6] ),
    .S(_01966_),
    .Z(_03003_));
 MUX2_X1 _09242_ (.A(_03002_),
    .B(_03003_),
    .S(_01964_),
    .Z(_03004_));
 MUX2_X1 _09243_ (.A(_03001_),
    .B(_03004_),
    .S(_02149_),
    .Z(_03005_));
 AOI221_X2 _09244_ (.A(_01860_),
    .B1(_02995_),
    .B2(_02998_),
    .C1(_03005_),
    .C2(_02722_),
    .ZN(_03006_));
 MUX2_X1 _09245_ (.A(\registers[0][6] ),
    .B(\registers[1][6] ),
    .S(_02043_),
    .Z(_03007_));
 NOR2_X1 _09246_ (.A1(_01913_),
    .A2(_03007_),
    .ZN(_03008_));
 MUX2_X1 _09247_ (.A(\registers[2][6] ),
    .B(\registers[3][6] ),
    .S(_02150_),
    .Z(_03009_));
 NOR3_X1 _09248_ (.A1(_01917_),
    .A2(_01918_),
    .A3(_03009_),
    .ZN(_03010_));
 MUX2_X1 _09249_ (.A(\registers[4][6] ),
    .B(\registers[5][6] ),
    .S(_01955_),
    .Z(_03011_));
 NOR3_X1 _09250_ (.A1(_01921_),
    .A2(_01986_),
    .A3(_03011_),
    .ZN(_03012_));
 MUX2_X1 _09251_ (.A(\registers[6][6] ),
    .B(\registers[7][6] ),
    .S(_01951_),
    .Z(_03013_));
 NOR2_X1 _09252_ (.A1(_01924_),
    .A2(_03013_),
    .ZN(_03014_));
 NOR4_X1 _09253_ (.A1(_03008_),
    .A2(_03010_),
    .A3(_03012_),
    .A4(_03014_),
    .ZN(_03015_));
 MUX2_X1 _09254_ (.A(\registers[12][6] ),
    .B(\registers[14][6] ),
    .S(_02156_),
    .Z(_03016_));
 MUX2_X1 _09255_ (.A(\registers[13][6] ),
    .B(\registers[15][6] ),
    .S(_02158_),
    .Z(_03017_));
 MUX2_X1 _09256_ (.A(_03016_),
    .B(_03017_),
    .S(_02160_),
    .Z(_03018_));
 MUX2_X1 _09257_ (.A(\registers[8][6] ),
    .B(\registers[10][6] ),
    .S(_02162_),
    .Z(_03019_));
 MUX2_X1 _09258_ (.A(\registers[9][6] ),
    .B(\registers[11][6] ),
    .S(_02164_),
    .Z(_03020_));
 MUX2_X1 _09259_ (.A(_03019_),
    .B(_03020_),
    .S(_01931_),
    .Z(_03021_));
 MUX2_X1 _09260_ (.A(_03018_),
    .B(_03021_),
    .S(_01936_),
    .Z(_03022_));
 OAI221_X1 _09261_ (.A(_02724_),
    .B1(_01912_),
    .B2(_03015_),
    .C1(_03022_),
    .C2(_01939_),
    .ZN(_03023_));
 OAI22_X1 _09262_ (.A1(_02989_),
    .A2(_02743_),
    .B1(_03006_),
    .B2(_03023_),
    .ZN(_00357_));
 INV_X1 _09263_ (.A(net34),
    .ZN(_03024_));
 MUX2_X1 _09264_ (.A(\registers[16][7] ),
    .B(\registers[17][7] ),
    .S(_01874_),
    .Z(_03025_));
 MUX2_X1 _09265_ (.A(\registers[22][7] ),
    .B(\registers[23][7] ),
    .S(_01898_),
    .Z(_03026_));
 OAI22_X1 _09266_ (.A1(_01865_),
    .A2(_03025_),
    .B1(_03026_),
    .B2(_01872_),
    .ZN(_03027_));
 MUX2_X1 _09267_ (.A(\registers[18][7] ),
    .B(\registers[19][7] ),
    .S(_02029_),
    .Z(_03028_));
 INV_X1 _09268_ (.A(_03028_),
    .ZN(_03029_));
 AOI21_X2 _09269_ (.A(_03027_),
    .B1(_03029_),
    .B2(_02709_),
    .ZN(_03030_));
 MUX2_X1 _09270_ (.A(\registers[20][7] ),
    .B(\registers[21][7] ),
    .S(_01869_),
    .Z(_03031_));
 INV_X1 _09271_ (.A(_03031_),
    .ZN(_03032_));
 AOI21_X1 _09272_ (.A(_02785_),
    .B1(_02711_),
    .B2(_03032_),
    .ZN(_03033_));
 MUX2_X1 _09273_ (.A(\registers[28][7] ),
    .B(\registers[30][7] ),
    .S(_01871_),
    .Z(_03034_));
 MUX2_X1 _09274_ (.A(\registers[29][7] ),
    .B(\registers[31][7] ),
    .S(_01960_),
    .Z(_03035_));
 MUX2_X1 _09275_ (.A(_03034_),
    .B(_03035_),
    .S(_01995_),
    .Z(_03036_));
 MUX2_X1 _09276_ (.A(\registers[24][7] ),
    .B(\registers[26][7] ),
    .S(_01962_),
    .Z(_03037_));
 MUX2_X1 _09277_ (.A(\registers[25][7] ),
    .B(\registers[27][7] ),
    .S(_01966_),
    .Z(_03038_));
 MUX2_X1 _09278_ (.A(_03037_),
    .B(_03038_),
    .S(_01964_),
    .Z(_03039_));
 MUX2_X1 _09279_ (.A(_03036_),
    .B(_03039_),
    .S(_02149_),
    .Z(_03040_));
 AOI221_X2 _09280_ (.A(_01860_),
    .B1(_03030_),
    .B2(_03033_),
    .C1(_03040_),
    .C2(_02722_),
    .ZN(_03041_));
 MUX2_X1 _09281_ (.A(\registers[0][7] ),
    .B(\registers[1][7] ),
    .S(_02043_),
    .Z(_03042_));
 NOR2_X1 _09282_ (.A1(_01866_),
    .A2(_03042_),
    .ZN(_03043_));
 MUX2_X1 _09283_ (.A(\registers[2][7] ),
    .B(\registers[3][7] ),
    .S(_02150_),
    .Z(_03044_));
 NOR3_X1 _09284_ (.A1(_01882_),
    .A2(_01863_),
    .A3(_03044_),
    .ZN(_03045_));
 MUX2_X1 _09285_ (.A(\registers[4][7] ),
    .B(\registers[5][7] ),
    .S(_01955_),
    .Z(_03046_));
 NOR3_X1 _09286_ (.A1(_01888_),
    .A2(_01986_),
    .A3(_03046_),
    .ZN(_03047_));
 MUX2_X1 _09287_ (.A(\registers[6][7] ),
    .B(\registers[7][7] ),
    .S(_01951_),
    .Z(_03048_));
 NOR2_X1 _09288_ (.A1(_01873_),
    .A2(_03048_),
    .ZN(_03049_));
 NOR4_X1 _09289_ (.A1(_03043_),
    .A2(_03045_),
    .A3(_03047_),
    .A4(_03049_),
    .ZN(_03050_));
 MUX2_X1 _09290_ (.A(\registers[12][7] ),
    .B(\registers[14][7] ),
    .S(_02156_),
    .Z(_03051_));
 MUX2_X1 _09291_ (.A(\registers[13][7] ),
    .B(\registers[15][7] ),
    .S(_02158_),
    .Z(_03052_));
 MUX2_X1 _09292_ (.A(_03051_),
    .B(_03052_),
    .S(_02030_),
    .Z(_03053_));
 MUX2_X1 _09293_ (.A(\registers[8][7] ),
    .B(\registers[10][7] ),
    .S(_02162_),
    .Z(_03054_));
 MUX2_X1 _09294_ (.A(\registers[9][7] ),
    .B(\registers[11][7] ),
    .S(_02164_),
    .Z(_03055_));
 MUX2_X1 _09295_ (.A(_03054_),
    .B(_03055_),
    .S(_02160_),
    .Z(_03056_));
 MUX2_X1 _09296_ (.A(_03053_),
    .B(_03056_),
    .S(_01936_),
    .Z(_03057_));
 OAI221_X1 _09297_ (.A(_02724_),
    .B1(_01912_),
    .B2(_03050_),
    .C1(_03057_),
    .C2(_01939_),
    .ZN(_03058_));
 OAI22_X1 _09298_ (.A1(_03024_),
    .A2(_02743_),
    .B1(_03041_),
    .B2(_03058_),
    .ZN(_00358_));
 INV_X1 _09299_ (.A(net35),
    .ZN(_03059_));
 MUX2_X1 _09300_ (.A(\registers[0][8] ),
    .B(\registers[1][8] ),
    .S(_01874_),
    .Z(_03060_));
 MUX2_X1 _09301_ (.A(\registers[6][8] ),
    .B(\registers[7][8] ),
    .S(_01898_),
    .Z(_03061_));
 OAI22_X1 _09302_ (.A1(_01865_),
    .A2(_03060_),
    .B1(_03061_),
    .B2(_01872_),
    .ZN(_03062_));
 MUX2_X1 _09303_ (.A(\registers[2][8] ),
    .B(\registers[3][8] ),
    .S(_02029_),
    .Z(_03063_));
 INV_X1 _09304_ (.A(_03063_),
    .ZN(_03064_));
 AOI21_X1 _09305_ (.A(_03062_),
    .B1(_03064_),
    .B2(_01883_),
    .ZN(_03065_));
 MUX2_X1 _09306_ (.A(\registers[4][8] ),
    .B(\registers[5][8] ),
    .S(_01869_),
    .Z(_03066_));
 INV_X1 _09307_ (.A(_03066_),
    .ZN(_03067_));
 AOI21_X1 _09308_ (.A(_02785_),
    .B1(_01890_),
    .B2(_03067_),
    .ZN(_03068_));
 MUX2_X1 _09309_ (.A(\registers[12][8] ),
    .B(\registers[14][8] ),
    .S(_01871_),
    .Z(_03069_));
 MUX2_X1 _09310_ (.A(\registers[13][8] ),
    .B(\registers[15][8] ),
    .S(_01960_),
    .Z(_03070_));
 MUX2_X1 _09311_ (.A(_03069_),
    .B(_03070_),
    .S(_01995_),
    .Z(_03071_));
 MUX2_X1 _09312_ (.A(\registers[8][8] ),
    .B(\registers[10][8] ),
    .S(_01962_),
    .Z(_03072_));
 MUX2_X1 _09313_ (.A(\registers[9][8] ),
    .B(\registers[11][8] ),
    .S(_01966_),
    .Z(_03073_));
 MUX2_X1 _09314_ (.A(_03072_),
    .B(_03073_),
    .S(_01964_),
    .Z(_03074_));
 MUX2_X2 _09315_ (.A(_03071_),
    .B(_03074_),
    .S(_02149_),
    .Z(_03075_));
 AOI221_X2 _09316_ (.A(_01858_),
    .B1(_03065_),
    .B2(_03068_),
    .C1(_03075_),
    .C2(_01887_),
    .ZN(_03076_));
 MUX2_X1 _09317_ (.A(\registers[28][8] ),
    .B(\registers[30][8] ),
    .S(_01881_),
    .Z(_03077_));
 MUX2_X1 _09318_ (.A(\registers[29][8] ),
    .B(\registers[31][8] ),
    .S(_01975_),
    .Z(_03078_));
 MUX2_X1 _09319_ (.A(_03077_),
    .B(_03078_),
    .S(_02144_),
    .Z(_03079_));
 MUX2_X1 _09320_ (.A(\registers[24][8] ),
    .B(\registers[26][8] ),
    .S(_01977_),
    .Z(_03080_));
 MUX2_X1 _09321_ (.A(\registers[25][8] ),
    .B(\registers[27][8] ),
    .S(_01981_),
    .Z(_03081_));
 MUX2_X1 _09322_ (.A(_03080_),
    .B(_03081_),
    .S(_01979_),
    .Z(_03082_));
 MUX2_X1 _09323_ (.A(_03079_),
    .B(_03082_),
    .S(_02039_),
    .Z(_03083_));
 MUX2_X1 _09324_ (.A(\registers[16][8] ),
    .B(\registers[17][8] ),
    .S(_01914_),
    .Z(_03084_));
 NOR2_X1 _09325_ (.A1(_02543_),
    .A2(_03084_),
    .ZN(_03085_));
 MUX2_X1 _09326_ (.A(\registers[18][8] ),
    .B(\registers[19][8] ),
    .S(_01899_),
    .Z(_03086_));
 NOR3_X1 _09327_ (.A1(_02546_),
    .A2(_02547_),
    .A3(_03086_),
    .ZN(_03087_));
 MUX2_X1 _09328_ (.A(\registers[20][8] ),
    .B(\registers[21][8] ),
    .S(_01878_),
    .Z(_03088_));
 NOR3_X1 _09329_ (.A1(_02550_),
    .A2(_01904_),
    .A3(_03088_),
    .ZN(_03089_));
 MUX2_X1 _09330_ (.A(\registers[22][8] ),
    .B(\registers[23][8] ),
    .S(_02035_),
    .Z(_03090_));
 NOR2_X1 _09331_ (.A1(_02553_),
    .A2(_03090_),
    .ZN(_03091_));
 NOR4_X2 _09332_ (.A1(_03085_),
    .A2(_03087_),
    .A3(_03089_),
    .A4(_03091_),
    .ZN(_03092_));
 OAI221_X1 _09333_ (.A(_01909_),
    .B1(_01973_),
    .B2(_03083_),
    .C1(_03092_),
    .C2(_01989_),
    .ZN(_03093_));
 OAI22_X1 _09334_ (.A1(_03059_),
    .A2(_02743_),
    .B1(_03076_),
    .B2(_03093_),
    .ZN(_00359_));
 INV_X1 _09335_ (.A(net36),
    .ZN(_03094_));
 MUX2_X1 _09336_ (.A(\registers[16][9] ),
    .B(\registers[17][9] ),
    .S(_01874_),
    .Z(_03095_));
 MUX2_X1 _09337_ (.A(\registers[22][9] ),
    .B(\registers[23][9] ),
    .S(_01898_),
    .Z(_03096_));
 OAI22_X1 _09338_ (.A1(_01865_),
    .A2(_03095_),
    .B1(_03096_),
    .B2(_01872_),
    .ZN(_03097_));
 MUX2_X1 _09339_ (.A(\registers[18][9] ),
    .B(\registers[19][9] ),
    .S(_02029_),
    .Z(_03098_));
 INV_X1 _09340_ (.A(_03098_),
    .ZN(_03099_));
 AOI21_X1 _09341_ (.A(_03097_),
    .B1(_03099_),
    .B2(_01883_),
    .ZN(_03100_));
 MUX2_X1 _09342_ (.A(\registers[20][9] ),
    .B(\registers[21][9] ),
    .S(_01869_),
    .Z(_03101_));
 INV_X1 _09343_ (.A(_03101_),
    .ZN(_03102_));
 AOI21_X1 _09344_ (.A(_02785_),
    .B1(_01890_),
    .B2(_03102_),
    .ZN(_03103_));
 MUX2_X1 _09345_ (.A(\registers[28][9] ),
    .B(\registers[30][9] ),
    .S(_01871_),
    .Z(_03104_));
 MUX2_X1 _09346_ (.A(\registers[29][9] ),
    .B(\registers[31][9] ),
    .S(_01960_),
    .Z(_03105_));
 MUX2_X1 _09347_ (.A(_03104_),
    .B(_03105_),
    .S(_01995_),
    .Z(_03106_));
 MUX2_X1 _09348_ (.A(\registers[24][9] ),
    .B(\registers[26][9] ),
    .S(_01962_),
    .Z(_03107_));
 MUX2_X1 _09349_ (.A(\registers[25][9] ),
    .B(\registers[27][9] ),
    .S(_01966_),
    .Z(_03108_));
 MUX2_X1 _09350_ (.A(_03107_),
    .B(_03108_),
    .S(_01964_),
    .Z(_03109_));
 MUX2_X1 _09351_ (.A(_03106_),
    .B(_03109_),
    .S(_02149_),
    .Z(_03110_));
 AOI221_X1 _09352_ (.A(_01859_),
    .B1(_03100_),
    .B2(_03103_),
    .C1(_03110_),
    .C2(_01887_),
    .ZN(_03111_));
 MUX2_X1 _09353_ (.A(\registers[0][9] ),
    .B(\registers[1][9] ),
    .S(_02043_),
    .Z(_03112_));
 NOR2_X1 _09354_ (.A1(_01866_),
    .A2(_03112_),
    .ZN(_03113_));
 MUX2_X1 _09355_ (.A(\registers[2][9] ),
    .B(\registers[3][9] ),
    .S(_02150_),
    .Z(_03114_));
 NOR3_X1 _09356_ (.A1(_01882_),
    .A2(_01863_),
    .A3(_03114_),
    .ZN(_03115_));
 MUX2_X1 _09357_ (.A(\registers[4][9] ),
    .B(\registers[5][9] ),
    .S(_01955_),
    .Z(_03116_));
 NOR3_X1 _09358_ (.A1(_01888_),
    .A2(_01986_),
    .A3(_03116_),
    .ZN(_03117_));
 MUX2_X1 _09359_ (.A(\registers[6][9] ),
    .B(\registers[7][9] ),
    .S(_01951_),
    .Z(_03118_));
 NOR2_X1 _09360_ (.A1(_01873_),
    .A2(_03118_),
    .ZN(_03119_));
 NOR4_X1 _09361_ (.A1(_03113_),
    .A2(_03115_),
    .A3(_03117_),
    .A4(_03119_),
    .ZN(_03120_));
 MUX2_X1 _09362_ (.A(\registers[12][9] ),
    .B(\registers[14][9] ),
    .S(_02156_),
    .Z(_03121_));
 MUX2_X1 _09363_ (.A(\registers[13][9] ),
    .B(\registers[15][9] ),
    .S(_02158_),
    .Z(_03122_));
 MUX2_X1 _09364_ (.A(_03121_),
    .B(_03122_),
    .S(_02030_),
    .Z(_03123_));
 MUX2_X1 _09365_ (.A(\registers[8][9] ),
    .B(\registers[10][9] ),
    .S(_02162_),
    .Z(_03124_));
 MUX2_X1 _09366_ (.A(\registers[9][9] ),
    .B(\registers[11][9] ),
    .S(_02164_),
    .Z(_03125_));
 MUX2_X1 _09367_ (.A(_03124_),
    .B(_03125_),
    .S(_02160_),
    .Z(_03126_));
 MUX2_X1 _09368_ (.A(_03123_),
    .B(_03126_),
    .S(_01987_),
    .Z(_03127_));
 OAI221_X1 _09369_ (.A(_01909_),
    .B1(_01911_),
    .B2(_03120_),
    .C1(_03127_),
    .C2(_01938_),
    .ZN(_03128_));
 OAI22_X1 _09370_ (.A1(_03094_),
    .A2(_01942_),
    .B1(_03111_),
    .B2(_03128_),
    .ZN(_00360_));
 CLKBUF_X3 _09371_ (.A(read_addr2[4]),
    .Z(_03129_));
 INV_X2 _09372_ (.A(_03129_),
    .ZN(_03130_));
 BUF_X4 _09373_ (.A(_03130_),
    .Z(_03131_));
 BUF_X4 _09374_ (.A(read_addr2[1]),
    .Z(_03132_));
 BUF_X16 _09375_ (.A(_03132_),
    .Z(_03133_));
 BUF_X4 _09376_ (.A(read_addr2[2]),
    .Z(_03134_));
 OR2_X1 _09377_ (.A1(_03133_),
    .A2(_03134_),
    .ZN(_03135_));
 BUF_X4 _09378_ (.A(_03135_),
    .Z(_03136_));
 BUF_X8 _09379_ (.A(_03136_),
    .Z(_03137_));
 BUF_X4 _09380_ (.A(read_addr2[0]),
    .Z(_03138_));
 BUF_X8 _09381_ (.A(_03138_),
    .Z(_03139_));
 BUF_X4 _09382_ (.A(_03139_),
    .Z(_03140_));
 MUX2_X1 _09383_ (.A(\registers[16][0] ),
    .B(\registers[17][0] ),
    .S(_03140_),
    .Z(_03141_));
 BUF_X8 _09384_ (.A(_03132_),
    .Z(_03142_));
 NAND2_X4 _09385_ (.A1(_03142_),
    .A2(_03134_),
    .ZN(_03143_));
 BUF_X4 _09386_ (.A(_03143_),
    .Z(_03144_));
 BUF_X4 _09387_ (.A(_03139_),
    .Z(_03145_));
 MUX2_X1 _09388_ (.A(\registers[22][0] ),
    .B(\registers[23][0] ),
    .S(_03145_),
    .Z(_03146_));
 OAI22_X1 _09389_ (.A1(_03137_),
    .A2(_03141_),
    .B1(_03144_),
    .B2(_03146_),
    .ZN(_03147_));
 BUF_X8 _09390_ (.A(_03138_),
    .Z(_03148_));
 BUF_X4 _09391_ (.A(_03148_),
    .Z(_03149_));
 MUX2_X1 _09392_ (.A(\registers[18][0] ),
    .B(\registers[19][0] ),
    .S(_03149_),
    .Z(_03150_));
 INV_X1 _09393_ (.A(_03150_),
    .ZN(_03151_));
 BUF_X16 _09394_ (.A(_03133_),
    .Z(_03152_));
 INV_X4 _09395_ (.A(_03152_),
    .ZN(_03153_));
 NOR2_X4 _09396_ (.A1(_03153_),
    .A2(_03134_),
    .ZN(_03154_));
 BUF_X4 _09397_ (.A(_03154_),
    .Z(_03155_));
 AOI21_X1 _09398_ (.A(_03147_),
    .B1(_03151_),
    .B2(_03155_),
    .ZN(_03156_));
 BUF_X2 _09399_ (.A(read_addr2[3]),
    .Z(_03157_));
 BUF_X4 _09400_ (.A(_03157_),
    .Z(_03158_));
 BUF_X16 _09401_ (.A(_03152_),
    .Z(_03159_));
 INV_X4 _09402_ (.A(_03134_),
    .ZN(_03160_));
 NOR2_X2 _09403_ (.A1(_03159_),
    .A2(_03160_),
    .ZN(_03161_));
 CLKBUF_X3 _09404_ (.A(_03161_),
    .Z(_03162_));
 BUF_X4 _09405_ (.A(_03139_),
    .Z(_03163_));
 MUX2_X1 _09406_ (.A(\registers[20][0] ),
    .B(\registers[21][0] ),
    .S(_03163_),
    .Z(_03164_));
 INV_X1 _09407_ (.A(_03164_),
    .ZN(_03165_));
 AOI21_X1 _09408_ (.A(_03158_),
    .B1(_03162_),
    .B2(_03165_),
    .ZN(_03166_));
 MUX2_X1 _09409_ (.A(\registers[28][0] ),
    .B(\registers[30][0] ),
    .S(_03152_),
    .Z(_03167_));
 MUX2_X1 _09410_ (.A(\registers[29][0] ),
    .B(\registers[31][0] ),
    .S(_03152_),
    .Z(_03168_));
 BUF_X4 _09411_ (.A(_03138_),
    .Z(_03169_));
 BUF_X4 _09412_ (.A(_03169_),
    .Z(_03170_));
 MUX2_X1 _09413_ (.A(_03167_),
    .B(_03168_),
    .S(_03170_),
    .Z(_03171_));
 MUX2_X1 _09414_ (.A(\registers[24][0] ),
    .B(\registers[26][0] ),
    .S(_03152_),
    .Z(_03172_));
 MUX2_X1 _09415_ (.A(\registers[25][0] ),
    .B(\registers[27][0] ),
    .S(_03152_),
    .Z(_03173_));
 MUX2_X1 _09416_ (.A(_03172_),
    .B(_03173_),
    .S(_03170_),
    .Z(_03174_));
 BUF_X4 _09417_ (.A(_03160_),
    .Z(_03175_));
 MUX2_X1 _09418_ (.A(_03171_),
    .B(_03174_),
    .S(_03175_),
    .Z(_03176_));
 BUF_X4 _09419_ (.A(_03158_),
    .Z(_03177_));
 AOI221_X2 _09420_ (.A(_03131_),
    .B1(_03156_),
    .B2(_03166_),
    .C1(_03176_),
    .C2(_03177_),
    .ZN(_03178_));
 AND2_X1 _09421_ (.A1(_01103_),
    .A2(net2),
    .ZN(_03179_));
 BUF_X2 _09422_ (.A(_03179_),
    .Z(_03180_));
 BUF_X4 _09423_ (.A(_03180_),
    .Z(_03181_));
 OR2_X2 _09424_ (.A1(_03157_),
    .A2(_03129_),
    .ZN(_03182_));
 BUF_X4 _09425_ (.A(_03182_),
    .Z(_03183_));
 BUF_X4 _09426_ (.A(_03137_),
    .Z(_03184_));
 BUF_X4 _09427_ (.A(_03140_),
    .Z(_03185_));
 MUX2_X1 _09428_ (.A(\registers[0][0] ),
    .B(\registers[1][0] ),
    .S(_03185_),
    .Z(_03186_));
 NOR2_X1 _09429_ (.A1(_03184_),
    .A2(_03186_),
    .ZN(_03187_));
 BUF_X4 _09430_ (.A(_03153_),
    .Z(_03188_));
 BUF_X4 _09431_ (.A(_03134_),
    .Z(_03189_));
 BUF_X4 _09432_ (.A(_03148_),
    .Z(_03190_));
 MUX2_X1 _09433_ (.A(\registers[2][0] ),
    .B(\registers[3][0] ),
    .S(_03190_),
    .Z(_03191_));
 NOR3_X1 _09434_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_03191_),
    .ZN(_03192_));
 BUF_X4 _09435_ (.A(_03159_),
    .Z(_03193_));
 BUF_X4 _09436_ (.A(_03139_),
    .Z(_03194_));
 MUX2_X1 _09437_ (.A(\registers[4][0] ),
    .B(\registers[5][0] ),
    .S(_03194_),
    .Z(_03195_));
 NOR3_X1 _09438_ (.A1(_03193_),
    .A2(_03175_),
    .A3(_03195_),
    .ZN(_03196_));
 BUF_X4 _09439_ (.A(_03144_),
    .Z(_03197_));
 MUX2_X1 _09440_ (.A(\registers[6][0] ),
    .B(\registers[7][0] ),
    .S(_03170_),
    .Z(_03198_));
 NOR2_X1 _09441_ (.A1(_03197_),
    .A2(_03198_),
    .ZN(_03199_));
 NOR4_X2 _09442_ (.A1(_03187_),
    .A2(_03192_),
    .A3(_03196_),
    .A4(_03199_),
    .ZN(_03200_));
 MUX2_X1 _09443_ (.A(\registers[12][0] ),
    .B(\registers[14][0] ),
    .S(_03159_),
    .Z(_03201_));
 MUX2_X1 _09444_ (.A(\registers[13][0] ),
    .B(\registers[15][0] ),
    .S(_03159_),
    .Z(_03202_));
 BUF_X4 _09445_ (.A(_03149_),
    .Z(_03203_));
 MUX2_X1 _09446_ (.A(_03201_),
    .B(_03202_),
    .S(_03203_),
    .Z(_03204_));
 MUX2_X1 _09447_ (.A(\registers[8][0] ),
    .B(\registers[10][0] ),
    .S(_03159_),
    .Z(_03205_));
 MUX2_X1 _09448_ (.A(\registers[9][0] ),
    .B(\registers[11][0] ),
    .S(_03159_),
    .Z(_03206_));
 MUX2_X1 _09449_ (.A(_03205_),
    .B(_03206_),
    .S(_03203_),
    .Z(_03207_));
 BUF_X4 _09450_ (.A(_03175_),
    .Z(_03208_));
 MUX2_X1 _09451_ (.A(_03204_),
    .B(_03207_),
    .S(_03208_),
    .Z(_03209_));
 NAND2_X2 _09452_ (.A1(_03158_),
    .A2(_03130_),
    .ZN(_03210_));
 BUF_X4 _09453_ (.A(_03210_),
    .Z(_03211_));
 OAI221_X2 _09454_ (.A(_03181_),
    .B1(_03183_),
    .B2(_03200_),
    .C1(_03209_),
    .C2(_03211_),
    .ZN(_03212_));
 INV_X1 _09455_ (.A(net2),
    .ZN(_03213_));
 NAND2_X2 _09456_ (.A1(_01416_),
    .A2(_03213_),
    .ZN(_03214_));
 INV_X1 _09457_ (.A(net37),
    .ZN(_03215_));
 OAI22_X1 _09458_ (.A1(_03178_),
    .A2(_03212_),
    .B1(_03214_),
    .B2(_03215_),
    .ZN(_00361_));
 INV_X1 _09459_ (.A(net38),
    .ZN(_03216_));
 CLKBUF_X3 _09460_ (.A(_03214_),
    .Z(_03217_));
 BUF_X4 _09461_ (.A(_03129_),
    .Z(_03218_));
 BUF_X4 _09462_ (.A(_03138_),
    .Z(_03219_));
 MUX2_X1 _09463_ (.A(\registers[0][10] ),
    .B(\registers[1][10] ),
    .S(_03219_),
    .Z(_03220_));
 MUX2_X1 _09464_ (.A(\registers[6][10] ),
    .B(\registers[7][10] ),
    .S(_03145_),
    .Z(_03221_));
 OAI22_X1 _09465_ (.A1(_03137_),
    .A2(_03220_),
    .B1(_03221_),
    .B2(_03144_),
    .ZN(_03222_));
 BUF_X4 _09466_ (.A(_03148_),
    .Z(_03223_));
 MUX2_X1 _09467_ (.A(\registers[2][10] ),
    .B(\registers[3][10] ),
    .S(_03223_),
    .Z(_03224_));
 INV_X1 _09468_ (.A(_03224_),
    .ZN(_03225_));
 AOI21_X1 _09469_ (.A(_03222_),
    .B1(_03225_),
    .B2(_03155_),
    .ZN(_03226_));
 BUF_X4 _09470_ (.A(_03139_),
    .Z(_03227_));
 MUX2_X1 _09471_ (.A(\registers[4][10] ),
    .B(\registers[5][10] ),
    .S(_03227_),
    .Z(_03228_));
 INV_X1 _09472_ (.A(_03228_),
    .ZN(_03229_));
 AOI21_X1 _09473_ (.A(_03158_),
    .B1(_03162_),
    .B2(_03229_),
    .ZN(_03230_));
 BUF_X8 _09474_ (.A(_03132_),
    .Z(_03231_));
 BUF_X4 _09475_ (.A(_03231_),
    .Z(_03232_));
 MUX2_X1 _09476_ (.A(\registers[12][10] ),
    .B(\registers[14][10] ),
    .S(_03232_),
    .Z(_03233_));
 BUF_X4 _09477_ (.A(_03231_),
    .Z(_03234_));
 MUX2_X1 _09478_ (.A(\registers[13][10] ),
    .B(\registers[15][10] ),
    .S(_03234_),
    .Z(_03235_));
 BUF_X4 _09479_ (.A(_03148_),
    .Z(_03236_));
 MUX2_X1 _09480_ (.A(_03233_),
    .B(_03235_),
    .S(_03236_),
    .Z(_03237_));
 BUF_X4 _09481_ (.A(_03231_),
    .Z(_03238_));
 MUX2_X1 _09482_ (.A(\registers[8][10] ),
    .B(\registers[10][10] ),
    .S(_03238_),
    .Z(_03239_));
 BUF_X4 _09483_ (.A(_03132_),
    .Z(_03240_));
 MUX2_X1 _09484_ (.A(\registers[9][10] ),
    .B(\registers[11][10] ),
    .S(_03240_),
    .Z(_03241_));
 MUX2_X1 _09485_ (.A(_03239_),
    .B(_03241_),
    .S(_03190_),
    .Z(_03242_));
 MUX2_X2 _09486_ (.A(_03237_),
    .B(_03242_),
    .S(_03175_),
    .Z(_03243_));
 AOI221_X2 _09487_ (.A(_03218_),
    .B1(_03226_),
    .B2(_03230_),
    .C1(_03243_),
    .C2(_03177_),
    .ZN(_03244_));
 NAND2_X1 _09488_ (.A1(_03158_),
    .A2(_03129_),
    .ZN(_03245_));
 CLKBUF_X3 _09489_ (.A(_03245_),
    .Z(_03246_));
 BUF_X8 _09490_ (.A(_03133_),
    .Z(_03247_));
 MUX2_X1 _09491_ (.A(\registers[28][10] ),
    .B(\registers[30][10] ),
    .S(_03247_),
    .Z(_03248_));
 BUF_X8 _09492_ (.A(_03133_),
    .Z(_03249_));
 MUX2_X1 _09493_ (.A(\registers[29][10] ),
    .B(\registers[31][10] ),
    .S(_03249_),
    .Z(_03250_));
 BUF_X4 _09494_ (.A(_03140_),
    .Z(_03251_));
 MUX2_X1 _09495_ (.A(_03248_),
    .B(_03250_),
    .S(_03251_),
    .Z(_03252_));
 BUF_X8 _09496_ (.A(_03133_),
    .Z(_03253_));
 MUX2_X1 _09497_ (.A(\registers[24][10] ),
    .B(\registers[26][10] ),
    .S(_03253_),
    .Z(_03254_));
 BUF_X4 _09498_ (.A(_03142_),
    .Z(_03255_));
 MUX2_X1 _09499_ (.A(\registers[25][10] ),
    .B(\registers[27][10] ),
    .S(_03255_),
    .Z(_03256_));
 MUX2_X1 _09500_ (.A(_03254_),
    .B(_03256_),
    .S(_03185_),
    .Z(_03257_));
 BUF_X4 _09501_ (.A(_03160_),
    .Z(_03258_));
 BUF_X4 _09502_ (.A(_03258_),
    .Z(_03259_));
 MUX2_X1 _09503_ (.A(_03252_),
    .B(_03257_),
    .S(_03259_),
    .Z(_03260_));
 CLKBUF_X3 _09504_ (.A(_03157_),
    .Z(_03261_));
 OR2_X1 _09505_ (.A1(_03261_),
    .A2(_03130_),
    .ZN(_03262_));
 CLKBUF_X3 _09506_ (.A(_03262_),
    .Z(_03263_));
 BUF_X4 _09507_ (.A(_03137_),
    .Z(_03264_));
 MUX2_X1 _09508_ (.A(\registers[16][10] ),
    .B(\registers[17][10] ),
    .S(_03185_),
    .Z(_03265_));
 NOR2_X1 _09509_ (.A1(_03264_),
    .A2(_03265_),
    .ZN(_03266_));
 BUF_X4 _09510_ (.A(_03153_),
    .Z(_03267_));
 BUF_X4 _09511_ (.A(_03134_),
    .Z(_03268_));
 MUX2_X1 _09512_ (.A(\registers[18][10] ),
    .B(\registers[19][10] ),
    .S(_03170_),
    .Z(_03269_));
 NOR3_X2 _09513_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_03269_),
    .ZN(_03270_));
 BUF_X4 _09514_ (.A(_03159_),
    .Z(_03271_));
 BUF_X4 _09515_ (.A(_03148_),
    .Z(_03272_));
 MUX2_X1 _09516_ (.A(\registers[20][10] ),
    .B(\registers[21][10] ),
    .S(_03272_),
    .Z(_03273_));
 NOR3_X1 _09517_ (.A1(_03271_),
    .A2(_03175_),
    .A3(_03273_),
    .ZN(_03274_));
 BUF_X4 _09518_ (.A(_03144_),
    .Z(_03275_));
 MUX2_X1 _09519_ (.A(\registers[22][10] ),
    .B(\registers[23][10] ),
    .S(_03170_),
    .Z(_03276_));
 NOR2_X1 _09520_ (.A1(_03275_),
    .A2(_03276_),
    .ZN(_03277_));
 NOR4_X2 _09521_ (.A1(_03266_),
    .A2(_03270_),
    .A3(_03274_),
    .A4(_03277_),
    .ZN(_03278_));
 OAI221_X1 _09522_ (.A(_03181_),
    .B1(_03246_),
    .B2(_03260_),
    .C1(_03263_),
    .C2(_03278_),
    .ZN(_03279_));
 OAI22_X1 _09523_ (.A1(_03216_),
    .A2(_03217_),
    .B1(_03244_),
    .B2(_03279_),
    .ZN(_00362_));
 INV_X1 _09524_ (.A(net39),
    .ZN(_03280_));
 MUX2_X1 _09525_ (.A(\registers[0][11] ),
    .B(\registers[1][11] ),
    .S(_03219_),
    .Z(_03281_));
 MUX2_X1 _09526_ (.A(\registers[6][11] ),
    .B(\registers[7][11] ),
    .S(_03145_),
    .Z(_03282_));
 OAI22_X1 _09527_ (.A1(_03137_),
    .A2(_03281_),
    .B1(_03282_),
    .B2(_03144_),
    .ZN(_03283_));
 MUX2_X1 _09528_ (.A(\registers[2][11] ),
    .B(\registers[3][11] ),
    .S(_03223_),
    .Z(_03284_));
 INV_X1 _09529_ (.A(_03284_),
    .ZN(_03285_));
 AOI21_X1 _09530_ (.A(_03283_),
    .B1(_03285_),
    .B2(_03155_),
    .ZN(_03286_));
 MUX2_X1 _09531_ (.A(\registers[4][11] ),
    .B(\registers[5][11] ),
    .S(_03227_),
    .Z(_03287_));
 INV_X1 _09532_ (.A(_03287_),
    .ZN(_03288_));
 AOI21_X1 _09533_ (.A(_03158_),
    .B1(_03162_),
    .B2(_03288_),
    .ZN(_03289_));
 MUX2_X1 _09534_ (.A(\registers[12][11] ),
    .B(\registers[14][11] ),
    .S(_03232_),
    .Z(_03290_));
 MUX2_X1 _09535_ (.A(\registers[13][11] ),
    .B(\registers[15][11] ),
    .S(_03234_),
    .Z(_03291_));
 MUX2_X1 _09536_ (.A(_03290_),
    .B(_03291_),
    .S(_03236_),
    .Z(_03292_));
 MUX2_X1 _09537_ (.A(\registers[8][11] ),
    .B(\registers[10][11] ),
    .S(_03238_),
    .Z(_03293_));
 MUX2_X1 _09538_ (.A(\registers[9][11] ),
    .B(\registers[11][11] ),
    .S(_03240_),
    .Z(_03294_));
 MUX2_X1 _09539_ (.A(_03293_),
    .B(_03294_),
    .S(_03190_),
    .Z(_03295_));
 MUX2_X2 _09540_ (.A(_03292_),
    .B(_03295_),
    .S(_03175_),
    .Z(_03296_));
 AOI221_X2 _09541_ (.A(_03218_),
    .B1(_03286_),
    .B2(_03289_),
    .C1(_03296_),
    .C2(_03177_),
    .ZN(_03297_));
 MUX2_X1 _09542_ (.A(\registers[28][11] ),
    .B(\registers[30][11] ),
    .S(_03247_),
    .Z(_03298_));
 MUX2_X1 _09543_ (.A(\registers[29][11] ),
    .B(\registers[31][11] ),
    .S(_03249_),
    .Z(_03299_));
 MUX2_X1 _09544_ (.A(_03298_),
    .B(_03299_),
    .S(_03251_),
    .Z(_03300_));
 MUX2_X1 _09545_ (.A(\registers[24][11] ),
    .B(\registers[26][11] ),
    .S(_03253_),
    .Z(_03301_));
 MUX2_X1 _09546_ (.A(\registers[25][11] ),
    .B(\registers[27][11] ),
    .S(_03255_),
    .Z(_03302_));
 MUX2_X1 _09547_ (.A(_03301_),
    .B(_03302_),
    .S(_03185_),
    .Z(_03303_));
 MUX2_X1 _09548_ (.A(_03300_),
    .B(_03303_),
    .S(_03259_),
    .Z(_03304_));
 BUF_X4 _09549_ (.A(_03137_),
    .Z(_03305_));
 BUF_X4 _09550_ (.A(_03194_),
    .Z(_03306_));
 MUX2_X1 _09551_ (.A(\registers[16][11] ),
    .B(\registers[17][11] ),
    .S(_03306_),
    .Z(_03307_));
 NOR2_X1 _09552_ (.A1(_03305_),
    .A2(_03307_),
    .ZN(_03308_));
 CLKBUF_X3 _09553_ (.A(_03153_),
    .Z(_03309_));
 CLKBUF_X3 _09554_ (.A(_03134_),
    .Z(_03310_));
 BUF_X4 _09555_ (.A(_03219_),
    .Z(_03311_));
 MUX2_X1 _09556_ (.A(\registers[18][11] ),
    .B(\registers[19][11] ),
    .S(_03311_),
    .Z(_03312_));
 NOR3_X1 _09557_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03312_),
    .ZN(_03313_));
 CLKBUF_X3 _09558_ (.A(_03159_),
    .Z(_03314_));
 BUF_X4 _09559_ (.A(_03160_),
    .Z(_03315_));
 MUX2_X1 _09560_ (.A(\registers[20][11] ),
    .B(\registers[21][11] ),
    .S(_03170_),
    .Z(_03316_));
 NOR3_X1 _09561_ (.A1(_03314_),
    .A2(_03315_),
    .A3(_03316_),
    .ZN(_03317_));
 BUF_X4 _09562_ (.A(_03144_),
    .Z(_03318_));
 BUF_X4 _09563_ (.A(_03219_),
    .Z(_03319_));
 MUX2_X1 _09564_ (.A(\registers[22][11] ),
    .B(\registers[23][11] ),
    .S(_03319_),
    .Z(_03320_));
 NOR2_X1 _09565_ (.A1(_03318_),
    .A2(_03320_),
    .ZN(_03321_));
 NOR4_X1 _09566_ (.A1(_03308_),
    .A2(_03313_),
    .A3(_03317_),
    .A4(_03321_),
    .ZN(_03322_));
 OAI221_X1 _09567_ (.A(_03181_),
    .B1(_03246_),
    .B2(_03304_),
    .C1(_03322_),
    .C2(_03263_),
    .ZN(_03323_));
 OAI22_X1 _09568_ (.A1(_03280_),
    .A2(_03217_),
    .B1(_03297_),
    .B2(_03323_),
    .ZN(_00363_));
 INV_X1 _09569_ (.A(net40),
    .ZN(_03324_));
 MUX2_X1 _09570_ (.A(\registers[0][12] ),
    .B(\registers[1][12] ),
    .S(_03219_),
    .Z(_03325_));
 MUX2_X1 _09571_ (.A(\registers[6][12] ),
    .B(\registers[7][12] ),
    .S(_03145_),
    .Z(_03326_));
 OAI22_X1 _09572_ (.A1(_03137_),
    .A2(_03325_),
    .B1(_03326_),
    .B2(_03144_),
    .ZN(_03327_));
 MUX2_X1 _09573_ (.A(\registers[2][12] ),
    .B(\registers[3][12] ),
    .S(_03223_),
    .Z(_03328_));
 INV_X1 _09574_ (.A(_03328_),
    .ZN(_03329_));
 AOI21_X1 _09575_ (.A(_03327_),
    .B1(_03329_),
    .B2(_03155_),
    .ZN(_03330_));
 CLKBUF_X3 _09576_ (.A(_03157_),
    .Z(_03331_));
 MUX2_X1 _09577_ (.A(\registers[4][12] ),
    .B(\registers[5][12] ),
    .S(_03227_),
    .Z(_03332_));
 INV_X1 _09578_ (.A(_03332_),
    .ZN(_03333_));
 AOI21_X1 _09579_ (.A(_03331_),
    .B1(_03162_),
    .B2(_03333_),
    .ZN(_03334_));
 MUX2_X1 _09580_ (.A(\registers[12][12] ),
    .B(\registers[14][12] ),
    .S(_03232_),
    .Z(_03335_));
 MUX2_X1 _09581_ (.A(\registers[13][12] ),
    .B(\registers[15][12] ),
    .S(_03234_),
    .Z(_03336_));
 MUX2_X1 _09582_ (.A(_03335_),
    .B(_03336_),
    .S(_03236_),
    .Z(_03337_));
 MUX2_X1 _09583_ (.A(\registers[8][12] ),
    .B(\registers[10][12] ),
    .S(_03238_),
    .Z(_03338_));
 MUX2_X1 _09584_ (.A(\registers[9][12] ),
    .B(\registers[11][12] ),
    .S(_03240_),
    .Z(_03339_));
 MUX2_X1 _09585_ (.A(_03338_),
    .B(_03339_),
    .S(_03190_),
    .Z(_03340_));
 MUX2_X2 _09586_ (.A(_03337_),
    .B(_03340_),
    .S(_03175_),
    .Z(_03341_));
 AOI221_X2 _09587_ (.A(_03218_),
    .B1(_03330_),
    .B2(_03334_),
    .C1(_03341_),
    .C2(_03177_),
    .ZN(_03342_));
 MUX2_X1 _09588_ (.A(\registers[28][12] ),
    .B(\registers[30][12] ),
    .S(_03247_),
    .Z(_03343_));
 MUX2_X1 _09589_ (.A(\registers[29][12] ),
    .B(\registers[31][12] ),
    .S(_03249_),
    .Z(_03344_));
 MUX2_X1 _09590_ (.A(_03343_),
    .B(_03344_),
    .S(_03251_),
    .Z(_03345_));
 MUX2_X1 _09591_ (.A(\registers[24][12] ),
    .B(\registers[26][12] ),
    .S(_03253_),
    .Z(_03346_));
 MUX2_X1 _09592_ (.A(\registers[25][12] ),
    .B(\registers[27][12] ),
    .S(_03255_),
    .Z(_03347_));
 MUX2_X1 _09593_ (.A(_03346_),
    .B(_03347_),
    .S(_03185_),
    .Z(_03348_));
 MUX2_X1 _09594_ (.A(_03345_),
    .B(_03348_),
    .S(_03259_),
    .Z(_03349_));
 MUX2_X1 _09595_ (.A(\registers[16][12] ),
    .B(\registers[17][12] ),
    .S(_03306_),
    .Z(_03350_));
 NOR2_X1 _09596_ (.A1(_03305_),
    .A2(_03350_),
    .ZN(_03351_));
 MUX2_X1 _09597_ (.A(\registers[18][12] ),
    .B(\registers[19][12] ),
    .S(_03311_),
    .Z(_03352_));
 NOR3_X1 _09598_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03352_),
    .ZN(_03353_));
 BUF_X4 _09599_ (.A(_03169_),
    .Z(_03354_));
 MUX2_X1 _09600_ (.A(\registers[20][12] ),
    .B(\registers[21][12] ),
    .S(_03354_),
    .Z(_03355_));
 NOR3_X1 _09601_ (.A1(_03314_),
    .A2(_03315_),
    .A3(_03355_),
    .ZN(_03356_));
 MUX2_X1 _09602_ (.A(\registers[22][12] ),
    .B(\registers[23][12] ),
    .S(_03319_),
    .Z(_03357_));
 NOR2_X1 _09603_ (.A1(_03318_),
    .A2(_03357_),
    .ZN(_03358_));
 NOR4_X1 _09604_ (.A1(_03351_),
    .A2(_03353_),
    .A3(_03356_),
    .A4(_03358_),
    .ZN(_03359_));
 OAI221_X1 _09605_ (.A(_03181_),
    .B1(_03246_),
    .B2(_03349_),
    .C1(_03359_),
    .C2(_03263_),
    .ZN(_03360_));
 OAI22_X1 _09606_ (.A1(_03324_),
    .A2(_03217_),
    .B1(_03342_),
    .B2(_03360_),
    .ZN(_00364_));
 INV_X1 _09607_ (.A(net41),
    .ZN(_03361_));
 MUX2_X1 _09608_ (.A(\registers[16][13] ),
    .B(\registers[17][13] ),
    .S(_03219_),
    .Z(_03362_));
 MUX2_X1 _09609_ (.A(\registers[22][13] ),
    .B(\registers[23][13] ),
    .S(_03145_),
    .Z(_03363_));
 OAI22_X1 _09610_ (.A1(_03137_),
    .A2(_03362_),
    .B1(_03363_),
    .B2(_03144_),
    .ZN(_03364_));
 MUX2_X1 _09611_ (.A(\registers[18][13] ),
    .B(\registers[19][13] ),
    .S(_03223_),
    .Z(_03365_));
 INV_X1 _09612_ (.A(_03365_),
    .ZN(_03366_));
 AOI21_X1 _09613_ (.A(_03364_),
    .B1(_03366_),
    .B2(_03155_),
    .ZN(_03367_));
 MUX2_X1 _09614_ (.A(\registers[20][13] ),
    .B(\registers[21][13] ),
    .S(_03227_),
    .Z(_03368_));
 INV_X1 _09615_ (.A(_03368_),
    .ZN(_03369_));
 AOI21_X1 _09616_ (.A(_03331_),
    .B1(_03162_),
    .B2(_03369_),
    .ZN(_03370_));
 BUF_X4 _09617_ (.A(_03231_),
    .Z(_03371_));
 MUX2_X1 _09618_ (.A(\registers[28][13] ),
    .B(\registers[30][13] ),
    .S(_03371_),
    .Z(_03372_));
 MUX2_X1 _09619_ (.A(\registers[29][13] ),
    .B(\registers[31][13] ),
    .S(_03234_),
    .Z(_03373_));
 MUX2_X1 _09620_ (.A(_03372_),
    .B(_03373_),
    .S(_03236_),
    .Z(_03374_));
 MUX2_X1 _09621_ (.A(\registers[24][13] ),
    .B(\registers[26][13] ),
    .S(_03238_),
    .Z(_03375_));
 MUX2_X1 _09622_ (.A(\registers[25][13] ),
    .B(\registers[27][13] ),
    .S(_03240_),
    .Z(_03376_));
 MUX2_X1 _09623_ (.A(_03375_),
    .B(_03376_),
    .S(_03190_),
    .Z(_03377_));
 MUX2_X1 _09624_ (.A(_03374_),
    .B(_03377_),
    .S(_03175_),
    .Z(_03378_));
 AOI221_X2 _09625_ (.A(_03131_),
    .B1(_03367_),
    .B2(_03370_),
    .C1(_03378_),
    .C2(_03177_),
    .ZN(_03379_));
 BUF_X4 _09626_ (.A(_03140_),
    .Z(_03380_));
 MUX2_X1 _09627_ (.A(\registers[0][13] ),
    .B(\registers[1][13] ),
    .S(_03380_),
    .Z(_03381_));
 NOR2_X1 _09628_ (.A1(_03184_),
    .A2(_03381_),
    .ZN(_03382_));
 MUX2_X1 _09629_ (.A(\registers[2][13] ),
    .B(\registers[3][13] ),
    .S(_03163_),
    .Z(_03383_));
 NOR3_X1 _09630_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_03383_),
    .ZN(_03384_));
 BUF_X4 _09631_ (.A(_03160_),
    .Z(_03385_));
 BUF_X4 _09632_ (.A(_03139_),
    .Z(_03386_));
 MUX2_X1 _09633_ (.A(\registers[4][13] ),
    .B(\registers[5][13] ),
    .S(_03386_),
    .Z(_03387_));
 NOR3_X1 _09634_ (.A1(_03193_),
    .A2(_03385_),
    .A3(_03387_),
    .ZN(_03388_));
 MUX2_X1 _09635_ (.A(\registers[6][13] ),
    .B(\registers[7][13] ),
    .S(_03272_),
    .Z(_03389_));
 NOR2_X1 _09636_ (.A1(_03197_),
    .A2(_03389_),
    .ZN(_03390_));
 NOR4_X2 _09637_ (.A1(_03382_),
    .A2(_03384_),
    .A3(_03388_),
    .A4(_03390_),
    .ZN(_03391_));
 BUF_X4 _09638_ (.A(_03240_),
    .Z(_03392_));
 MUX2_X1 _09639_ (.A(\registers[12][13] ),
    .B(\registers[14][13] ),
    .S(_03392_),
    .Z(_03393_));
 BUF_X4 _09640_ (.A(_03240_),
    .Z(_03394_));
 MUX2_X1 _09641_ (.A(\registers[13][13] ),
    .B(\registers[15][13] ),
    .S(_03394_),
    .Z(_03395_));
 BUF_X4 _09642_ (.A(_03190_),
    .Z(_03396_));
 MUX2_X1 _09643_ (.A(_03393_),
    .B(_03395_),
    .S(_03396_),
    .Z(_03397_));
 BUF_X4 _09644_ (.A(_03240_),
    .Z(_03398_));
 MUX2_X1 _09645_ (.A(\registers[8][13] ),
    .B(\registers[10][13] ),
    .S(_03398_),
    .Z(_03399_));
 BUF_X4 _09646_ (.A(_03240_),
    .Z(_03400_));
 MUX2_X1 _09647_ (.A(\registers[9][13] ),
    .B(\registers[11][13] ),
    .S(_03400_),
    .Z(_03401_));
 MUX2_X1 _09648_ (.A(_03399_),
    .B(_03401_),
    .S(_03203_),
    .Z(_03402_));
 MUX2_X2 _09649_ (.A(_03397_),
    .B(_03402_),
    .S(_03208_),
    .Z(_03403_));
 OAI221_X2 _09650_ (.A(_03181_),
    .B1(_03183_),
    .B2(_03391_),
    .C1(_03403_),
    .C2(_03211_),
    .ZN(_03404_));
 OAI22_X1 _09651_ (.A1(_03361_),
    .A2(_03217_),
    .B1(_03379_),
    .B2(_03404_),
    .ZN(_00365_));
 INV_X1 _09652_ (.A(net42),
    .ZN(_03405_));
 BUF_X4 _09653_ (.A(_03136_),
    .Z(_03406_));
 MUX2_X1 _09654_ (.A(\registers[0][14] ),
    .B(\registers[1][14] ),
    .S(_03219_),
    .Z(_03407_));
 BUF_X4 _09655_ (.A(_03138_),
    .Z(_03408_));
 MUX2_X1 _09656_ (.A(\registers[6][14] ),
    .B(\registers[7][14] ),
    .S(_03408_),
    .Z(_03409_));
 BUF_X4 _09657_ (.A(_03143_),
    .Z(_03410_));
 OAI22_X1 _09658_ (.A1(_03406_),
    .A2(_03407_),
    .B1(_03409_),
    .B2(_03410_),
    .ZN(_03411_));
 BUF_X4 _09659_ (.A(_03148_),
    .Z(_03412_));
 MUX2_X1 _09660_ (.A(\registers[2][14] ),
    .B(\registers[3][14] ),
    .S(_03412_),
    .Z(_03413_));
 INV_X1 _09661_ (.A(_03413_),
    .ZN(_03414_));
 AOI21_X1 _09662_ (.A(_03411_),
    .B1(_03414_),
    .B2(_03155_),
    .ZN(_03415_));
 MUX2_X1 _09663_ (.A(\registers[4][14] ),
    .B(\registers[5][14] ),
    .S(_03227_),
    .Z(_03416_));
 INV_X1 _09664_ (.A(_03416_),
    .ZN(_03417_));
 AOI21_X1 _09665_ (.A(_03331_),
    .B1(_03162_),
    .B2(_03417_),
    .ZN(_03418_));
 MUX2_X1 _09666_ (.A(\registers[12][14] ),
    .B(\registers[14][14] ),
    .S(_03371_),
    .Z(_03419_));
 BUF_X4 _09667_ (.A(_03231_),
    .Z(_03420_));
 MUX2_X1 _09668_ (.A(\registers[13][14] ),
    .B(\registers[15][14] ),
    .S(_03420_),
    .Z(_03421_));
 MUX2_X1 _09669_ (.A(_03419_),
    .B(_03421_),
    .S(_03236_),
    .Z(_03422_));
 MUX2_X1 _09670_ (.A(\registers[8][14] ),
    .B(\registers[10][14] ),
    .S(_03238_),
    .Z(_03423_));
 MUX2_X1 _09671_ (.A(\registers[9][14] ),
    .B(\registers[11][14] ),
    .S(_03240_),
    .Z(_03424_));
 MUX2_X1 _09672_ (.A(_03423_),
    .B(_03424_),
    .S(_03190_),
    .Z(_03425_));
 MUX2_X2 _09673_ (.A(_03422_),
    .B(_03425_),
    .S(_03175_),
    .Z(_03426_));
 AOI221_X1 _09674_ (.A(_03218_),
    .B1(_03415_),
    .B2(_03418_),
    .C1(_03426_),
    .C2(_03177_),
    .ZN(_03427_));
 MUX2_X1 _09675_ (.A(\registers[28][14] ),
    .B(\registers[30][14] ),
    .S(_03247_),
    .Z(_03428_));
 MUX2_X1 _09676_ (.A(\registers[29][14] ),
    .B(\registers[31][14] ),
    .S(_03249_),
    .Z(_03429_));
 MUX2_X1 _09677_ (.A(_03428_),
    .B(_03429_),
    .S(_03251_),
    .Z(_03430_));
 MUX2_X1 _09678_ (.A(\registers[24][14] ),
    .B(\registers[26][14] ),
    .S(_03253_),
    .Z(_03431_));
 MUX2_X1 _09679_ (.A(\registers[25][14] ),
    .B(\registers[27][14] ),
    .S(_03255_),
    .Z(_03432_));
 MUX2_X1 _09680_ (.A(_03431_),
    .B(_03432_),
    .S(_03185_),
    .Z(_03433_));
 MUX2_X1 _09681_ (.A(_03430_),
    .B(_03433_),
    .S(_03259_),
    .Z(_03434_));
 MUX2_X1 _09682_ (.A(\registers[16][14] ),
    .B(\registers[17][14] ),
    .S(_03306_),
    .Z(_03435_));
 NOR2_X1 _09683_ (.A1(_03305_),
    .A2(_03435_),
    .ZN(_03436_));
 MUX2_X1 _09684_ (.A(\registers[18][14] ),
    .B(\registers[19][14] ),
    .S(_03311_),
    .Z(_03437_));
 NOR3_X1 _09685_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03437_),
    .ZN(_03438_));
 MUX2_X1 _09686_ (.A(\registers[20][14] ),
    .B(\registers[21][14] ),
    .S(_03354_),
    .Z(_03439_));
 NOR3_X1 _09687_ (.A1(_03314_),
    .A2(_03315_),
    .A3(_03439_),
    .ZN(_03440_));
 MUX2_X1 _09688_ (.A(\registers[22][14] ),
    .B(\registers[23][14] ),
    .S(_03319_),
    .Z(_03441_));
 NOR2_X1 _09689_ (.A1(_03318_),
    .A2(_03441_),
    .ZN(_03442_));
 NOR4_X1 _09690_ (.A1(_03436_),
    .A2(_03438_),
    .A3(_03440_),
    .A4(_03442_),
    .ZN(_03443_));
 OAI221_X1 _09691_ (.A(_03181_),
    .B1(_03246_),
    .B2(_03434_),
    .C1(_03443_),
    .C2(_03263_),
    .ZN(_03444_));
 OAI22_X1 _09692_ (.A1(_03405_),
    .A2(_03217_),
    .B1(_03427_),
    .B2(_03444_),
    .ZN(_00366_));
 INV_X1 _09693_ (.A(net43),
    .ZN(_03445_));
 MUX2_X1 _09694_ (.A(\registers[0][15] ),
    .B(\registers[1][15] ),
    .S(_03219_),
    .Z(_03446_));
 MUX2_X1 _09695_ (.A(\registers[6][15] ),
    .B(\registers[7][15] ),
    .S(_03408_),
    .Z(_03447_));
 OAI22_X1 _09696_ (.A1(_03406_),
    .A2(_03446_),
    .B1(_03447_),
    .B2(_03410_),
    .ZN(_03448_));
 MUX2_X1 _09697_ (.A(\registers[2][15] ),
    .B(\registers[3][15] ),
    .S(_03412_),
    .Z(_03449_));
 INV_X1 _09698_ (.A(_03449_),
    .ZN(_03450_));
 AOI21_X1 _09699_ (.A(_03448_),
    .B1(_03450_),
    .B2(_03155_),
    .ZN(_03451_));
 MUX2_X1 _09700_ (.A(\registers[4][15] ),
    .B(\registers[5][15] ),
    .S(_03227_),
    .Z(_03452_));
 INV_X1 _09701_ (.A(_03452_),
    .ZN(_03453_));
 AOI21_X1 _09702_ (.A(_03331_),
    .B1(_03162_),
    .B2(_03453_),
    .ZN(_03454_));
 MUX2_X1 _09703_ (.A(\registers[12][15] ),
    .B(\registers[14][15] ),
    .S(_03371_),
    .Z(_03455_));
 MUX2_X1 _09704_ (.A(\registers[13][15] ),
    .B(\registers[15][15] ),
    .S(_03420_),
    .Z(_03456_));
 MUX2_X1 _09705_ (.A(_03455_),
    .B(_03456_),
    .S(_03236_),
    .Z(_03457_));
 BUF_X4 _09706_ (.A(_03231_),
    .Z(_03458_));
 MUX2_X1 _09707_ (.A(\registers[8][15] ),
    .B(\registers[10][15] ),
    .S(_03458_),
    .Z(_03459_));
 MUX2_X1 _09708_ (.A(\registers[9][15] ),
    .B(\registers[11][15] ),
    .S(_03240_),
    .Z(_03460_));
 MUX2_X1 _09709_ (.A(_03459_),
    .B(_03460_),
    .S(_03190_),
    .Z(_03461_));
 BUF_X4 _09710_ (.A(_03160_),
    .Z(_03462_));
 MUX2_X2 _09711_ (.A(_03457_),
    .B(_03461_),
    .S(_03462_),
    .Z(_03463_));
 AOI221_X2 _09712_ (.A(_03218_),
    .B1(_03451_),
    .B2(_03454_),
    .C1(_03463_),
    .C2(_03177_),
    .ZN(_03464_));
 MUX2_X1 _09713_ (.A(\registers[28][15] ),
    .B(\registers[30][15] ),
    .S(_03247_),
    .Z(_03465_));
 MUX2_X1 _09714_ (.A(\registers[29][15] ),
    .B(\registers[31][15] ),
    .S(_03249_),
    .Z(_03466_));
 MUX2_X1 _09715_ (.A(_03465_),
    .B(_03466_),
    .S(_03251_),
    .Z(_03467_));
 MUX2_X1 _09716_ (.A(\registers[24][15] ),
    .B(\registers[26][15] ),
    .S(_03253_),
    .Z(_03468_));
 MUX2_X1 _09717_ (.A(\registers[25][15] ),
    .B(\registers[27][15] ),
    .S(_03255_),
    .Z(_03469_));
 MUX2_X1 _09718_ (.A(_03468_),
    .B(_03469_),
    .S(_03185_),
    .Z(_03470_));
 MUX2_X1 _09719_ (.A(_03467_),
    .B(_03470_),
    .S(_03259_),
    .Z(_03471_));
 MUX2_X1 _09720_ (.A(\registers[16][15] ),
    .B(\registers[17][15] ),
    .S(_03306_),
    .Z(_03472_));
 NOR2_X1 _09721_ (.A1(_03305_),
    .A2(_03472_),
    .ZN(_03473_));
 MUX2_X1 _09722_ (.A(\registers[18][15] ),
    .B(\registers[19][15] ),
    .S(_03311_),
    .Z(_03474_));
 NOR3_X1 _09723_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03474_),
    .ZN(_03475_));
 MUX2_X1 _09724_ (.A(\registers[20][15] ),
    .B(\registers[21][15] ),
    .S(_03354_),
    .Z(_03476_));
 NOR3_X1 _09725_ (.A1(_03314_),
    .A2(_03315_),
    .A3(_03476_),
    .ZN(_03477_));
 MUX2_X1 _09726_ (.A(\registers[22][15] ),
    .B(\registers[23][15] ),
    .S(_03319_),
    .Z(_03478_));
 NOR2_X1 _09727_ (.A1(_03318_),
    .A2(_03478_),
    .ZN(_03479_));
 NOR4_X2 _09728_ (.A1(_03473_),
    .A2(_03475_),
    .A3(_03477_),
    .A4(_03479_),
    .ZN(_03480_));
 OAI221_X1 _09729_ (.A(_03181_),
    .B1(_03246_),
    .B2(_03471_),
    .C1(_03480_),
    .C2(_03263_),
    .ZN(_03481_));
 OAI22_X1 _09730_ (.A1(_03445_),
    .A2(_03217_),
    .B1(_03464_),
    .B2(_03481_),
    .ZN(_00367_));
 INV_X1 _09731_ (.A(net44),
    .ZN(_03482_));
 BUF_X4 _09732_ (.A(_03139_),
    .Z(_03483_));
 MUX2_X1 _09733_ (.A(\registers[0][16] ),
    .B(\registers[1][16] ),
    .S(_03483_),
    .Z(_03484_));
 MUX2_X1 _09734_ (.A(\registers[6][16] ),
    .B(\registers[7][16] ),
    .S(_03408_),
    .Z(_03485_));
 OAI22_X1 _09735_ (.A1(_03406_),
    .A2(_03484_),
    .B1(_03485_),
    .B2(_03410_),
    .ZN(_03486_));
 MUX2_X1 _09736_ (.A(\registers[2][16] ),
    .B(\registers[3][16] ),
    .S(_03412_),
    .Z(_03487_));
 INV_X1 _09737_ (.A(_03487_),
    .ZN(_03488_));
 AOI21_X1 _09738_ (.A(_03486_),
    .B1(_03488_),
    .B2(_03155_),
    .ZN(_03489_));
 MUX2_X1 _09739_ (.A(\registers[4][16] ),
    .B(\registers[5][16] ),
    .S(_03227_),
    .Z(_03490_));
 INV_X1 _09740_ (.A(_03490_),
    .ZN(_03491_));
 AOI21_X1 _09741_ (.A(_03331_),
    .B1(_03162_),
    .B2(_03491_),
    .ZN(_03492_));
 MUX2_X1 _09742_ (.A(\registers[12][16] ),
    .B(\registers[14][16] ),
    .S(_03371_),
    .Z(_03493_));
 MUX2_X1 _09743_ (.A(\registers[13][16] ),
    .B(\registers[15][16] ),
    .S(_03420_),
    .Z(_03494_));
 MUX2_X1 _09744_ (.A(_03493_),
    .B(_03494_),
    .S(_03236_),
    .Z(_03495_));
 MUX2_X1 _09745_ (.A(\registers[8][16] ),
    .B(\registers[10][16] ),
    .S(_03458_),
    .Z(_03496_));
 BUF_X4 _09746_ (.A(_03133_),
    .Z(_03497_));
 MUX2_X1 _09747_ (.A(\registers[9][16] ),
    .B(\registers[11][16] ),
    .S(_03497_),
    .Z(_03498_));
 MUX2_X1 _09748_ (.A(_03496_),
    .B(_03498_),
    .S(_03190_),
    .Z(_03499_));
 MUX2_X2 _09749_ (.A(_03495_),
    .B(_03499_),
    .S(_03462_),
    .Z(_03500_));
 AOI221_X2 _09750_ (.A(_03218_),
    .B1(_03489_),
    .B2(_03492_),
    .C1(_03500_),
    .C2(_03177_),
    .ZN(_03501_));
 MUX2_X1 _09751_ (.A(\registers[28][16] ),
    .B(\registers[30][16] ),
    .S(_03247_),
    .Z(_03502_));
 MUX2_X1 _09752_ (.A(\registers[29][16] ),
    .B(\registers[31][16] ),
    .S(_03249_),
    .Z(_03503_));
 BUF_X4 _09753_ (.A(_03140_),
    .Z(_03504_));
 MUX2_X1 _09754_ (.A(_03502_),
    .B(_03503_),
    .S(_03504_),
    .Z(_03505_));
 MUX2_X1 _09755_ (.A(\registers[24][16] ),
    .B(\registers[26][16] ),
    .S(_03253_),
    .Z(_03506_));
 MUX2_X1 _09756_ (.A(\registers[25][16] ),
    .B(\registers[27][16] ),
    .S(_03255_),
    .Z(_03507_));
 BUF_X4 _09757_ (.A(_03140_),
    .Z(_03508_));
 MUX2_X1 _09758_ (.A(_03506_),
    .B(_03507_),
    .S(_03508_),
    .Z(_03509_));
 MUX2_X1 _09759_ (.A(_03505_),
    .B(_03509_),
    .S(_03259_),
    .Z(_03510_));
 MUX2_X1 _09760_ (.A(\registers[16][16] ),
    .B(\registers[17][16] ),
    .S(_03306_),
    .Z(_03511_));
 NOR2_X1 _09761_ (.A1(_03305_),
    .A2(_03511_),
    .ZN(_03512_));
 MUX2_X1 _09762_ (.A(\registers[18][16] ),
    .B(\registers[19][16] ),
    .S(_03311_),
    .Z(_03513_));
 NOR3_X1 _09763_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03513_),
    .ZN(_03514_));
 MUX2_X1 _09764_ (.A(\registers[20][16] ),
    .B(\registers[21][16] ),
    .S(_03354_),
    .Z(_03515_));
 NOR3_X1 _09765_ (.A1(_03314_),
    .A2(_03315_),
    .A3(_03515_),
    .ZN(_03516_));
 BUF_X4 _09766_ (.A(_03219_),
    .Z(_03517_));
 MUX2_X1 _09767_ (.A(\registers[22][16] ),
    .B(\registers[23][16] ),
    .S(_03517_),
    .Z(_03518_));
 NOR2_X1 _09768_ (.A1(_03318_),
    .A2(_03518_),
    .ZN(_03519_));
 NOR4_X1 _09769_ (.A1(_03512_),
    .A2(_03514_),
    .A3(_03516_),
    .A4(_03519_),
    .ZN(_03520_));
 OAI221_X1 _09770_ (.A(_03181_),
    .B1(_03246_),
    .B2(_03510_),
    .C1(_03520_),
    .C2(_03263_),
    .ZN(_03521_));
 OAI22_X1 _09771_ (.A1(_03482_),
    .A2(_03217_),
    .B1(_03501_),
    .B2(_03521_),
    .ZN(_00368_));
 INV_X1 _09772_ (.A(net45),
    .ZN(_03522_));
 MUX2_X1 _09773_ (.A(\registers[0][17] ),
    .B(\registers[1][17] ),
    .S(_03483_),
    .Z(_03523_));
 MUX2_X1 _09774_ (.A(\registers[6][17] ),
    .B(\registers[7][17] ),
    .S(_03408_),
    .Z(_03524_));
 OAI22_X1 _09775_ (.A1(_03406_),
    .A2(_03523_),
    .B1(_03524_),
    .B2(_03410_),
    .ZN(_03525_));
 MUX2_X1 _09776_ (.A(\registers[2][17] ),
    .B(\registers[3][17] ),
    .S(_03412_),
    .Z(_03526_));
 INV_X1 _09777_ (.A(_03526_),
    .ZN(_03527_));
 AOI21_X1 _09778_ (.A(_03525_),
    .B1(_03527_),
    .B2(_03155_),
    .ZN(_03528_));
 BUF_X4 _09779_ (.A(_03139_),
    .Z(_03529_));
 MUX2_X1 _09780_ (.A(\registers[4][17] ),
    .B(\registers[5][17] ),
    .S(_03529_),
    .Z(_03530_));
 INV_X1 _09781_ (.A(_03530_),
    .ZN(_03531_));
 AOI21_X1 _09782_ (.A(_03331_),
    .B1(_03162_),
    .B2(_03531_),
    .ZN(_03532_));
 MUX2_X1 _09783_ (.A(\registers[12][17] ),
    .B(\registers[14][17] ),
    .S(_03371_),
    .Z(_03533_));
 MUX2_X1 _09784_ (.A(\registers[13][17] ),
    .B(\registers[15][17] ),
    .S(_03420_),
    .Z(_03534_));
 BUF_X4 _09785_ (.A(_03148_),
    .Z(_03535_));
 MUX2_X1 _09786_ (.A(_03533_),
    .B(_03534_),
    .S(_03535_),
    .Z(_03536_));
 MUX2_X1 _09787_ (.A(\registers[8][17] ),
    .B(\registers[10][17] ),
    .S(_03458_),
    .Z(_03537_));
 MUX2_X1 _09788_ (.A(\registers[9][17] ),
    .B(\registers[11][17] ),
    .S(_03497_),
    .Z(_03538_));
 MUX2_X1 _09789_ (.A(_03537_),
    .B(_03538_),
    .S(_03190_),
    .Z(_03539_));
 MUX2_X2 _09790_ (.A(_03536_),
    .B(_03539_),
    .S(_03462_),
    .Z(_03540_));
 AOI221_X2 _09791_ (.A(_03218_),
    .B1(_03528_),
    .B2(_03532_),
    .C1(_03540_),
    .C2(_03177_),
    .ZN(_03541_));
 BUF_X4 _09792_ (.A(_03133_),
    .Z(_03542_));
 MUX2_X1 _09793_ (.A(\registers[28][17] ),
    .B(\registers[30][17] ),
    .S(_03542_),
    .Z(_03543_));
 BUF_X4 _09794_ (.A(_03133_),
    .Z(_03544_));
 MUX2_X1 _09795_ (.A(\registers[29][17] ),
    .B(\registers[31][17] ),
    .S(_03544_),
    .Z(_03545_));
 MUX2_X1 _09796_ (.A(_03543_),
    .B(_03545_),
    .S(_03504_),
    .Z(_03546_));
 BUF_X8 _09797_ (.A(_03133_),
    .Z(_03547_));
 MUX2_X1 _09798_ (.A(\registers[24][17] ),
    .B(\registers[26][17] ),
    .S(_03547_),
    .Z(_03548_));
 BUF_X8 _09799_ (.A(_03133_),
    .Z(_03549_));
 MUX2_X1 _09800_ (.A(\registers[25][17] ),
    .B(\registers[27][17] ),
    .S(_03549_),
    .Z(_03550_));
 MUX2_X1 _09801_ (.A(_03548_),
    .B(_03550_),
    .S(_03508_),
    .Z(_03551_));
 MUX2_X1 _09802_ (.A(_03546_),
    .B(_03551_),
    .S(_03259_),
    .Z(_03552_));
 MUX2_X1 _09803_ (.A(\registers[16][17] ),
    .B(\registers[17][17] ),
    .S(_03306_),
    .Z(_03553_));
 NOR2_X1 _09804_ (.A1(_03305_),
    .A2(_03553_),
    .ZN(_03554_));
 BUF_X4 _09805_ (.A(_03219_),
    .Z(_03555_));
 MUX2_X1 _09806_ (.A(\registers[18][17] ),
    .B(\registers[19][17] ),
    .S(_03555_),
    .Z(_03556_));
 NOR3_X1 _09807_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03556_),
    .ZN(_03557_));
 MUX2_X1 _09808_ (.A(\registers[20][17] ),
    .B(\registers[21][17] ),
    .S(_03354_),
    .Z(_03558_));
 NOR3_X1 _09809_ (.A1(_03314_),
    .A2(_03315_),
    .A3(_03558_),
    .ZN(_03559_));
 MUX2_X1 _09810_ (.A(\registers[22][17] ),
    .B(\registers[23][17] ),
    .S(_03517_),
    .Z(_03560_));
 NOR2_X1 _09811_ (.A1(_03318_),
    .A2(_03560_),
    .ZN(_03561_));
 NOR4_X1 _09812_ (.A1(_03554_),
    .A2(_03557_),
    .A3(_03559_),
    .A4(_03561_),
    .ZN(_03562_));
 OAI221_X1 _09813_ (.A(_03181_),
    .B1(_03246_),
    .B2(_03552_),
    .C1(_03562_),
    .C2(_03263_),
    .ZN(_03563_));
 OAI22_X1 _09814_ (.A1(_03522_),
    .A2(_03217_),
    .B1(_03541_),
    .B2(_03563_),
    .ZN(_00369_));
 INV_X1 _09815_ (.A(net46),
    .ZN(_03564_));
 MUX2_X1 _09816_ (.A(\registers[0][18] ),
    .B(\registers[1][18] ),
    .S(_03483_),
    .Z(_03565_));
 MUX2_X1 _09817_ (.A(\registers[6][18] ),
    .B(\registers[7][18] ),
    .S(_03408_),
    .Z(_03566_));
 OAI22_X1 _09818_ (.A1(_03406_),
    .A2(_03565_),
    .B1(_03566_),
    .B2(_03410_),
    .ZN(_03567_));
 MUX2_X1 _09819_ (.A(\registers[2][18] ),
    .B(\registers[3][18] ),
    .S(_03412_),
    .Z(_03568_));
 INV_X1 _09820_ (.A(_03568_),
    .ZN(_03569_));
 AOI21_X1 _09821_ (.A(_03567_),
    .B1(_03569_),
    .B2(_03155_),
    .ZN(_03570_));
 MUX2_X1 _09822_ (.A(\registers[4][18] ),
    .B(\registers[5][18] ),
    .S(_03529_),
    .Z(_03571_));
 INV_X1 _09823_ (.A(_03571_),
    .ZN(_03572_));
 AOI21_X1 _09824_ (.A(_03331_),
    .B1(_03162_),
    .B2(_03572_),
    .ZN(_03573_));
 MUX2_X1 _09825_ (.A(\registers[12][18] ),
    .B(\registers[14][18] ),
    .S(_03371_),
    .Z(_03574_));
 MUX2_X1 _09826_ (.A(\registers[13][18] ),
    .B(\registers[15][18] ),
    .S(_03420_),
    .Z(_03575_));
 MUX2_X1 _09827_ (.A(_03574_),
    .B(_03575_),
    .S(_03535_),
    .Z(_03576_));
 MUX2_X1 _09828_ (.A(\registers[8][18] ),
    .B(\registers[10][18] ),
    .S(_03458_),
    .Z(_03577_));
 MUX2_X1 _09829_ (.A(\registers[9][18] ),
    .B(\registers[11][18] ),
    .S(_03497_),
    .Z(_03578_));
 BUF_X4 _09830_ (.A(_03169_),
    .Z(_03579_));
 MUX2_X1 _09831_ (.A(_03577_),
    .B(_03578_),
    .S(_03579_),
    .Z(_03580_));
 MUX2_X2 _09832_ (.A(_03576_),
    .B(_03580_),
    .S(_03462_),
    .Z(_03581_));
 AOI221_X2 _09833_ (.A(_03218_),
    .B1(_03570_),
    .B2(_03573_),
    .C1(_03581_),
    .C2(_03177_),
    .ZN(_03582_));
 MUX2_X1 _09834_ (.A(\registers[28][18] ),
    .B(\registers[30][18] ),
    .S(_03542_),
    .Z(_03583_));
 MUX2_X1 _09835_ (.A(\registers[29][18] ),
    .B(\registers[31][18] ),
    .S(_03544_),
    .Z(_03584_));
 MUX2_X1 _09836_ (.A(_03583_),
    .B(_03584_),
    .S(_03504_),
    .Z(_03585_));
 MUX2_X1 _09837_ (.A(\registers[24][18] ),
    .B(\registers[26][18] ),
    .S(_03547_),
    .Z(_03586_));
 MUX2_X1 _09838_ (.A(\registers[25][18] ),
    .B(\registers[27][18] ),
    .S(_03549_),
    .Z(_03587_));
 MUX2_X1 _09839_ (.A(_03586_),
    .B(_03587_),
    .S(_03508_),
    .Z(_03588_));
 MUX2_X1 _09840_ (.A(_03585_),
    .B(_03588_),
    .S(_03259_),
    .Z(_03589_));
 BUF_X4 _09841_ (.A(_03194_),
    .Z(_03590_));
 MUX2_X1 _09842_ (.A(\registers[16][18] ),
    .B(\registers[17][18] ),
    .S(_03590_),
    .Z(_03591_));
 NOR2_X1 _09843_ (.A1(_03305_),
    .A2(_03591_),
    .ZN(_03592_));
 MUX2_X1 _09844_ (.A(\registers[18][18] ),
    .B(\registers[19][18] ),
    .S(_03555_),
    .Z(_03593_));
 NOR3_X1 _09845_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03593_),
    .ZN(_03594_));
 MUX2_X1 _09846_ (.A(\registers[20][18] ),
    .B(\registers[21][18] ),
    .S(_03354_),
    .Z(_03595_));
 NOR3_X1 _09847_ (.A1(_03314_),
    .A2(_03315_),
    .A3(_03595_),
    .ZN(_03596_));
 MUX2_X1 _09848_ (.A(\registers[22][18] ),
    .B(\registers[23][18] ),
    .S(_03517_),
    .Z(_03597_));
 NOR2_X1 _09849_ (.A1(_03318_),
    .A2(_03597_),
    .ZN(_03598_));
 NOR4_X2 _09850_ (.A1(_03592_),
    .A2(_03594_),
    .A3(_03596_),
    .A4(_03598_),
    .ZN(_03599_));
 OAI221_X1 _09851_ (.A(_03181_),
    .B1(_03246_),
    .B2(_03589_),
    .C1(_03599_),
    .C2(_03263_),
    .ZN(_03600_));
 OAI22_X1 _09852_ (.A1(_03564_),
    .A2(_03217_),
    .B1(_03582_),
    .B2(_03600_),
    .ZN(_00370_));
 INV_X1 _09853_ (.A(net47),
    .ZN(_03601_));
 MUX2_X1 _09854_ (.A(\registers[0][19] ),
    .B(\registers[1][19] ),
    .S(_03483_),
    .Z(_03602_));
 MUX2_X1 _09855_ (.A(\registers[6][19] ),
    .B(\registers[7][19] ),
    .S(_03408_),
    .Z(_03603_));
 OAI22_X1 _09856_ (.A1(_03406_),
    .A2(_03602_),
    .B1(_03603_),
    .B2(_03410_),
    .ZN(_03604_));
 MUX2_X1 _09857_ (.A(\registers[2][19] ),
    .B(\registers[3][19] ),
    .S(_03412_),
    .Z(_03605_));
 INV_X1 _09858_ (.A(_03605_),
    .ZN(_03606_));
 BUF_X4 _09859_ (.A(_03154_),
    .Z(_03607_));
 AOI21_X1 _09860_ (.A(_03604_),
    .B1(_03606_),
    .B2(_03607_),
    .ZN(_03608_));
 CLKBUF_X3 _09861_ (.A(_03161_),
    .Z(_03609_));
 MUX2_X1 _09862_ (.A(\registers[4][19] ),
    .B(\registers[5][19] ),
    .S(_03529_),
    .Z(_03610_));
 INV_X1 _09863_ (.A(_03610_),
    .ZN(_03611_));
 AOI21_X1 _09864_ (.A(_03331_),
    .B1(_03609_),
    .B2(_03611_),
    .ZN(_03612_));
 MUX2_X1 _09865_ (.A(\registers[12][19] ),
    .B(\registers[14][19] ),
    .S(_03371_),
    .Z(_03613_));
 MUX2_X1 _09866_ (.A(\registers[13][19] ),
    .B(\registers[15][19] ),
    .S(_03420_),
    .Z(_03614_));
 MUX2_X1 _09867_ (.A(_03613_),
    .B(_03614_),
    .S(_03535_),
    .Z(_03615_));
 MUX2_X1 _09868_ (.A(\registers[8][19] ),
    .B(\registers[10][19] ),
    .S(_03458_),
    .Z(_03616_));
 MUX2_X1 _09869_ (.A(\registers[9][19] ),
    .B(\registers[11][19] ),
    .S(_03497_),
    .Z(_03617_));
 MUX2_X1 _09870_ (.A(_03616_),
    .B(_03617_),
    .S(_03579_),
    .Z(_03618_));
 MUX2_X2 _09871_ (.A(_03615_),
    .B(_03618_),
    .S(_03462_),
    .Z(_03619_));
 BUF_X4 _09872_ (.A(_03158_),
    .Z(_03620_));
 AOI221_X2 _09873_ (.A(_03218_),
    .B1(_03608_),
    .B2(_03612_),
    .C1(_03619_),
    .C2(_03620_),
    .ZN(_03621_));
 BUF_X4 _09874_ (.A(_03180_),
    .Z(_03622_));
 MUX2_X1 _09875_ (.A(\registers[28][19] ),
    .B(\registers[30][19] ),
    .S(_03542_),
    .Z(_03623_));
 MUX2_X1 _09876_ (.A(\registers[29][19] ),
    .B(\registers[31][19] ),
    .S(_03544_),
    .Z(_03624_));
 MUX2_X1 _09877_ (.A(_03623_),
    .B(_03624_),
    .S(_03504_),
    .Z(_03625_));
 MUX2_X1 _09878_ (.A(\registers[24][19] ),
    .B(\registers[26][19] ),
    .S(_03547_),
    .Z(_03626_));
 MUX2_X1 _09879_ (.A(\registers[25][19] ),
    .B(\registers[27][19] ),
    .S(_03549_),
    .Z(_03627_));
 MUX2_X1 _09880_ (.A(_03626_),
    .B(_03627_),
    .S(_03508_),
    .Z(_03628_));
 BUF_X4 _09881_ (.A(_03258_),
    .Z(_03629_));
 MUX2_X1 _09882_ (.A(_03625_),
    .B(_03628_),
    .S(_03629_),
    .Z(_03630_));
 MUX2_X1 _09883_ (.A(\registers[16][19] ),
    .B(\registers[17][19] ),
    .S(_03590_),
    .Z(_03631_));
 NOR2_X1 _09884_ (.A1(_03305_),
    .A2(_03631_),
    .ZN(_03632_));
 MUX2_X1 _09885_ (.A(\registers[18][19] ),
    .B(\registers[19][19] ),
    .S(_03555_),
    .Z(_03633_));
 NOR3_X1 _09886_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03633_),
    .ZN(_03634_));
 MUX2_X1 _09887_ (.A(\registers[20][19] ),
    .B(\registers[21][19] ),
    .S(_03354_),
    .Z(_03635_));
 NOR3_X1 _09888_ (.A1(_03314_),
    .A2(_03315_),
    .A3(_03635_),
    .ZN(_03636_));
 MUX2_X1 _09889_ (.A(\registers[22][19] ),
    .B(\registers[23][19] ),
    .S(_03517_),
    .Z(_03637_));
 NOR2_X1 _09890_ (.A1(_03318_),
    .A2(_03637_),
    .ZN(_03638_));
 NOR4_X2 _09891_ (.A1(_03632_),
    .A2(_03634_),
    .A3(_03636_),
    .A4(_03638_),
    .ZN(_03639_));
 OAI221_X1 _09892_ (.A(_03622_),
    .B1(_03246_),
    .B2(_03630_),
    .C1(_03639_),
    .C2(_03263_),
    .ZN(_03640_));
 OAI22_X1 _09893_ (.A1(_03601_),
    .A2(_03217_),
    .B1(_03621_),
    .B2(_03640_),
    .ZN(_00371_));
 INV_X1 _09894_ (.A(net48),
    .ZN(_03641_));
 CLKBUF_X3 _09895_ (.A(_03214_),
    .Z(_03642_));
 MUX2_X1 _09896_ (.A(\registers[16][1] ),
    .B(\registers[17][1] ),
    .S(_03483_),
    .Z(_03643_));
 MUX2_X1 _09897_ (.A(\registers[22][1] ),
    .B(\registers[23][1] ),
    .S(_03408_),
    .Z(_03644_));
 OAI22_X1 _09898_ (.A1(_03406_),
    .A2(_03643_),
    .B1(_03644_),
    .B2(_03410_),
    .ZN(_03645_));
 MUX2_X1 _09899_ (.A(\registers[18][1] ),
    .B(\registers[19][1] ),
    .S(_03412_),
    .Z(_03646_));
 INV_X1 _09900_ (.A(_03646_),
    .ZN(_03647_));
 AOI21_X1 _09901_ (.A(_03645_),
    .B1(_03647_),
    .B2(_03607_),
    .ZN(_03648_));
 MUX2_X1 _09902_ (.A(\registers[20][1] ),
    .B(\registers[21][1] ),
    .S(_03529_),
    .Z(_03649_));
 INV_X1 _09903_ (.A(_03649_),
    .ZN(_03650_));
 AOI21_X1 _09904_ (.A(_03331_),
    .B1(_03609_),
    .B2(_03650_),
    .ZN(_03651_));
 MUX2_X1 _09905_ (.A(\registers[28][1] ),
    .B(\registers[30][1] ),
    .S(_03371_),
    .Z(_03652_));
 MUX2_X1 _09906_ (.A(\registers[29][1] ),
    .B(\registers[31][1] ),
    .S(_03420_),
    .Z(_03653_));
 MUX2_X1 _09907_ (.A(_03652_),
    .B(_03653_),
    .S(_03535_),
    .Z(_03654_));
 MUX2_X1 _09908_ (.A(\registers[24][1] ),
    .B(\registers[26][1] ),
    .S(_03458_),
    .Z(_03655_));
 MUX2_X1 _09909_ (.A(\registers[25][1] ),
    .B(\registers[27][1] ),
    .S(_03497_),
    .Z(_03656_));
 MUX2_X1 _09910_ (.A(_03655_),
    .B(_03656_),
    .S(_03579_),
    .Z(_03657_));
 MUX2_X1 _09911_ (.A(_03654_),
    .B(_03657_),
    .S(_03462_),
    .Z(_03658_));
 AOI221_X1 _09912_ (.A(_03131_),
    .B1(_03648_),
    .B2(_03651_),
    .C1(_03658_),
    .C2(_03620_),
    .ZN(_03659_));
 MUX2_X1 _09913_ (.A(\registers[0][1] ),
    .B(\registers[1][1] ),
    .S(_03380_),
    .Z(_03660_));
 NOR2_X1 _09914_ (.A1(_03184_),
    .A2(_03660_),
    .ZN(_03661_));
 MUX2_X1 _09915_ (.A(\registers[2][1] ),
    .B(\registers[3][1] ),
    .S(_03163_),
    .Z(_03662_));
 NOR3_X1 _09916_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_03662_),
    .ZN(_03663_));
 MUX2_X1 _09917_ (.A(\registers[4][1] ),
    .B(\registers[5][1] ),
    .S(_03386_),
    .Z(_03664_));
 NOR3_X1 _09918_ (.A1(_03193_),
    .A2(_03385_),
    .A3(_03664_),
    .ZN(_03665_));
 MUX2_X1 _09919_ (.A(\registers[6][1] ),
    .B(\registers[7][1] ),
    .S(_03272_),
    .Z(_03666_));
 NOR2_X1 _09920_ (.A1(_03197_),
    .A2(_03666_),
    .ZN(_03667_));
 NOR4_X2 _09921_ (.A1(_03661_),
    .A2(_03663_),
    .A3(_03665_),
    .A4(_03667_),
    .ZN(_03668_));
 MUX2_X1 _09922_ (.A(\registers[12][1] ),
    .B(\registers[14][1] ),
    .S(_03392_),
    .Z(_03669_));
 MUX2_X1 _09923_ (.A(\registers[13][1] ),
    .B(\registers[15][1] ),
    .S(_03394_),
    .Z(_03670_));
 MUX2_X1 _09924_ (.A(_03669_),
    .B(_03670_),
    .S(_03396_),
    .Z(_03671_));
 MUX2_X1 _09925_ (.A(\registers[8][1] ),
    .B(\registers[10][1] ),
    .S(_03398_),
    .Z(_03672_));
 MUX2_X1 _09926_ (.A(\registers[9][1] ),
    .B(\registers[11][1] ),
    .S(_03400_),
    .Z(_03673_));
 MUX2_X1 _09927_ (.A(_03672_),
    .B(_03673_),
    .S(_03203_),
    .Z(_03674_));
 MUX2_X2 _09928_ (.A(_03671_),
    .B(_03674_),
    .S(_03208_),
    .Z(_03675_));
 OAI221_X2 _09929_ (.A(_03622_),
    .B1(_03183_),
    .B2(_03668_),
    .C1(_03675_),
    .C2(_03211_),
    .ZN(_03676_));
 OAI22_X1 _09930_ (.A1(_03641_),
    .A2(_03642_),
    .B1(_03659_),
    .B2(_03676_),
    .ZN(_00372_));
 INV_X1 _09931_ (.A(net49),
    .ZN(_03677_));
 MUX2_X1 _09932_ (.A(\registers[0][20] ),
    .B(\registers[1][20] ),
    .S(_03483_),
    .Z(_03678_));
 MUX2_X1 _09933_ (.A(\registers[6][20] ),
    .B(\registers[7][20] ),
    .S(_03408_),
    .Z(_03679_));
 OAI22_X1 _09934_ (.A1(_03406_),
    .A2(_03678_),
    .B1(_03679_),
    .B2(_03410_),
    .ZN(_03680_));
 MUX2_X1 _09935_ (.A(\registers[2][20] ),
    .B(\registers[3][20] ),
    .S(_03412_),
    .Z(_03681_));
 INV_X1 _09936_ (.A(_03681_),
    .ZN(_03682_));
 AOI21_X1 _09937_ (.A(_03680_),
    .B1(_03682_),
    .B2(_03607_),
    .ZN(_03683_));
 MUX2_X1 _09938_ (.A(\registers[4][20] ),
    .B(\registers[5][20] ),
    .S(_03529_),
    .Z(_03684_));
 INV_X1 _09939_ (.A(_03684_),
    .ZN(_03685_));
 AOI21_X1 _09940_ (.A(_03331_),
    .B1(_03609_),
    .B2(_03685_),
    .ZN(_03686_));
 MUX2_X1 _09941_ (.A(\registers[12][20] ),
    .B(\registers[14][20] ),
    .S(_03371_),
    .Z(_03687_));
 MUX2_X1 _09942_ (.A(\registers[13][20] ),
    .B(\registers[15][20] ),
    .S(_03420_),
    .Z(_03688_));
 MUX2_X1 _09943_ (.A(_03687_),
    .B(_03688_),
    .S(_03535_),
    .Z(_03689_));
 MUX2_X1 _09944_ (.A(\registers[8][20] ),
    .B(\registers[10][20] ),
    .S(_03458_),
    .Z(_03690_));
 MUX2_X1 _09945_ (.A(\registers[9][20] ),
    .B(\registers[11][20] ),
    .S(_03497_),
    .Z(_03691_));
 MUX2_X1 _09946_ (.A(_03690_),
    .B(_03691_),
    .S(_03579_),
    .Z(_03692_));
 MUX2_X2 _09947_ (.A(_03689_),
    .B(_03692_),
    .S(_03462_),
    .Z(_03693_));
 AOI221_X2 _09948_ (.A(_03218_),
    .B1(_03683_),
    .B2(_03686_),
    .C1(_03693_),
    .C2(_03620_),
    .ZN(_03694_));
 MUX2_X1 _09949_ (.A(\registers[28][20] ),
    .B(\registers[30][20] ),
    .S(_03542_),
    .Z(_03695_));
 MUX2_X1 _09950_ (.A(\registers[29][20] ),
    .B(\registers[31][20] ),
    .S(_03544_),
    .Z(_03696_));
 MUX2_X1 _09951_ (.A(_03695_),
    .B(_03696_),
    .S(_03504_),
    .Z(_03697_));
 MUX2_X1 _09952_ (.A(\registers[24][20] ),
    .B(\registers[26][20] ),
    .S(_03547_),
    .Z(_03698_));
 MUX2_X1 _09953_ (.A(\registers[25][20] ),
    .B(\registers[27][20] ),
    .S(_03549_),
    .Z(_03699_));
 MUX2_X1 _09954_ (.A(_03698_),
    .B(_03699_),
    .S(_03508_),
    .Z(_03700_));
 MUX2_X1 _09955_ (.A(_03697_),
    .B(_03700_),
    .S(_03629_),
    .Z(_03701_));
 MUX2_X1 _09956_ (.A(\registers[16][20] ),
    .B(\registers[17][20] ),
    .S(_03590_),
    .Z(_03702_));
 NOR2_X1 _09957_ (.A1(_03305_),
    .A2(_03702_),
    .ZN(_03703_));
 MUX2_X1 _09958_ (.A(\registers[18][20] ),
    .B(\registers[19][20] ),
    .S(_03555_),
    .Z(_03704_));
 NOR3_X1 _09959_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03704_),
    .ZN(_03705_));
 BUF_X4 _09960_ (.A(_03258_),
    .Z(_03706_));
 MUX2_X1 _09961_ (.A(\registers[20][20] ),
    .B(\registers[21][20] ),
    .S(_03354_),
    .Z(_03707_));
 NOR3_X1 _09962_ (.A1(_03314_),
    .A2(_03706_),
    .A3(_03707_),
    .ZN(_03708_));
 MUX2_X1 _09963_ (.A(\registers[22][20] ),
    .B(\registers[23][20] ),
    .S(_03517_),
    .Z(_03709_));
 NOR2_X1 _09964_ (.A1(_03318_),
    .A2(_03709_),
    .ZN(_03710_));
 NOR4_X2 _09965_ (.A1(_03703_),
    .A2(_03705_),
    .A3(_03708_),
    .A4(_03710_),
    .ZN(_03711_));
 OAI221_X1 _09966_ (.A(_03622_),
    .B1(_03246_),
    .B2(_03701_),
    .C1(_03711_),
    .C2(_03263_),
    .ZN(_03712_));
 OAI22_X1 _09967_ (.A1(_03677_),
    .A2(_03642_),
    .B1(_03694_),
    .B2(_03712_),
    .ZN(_00373_));
 INV_X1 _09968_ (.A(net50),
    .ZN(_03713_));
 BUF_X4 _09969_ (.A(_03129_),
    .Z(_03714_));
 MUX2_X1 _09970_ (.A(\registers[0][21] ),
    .B(\registers[1][21] ),
    .S(_03483_),
    .Z(_03715_));
 MUX2_X1 _09971_ (.A(\registers[6][21] ),
    .B(\registers[7][21] ),
    .S(_03408_),
    .Z(_03716_));
 OAI22_X1 _09972_ (.A1(_03406_),
    .A2(_03715_),
    .B1(_03716_),
    .B2(_03410_),
    .ZN(_03717_));
 MUX2_X1 _09973_ (.A(\registers[2][21] ),
    .B(\registers[3][21] ),
    .S(_03412_),
    .Z(_03718_));
 INV_X1 _09974_ (.A(_03718_),
    .ZN(_03719_));
 AOI21_X1 _09975_ (.A(_03717_),
    .B1(_03719_),
    .B2(_03607_),
    .ZN(_03720_));
 CLKBUF_X3 _09976_ (.A(_03157_),
    .Z(_03721_));
 MUX2_X1 _09977_ (.A(\registers[4][21] ),
    .B(\registers[5][21] ),
    .S(_03529_),
    .Z(_03722_));
 INV_X1 _09978_ (.A(_03722_),
    .ZN(_03723_));
 AOI21_X1 _09979_ (.A(_03721_),
    .B1(_03609_),
    .B2(_03723_),
    .ZN(_03724_));
 MUX2_X1 _09980_ (.A(\registers[12][21] ),
    .B(\registers[14][21] ),
    .S(_03371_),
    .Z(_03725_));
 MUX2_X1 _09981_ (.A(\registers[13][21] ),
    .B(\registers[15][21] ),
    .S(_03420_),
    .Z(_03726_));
 MUX2_X1 _09982_ (.A(_03725_),
    .B(_03726_),
    .S(_03535_),
    .Z(_03727_));
 MUX2_X1 _09983_ (.A(\registers[8][21] ),
    .B(\registers[10][21] ),
    .S(_03458_),
    .Z(_03728_));
 MUX2_X1 _09984_ (.A(\registers[9][21] ),
    .B(\registers[11][21] ),
    .S(_03497_),
    .Z(_03729_));
 MUX2_X1 _09985_ (.A(_03728_),
    .B(_03729_),
    .S(_03579_),
    .Z(_03730_));
 MUX2_X2 _09986_ (.A(_03727_),
    .B(_03730_),
    .S(_03462_),
    .Z(_03731_));
 AOI221_X2 _09987_ (.A(_03714_),
    .B1(_03720_),
    .B2(_03724_),
    .C1(_03731_),
    .C2(_03620_),
    .ZN(_03732_));
 CLKBUF_X3 _09988_ (.A(_03245_),
    .Z(_03733_));
 MUX2_X1 _09989_ (.A(\registers[28][21] ),
    .B(\registers[30][21] ),
    .S(_03542_),
    .Z(_03734_));
 MUX2_X1 _09990_ (.A(\registers[29][21] ),
    .B(\registers[31][21] ),
    .S(_03544_),
    .Z(_03735_));
 MUX2_X1 _09991_ (.A(_03734_),
    .B(_03735_),
    .S(_03504_),
    .Z(_03736_));
 MUX2_X1 _09992_ (.A(\registers[24][21] ),
    .B(\registers[26][21] ),
    .S(_03547_),
    .Z(_03737_));
 MUX2_X1 _09993_ (.A(\registers[25][21] ),
    .B(\registers[27][21] ),
    .S(_03549_),
    .Z(_03738_));
 MUX2_X1 _09994_ (.A(_03737_),
    .B(_03738_),
    .S(_03508_),
    .Z(_03739_));
 MUX2_X1 _09995_ (.A(_03736_),
    .B(_03739_),
    .S(_03629_),
    .Z(_03740_));
 MUX2_X1 _09996_ (.A(\registers[16][21] ),
    .B(\registers[17][21] ),
    .S(_03590_),
    .Z(_03741_));
 NOR2_X1 _09997_ (.A1(_03305_),
    .A2(_03741_),
    .ZN(_03742_));
 MUX2_X1 _09998_ (.A(\registers[18][21] ),
    .B(\registers[19][21] ),
    .S(_03555_),
    .Z(_03743_));
 NOR3_X1 _09999_ (.A1(_03309_),
    .A2(_03310_),
    .A3(_03743_),
    .ZN(_03744_));
 MUX2_X1 _10000_ (.A(\registers[20][21] ),
    .B(\registers[21][21] ),
    .S(_03354_),
    .Z(_03745_));
 NOR3_X1 _10001_ (.A1(_03314_),
    .A2(_03706_),
    .A3(_03745_),
    .ZN(_03746_));
 MUX2_X1 _10002_ (.A(\registers[22][21] ),
    .B(\registers[23][21] ),
    .S(_03517_),
    .Z(_03747_));
 NOR2_X1 _10003_ (.A1(_03318_),
    .A2(_03747_),
    .ZN(_03748_));
 NOR4_X1 _10004_ (.A1(_03742_),
    .A2(_03744_),
    .A3(_03746_),
    .A4(_03748_),
    .ZN(_03749_));
 CLKBUF_X3 _10005_ (.A(_03262_),
    .Z(_03750_));
 OAI221_X1 _10006_ (.A(_03622_),
    .B1(_03733_),
    .B2(_03740_),
    .C1(_03749_),
    .C2(_03750_),
    .ZN(_03751_));
 OAI22_X1 _10007_ (.A1(_03713_),
    .A2(_03642_),
    .B1(_03732_),
    .B2(_03751_),
    .ZN(_00374_));
 INV_X1 _10008_ (.A(net51),
    .ZN(_03752_));
 MUX2_X1 _10009_ (.A(\registers[16][22] ),
    .B(\registers[17][22] ),
    .S(_03483_),
    .Z(_03753_));
 MUX2_X1 _10010_ (.A(\registers[22][22] ),
    .B(\registers[23][22] ),
    .S(_03408_),
    .Z(_03754_));
 OAI22_X1 _10011_ (.A1(_03406_),
    .A2(_03753_),
    .B1(_03754_),
    .B2(_03410_),
    .ZN(_03755_));
 MUX2_X1 _10012_ (.A(\registers[18][22] ),
    .B(\registers[19][22] ),
    .S(_03412_),
    .Z(_03756_));
 INV_X1 _10013_ (.A(_03756_),
    .ZN(_03757_));
 AOI21_X1 _10014_ (.A(_03755_),
    .B1(_03757_),
    .B2(_03607_),
    .ZN(_03758_));
 MUX2_X1 _10015_ (.A(\registers[20][22] ),
    .B(\registers[21][22] ),
    .S(_03529_),
    .Z(_03759_));
 INV_X1 _10016_ (.A(_03759_),
    .ZN(_03760_));
 AOI21_X1 _10017_ (.A(_03721_),
    .B1(_03609_),
    .B2(_03760_),
    .ZN(_03761_));
 BUF_X4 _10018_ (.A(_03231_),
    .Z(_03762_));
 MUX2_X1 _10019_ (.A(\registers[28][22] ),
    .B(\registers[30][22] ),
    .S(_03762_),
    .Z(_03763_));
 MUX2_X1 _10020_ (.A(\registers[29][22] ),
    .B(\registers[31][22] ),
    .S(_03420_),
    .Z(_03764_));
 MUX2_X1 _10021_ (.A(_03763_),
    .B(_03764_),
    .S(_03535_),
    .Z(_03765_));
 MUX2_X1 _10022_ (.A(\registers[24][22] ),
    .B(\registers[26][22] ),
    .S(_03458_),
    .Z(_03766_));
 MUX2_X1 _10023_ (.A(\registers[25][22] ),
    .B(\registers[27][22] ),
    .S(_03497_),
    .Z(_03767_));
 MUX2_X1 _10024_ (.A(_03766_),
    .B(_03767_),
    .S(_03579_),
    .Z(_03768_));
 MUX2_X1 _10025_ (.A(_03765_),
    .B(_03768_),
    .S(_03462_),
    .Z(_03769_));
 AOI221_X1 _10026_ (.A(_03131_),
    .B1(_03758_),
    .B2(_03761_),
    .C1(_03769_),
    .C2(_03620_),
    .ZN(_03770_));
 MUX2_X1 _10027_ (.A(\registers[0][22] ),
    .B(\registers[1][22] ),
    .S(_03380_),
    .Z(_03771_));
 NOR2_X1 _10028_ (.A1(_03184_),
    .A2(_03771_),
    .ZN(_03772_));
 MUX2_X1 _10029_ (.A(\registers[2][22] ),
    .B(\registers[3][22] ),
    .S(_03163_),
    .Z(_03773_));
 NOR3_X1 _10030_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_03773_),
    .ZN(_03774_));
 MUX2_X1 _10031_ (.A(\registers[4][22] ),
    .B(\registers[5][22] ),
    .S(_03386_),
    .Z(_03775_));
 NOR3_X1 _10032_ (.A1(_03193_),
    .A2(_03385_),
    .A3(_03775_),
    .ZN(_03776_));
 MUX2_X1 _10033_ (.A(\registers[6][22] ),
    .B(\registers[7][22] ),
    .S(_03272_),
    .Z(_03777_));
 NOR2_X1 _10034_ (.A1(_03197_),
    .A2(_03777_),
    .ZN(_03778_));
 NOR4_X2 _10035_ (.A1(_03772_),
    .A2(_03774_),
    .A3(_03776_),
    .A4(_03778_),
    .ZN(_03779_));
 MUX2_X1 _10036_ (.A(\registers[12][22] ),
    .B(\registers[14][22] ),
    .S(_03392_),
    .Z(_03780_));
 MUX2_X1 _10037_ (.A(\registers[13][22] ),
    .B(\registers[15][22] ),
    .S(_03394_),
    .Z(_03781_));
 MUX2_X1 _10038_ (.A(_03780_),
    .B(_03781_),
    .S(_03396_),
    .Z(_03782_));
 MUX2_X1 _10039_ (.A(\registers[8][22] ),
    .B(\registers[10][22] ),
    .S(_03398_),
    .Z(_03783_));
 MUX2_X1 _10040_ (.A(\registers[9][22] ),
    .B(\registers[11][22] ),
    .S(_03400_),
    .Z(_03784_));
 MUX2_X1 _10041_ (.A(_03783_),
    .B(_03784_),
    .S(_03203_),
    .Z(_03785_));
 MUX2_X2 _10042_ (.A(_03782_),
    .B(_03785_),
    .S(_03208_),
    .Z(_03786_));
 OAI221_X2 _10043_ (.A(_03622_),
    .B1(_03183_),
    .B2(_03779_),
    .C1(_03786_),
    .C2(_03211_),
    .ZN(_03787_));
 OAI22_X1 _10044_ (.A1(_03752_),
    .A2(_03642_),
    .B1(_03770_),
    .B2(_03787_),
    .ZN(_00375_));
 INV_X1 _10045_ (.A(net52),
    .ZN(_03788_));
 BUF_X4 _10046_ (.A(_03136_),
    .Z(_03789_));
 MUX2_X1 _10047_ (.A(\registers[16][23] ),
    .B(\registers[17][23] ),
    .S(_03483_),
    .Z(_03790_));
 BUF_X4 _10048_ (.A(_03138_),
    .Z(_03791_));
 MUX2_X1 _10049_ (.A(\registers[22][23] ),
    .B(\registers[23][23] ),
    .S(_03791_),
    .Z(_03792_));
 BUF_X4 _10050_ (.A(_03143_),
    .Z(_03793_));
 OAI22_X1 _10051_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03792_),
    .B2(_03793_),
    .ZN(_03794_));
 BUF_X4 _10052_ (.A(_03148_),
    .Z(_03795_));
 MUX2_X1 _10053_ (.A(\registers[18][23] ),
    .B(\registers[19][23] ),
    .S(_03795_),
    .Z(_03796_));
 INV_X1 _10054_ (.A(_03796_),
    .ZN(_03797_));
 AOI21_X1 _10055_ (.A(_03794_),
    .B1(_03797_),
    .B2(_03607_),
    .ZN(_03798_));
 MUX2_X1 _10056_ (.A(\registers[20][23] ),
    .B(\registers[21][23] ),
    .S(_03529_),
    .Z(_03799_));
 INV_X1 _10057_ (.A(_03799_),
    .ZN(_03800_));
 AOI21_X1 _10058_ (.A(_03721_),
    .B1(_03609_),
    .B2(_03800_),
    .ZN(_03801_));
 MUX2_X1 _10059_ (.A(\registers[28][23] ),
    .B(\registers[30][23] ),
    .S(_03762_),
    .Z(_03802_));
 BUF_X4 _10060_ (.A(_03231_),
    .Z(_03803_));
 MUX2_X1 _10061_ (.A(\registers[29][23] ),
    .B(\registers[31][23] ),
    .S(_03803_),
    .Z(_03804_));
 MUX2_X1 _10062_ (.A(_03802_),
    .B(_03804_),
    .S(_03535_),
    .Z(_03805_));
 MUX2_X1 _10063_ (.A(\registers[24][23] ),
    .B(\registers[26][23] ),
    .S(_03458_),
    .Z(_03806_));
 MUX2_X1 _10064_ (.A(\registers[25][23] ),
    .B(\registers[27][23] ),
    .S(_03497_),
    .Z(_03807_));
 MUX2_X1 _10065_ (.A(_03806_),
    .B(_03807_),
    .S(_03579_),
    .Z(_03808_));
 MUX2_X1 _10066_ (.A(_03805_),
    .B(_03808_),
    .S(_03462_),
    .Z(_03809_));
 AOI221_X1 _10067_ (.A(_03131_),
    .B1(_03798_),
    .B2(_03801_),
    .C1(_03809_),
    .C2(_03620_),
    .ZN(_03810_));
 MUX2_X1 _10068_ (.A(\registers[0][23] ),
    .B(\registers[1][23] ),
    .S(_03380_),
    .Z(_03811_));
 NOR2_X1 _10069_ (.A1(_03184_),
    .A2(_03811_),
    .ZN(_03812_));
 MUX2_X1 _10070_ (.A(\registers[2][23] ),
    .B(\registers[3][23] ),
    .S(_03163_),
    .Z(_03813_));
 NOR3_X1 _10071_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_03813_),
    .ZN(_03814_));
 MUX2_X1 _10072_ (.A(\registers[4][23] ),
    .B(\registers[5][23] ),
    .S(_03386_),
    .Z(_03815_));
 NOR3_X1 _10073_ (.A1(_03193_),
    .A2(_03385_),
    .A3(_03815_),
    .ZN(_03816_));
 MUX2_X1 _10074_ (.A(\registers[6][23] ),
    .B(\registers[7][23] ),
    .S(_03272_),
    .Z(_03817_));
 NOR2_X1 _10075_ (.A1(_03197_),
    .A2(_03817_),
    .ZN(_03818_));
 NOR4_X2 _10076_ (.A1(_03812_),
    .A2(_03814_),
    .A3(_03816_),
    .A4(_03818_),
    .ZN(_03819_));
 MUX2_X1 _10077_ (.A(\registers[12][23] ),
    .B(\registers[14][23] ),
    .S(_03392_),
    .Z(_03820_));
 MUX2_X1 _10078_ (.A(\registers[13][23] ),
    .B(\registers[15][23] ),
    .S(_03394_),
    .Z(_03821_));
 MUX2_X1 _10079_ (.A(_03820_),
    .B(_03821_),
    .S(_03396_),
    .Z(_03822_));
 MUX2_X1 _10080_ (.A(\registers[8][23] ),
    .B(\registers[10][23] ),
    .S(_03398_),
    .Z(_03823_));
 MUX2_X1 _10081_ (.A(\registers[9][23] ),
    .B(\registers[11][23] ),
    .S(_03400_),
    .Z(_03824_));
 MUX2_X1 _10082_ (.A(_03823_),
    .B(_03824_),
    .S(_03203_),
    .Z(_03825_));
 MUX2_X2 _10083_ (.A(_03822_),
    .B(_03825_),
    .S(_03208_),
    .Z(_03826_));
 OAI221_X2 _10084_ (.A(_03622_),
    .B1(_03183_),
    .B2(_03819_),
    .C1(_03826_),
    .C2(_03211_),
    .ZN(_03827_));
 OAI22_X1 _10085_ (.A1(_03788_),
    .A2(_03642_),
    .B1(_03810_),
    .B2(_03827_),
    .ZN(_00376_));
 INV_X1 _10086_ (.A(net53),
    .ZN(_03828_));
 MUX2_X1 _10087_ (.A(\registers[16][24] ),
    .B(\registers[17][24] ),
    .S(_03483_),
    .Z(_03829_));
 MUX2_X1 _10088_ (.A(\registers[22][24] ),
    .B(\registers[23][24] ),
    .S(_03791_),
    .Z(_03830_));
 OAI22_X1 _10089_ (.A1(_03789_),
    .A2(_03829_),
    .B1(_03830_),
    .B2(_03793_),
    .ZN(_03831_));
 MUX2_X1 _10090_ (.A(\registers[18][24] ),
    .B(\registers[19][24] ),
    .S(_03795_),
    .Z(_03832_));
 INV_X1 _10091_ (.A(_03832_),
    .ZN(_03833_));
 AOI21_X1 _10092_ (.A(_03831_),
    .B1(_03833_),
    .B2(_03607_),
    .ZN(_03834_));
 MUX2_X1 _10093_ (.A(\registers[20][24] ),
    .B(\registers[21][24] ),
    .S(_03529_),
    .Z(_03835_));
 INV_X1 _10094_ (.A(_03835_),
    .ZN(_03836_));
 AOI21_X1 _10095_ (.A(_03721_),
    .B1(_03609_),
    .B2(_03836_),
    .ZN(_03837_));
 MUX2_X1 _10096_ (.A(\registers[28][24] ),
    .B(\registers[30][24] ),
    .S(_03762_),
    .Z(_03838_));
 MUX2_X1 _10097_ (.A(\registers[29][24] ),
    .B(\registers[31][24] ),
    .S(_03803_),
    .Z(_03839_));
 MUX2_X1 _10098_ (.A(_03838_),
    .B(_03839_),
    .S(_03535_),
    .Z(_03840_));
 BUF_X4 _10099_ (.A(_03231_),
    .Z(_03841_));
 MUX2_X1 _10100_ (.A(\registers[24][24] ),
    .B(\registers[26][24] ),
    .S(_03841_),
    .Z(_03842_));
 MUX2_X1 _10101_ (.A(\registers[25][24] ),
    .B(\registers[27][24] ),
    .S(_03497_),
    .Z(_03843_));
 MUX2_X1 _10102_ (.A(_03842_),
    .B(_03843_),
    .S(_03579_),
    .Z(_03844_));
 BUF_X4 _10103_ (.A(_03160_),
    .Z(_03845_));
 MUX2_X1 _10104_ (.A(_03840_),
    .B(_03844_),
    .S(_03845_),
    .Z(_03846_));
 AOI221_X1 _10105_ (.A(_03131_),
    .B1(_03834_),
    .B2(_03837_),
    .C1(_03846_),
    .C2(_03620_),
    .ZN(_03847_));
 MUX2_X1 _10106_ (.A(\registers[0][24] ),
    .B(\registers[1][24] ),
    .S(_03380_),
    .Z(_03848_));
 NOR2_X1 _10107_ (.A1(_03184_),
    .A2(_03848_),
    .ZN(_03849_));
 MUX2_X1 _10108_ (.A(\registers[2][24] ),
    .B(\registers[3][24] ),
    .S(_03163_),
    .Z(_03850_));
 NOR3_X1 _10109_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_03850_),
    .ZN(_03851_));
 MUX2_X1 _10110_ (.A(\registers[4][24] ),
    .B(\registers[5][24] ),
    .S(_03386_),
    .Z(_03852_));
 NOR3_X1 _10111_ (.A1(_03193_),
    .A2(_03258_),
    .A3(_03852_),
    .ZN(_03853_));
 MUX2_X1 _10112_ (.A(\registers[6][24] ),
    .B(\registers[7][24] ),
    .S(_03272_),
    .Z(_03854_));
 NOR2_X1 _10113_ (.A1(_03197_),
    .A2(_03854_),
    .ZN(_03855_));
 NOR4_X2 _10114_ (.A1(_03849_),
    .A2(_03851_),
    .A3(_03853_),
    .A4(_03855_),
    .ZN(_03856_));
 MUX2_X1 _10115_ (.A(\registers[12][24] ),
    .B(\registers[14][24] ),
    .S(_03392_),
    .Z(_03857_));
 MUX2_X1 _10116_ (.A(\registers[13][24] ),
    .B(\registers[15][24] ),
    .S(_03394_),
    .Z(_03858_));
 MUX2_X1 _10117_ (.A(_03857_),
    .B(_03858_),
    .S(_03396_),
    .Z(_03859_));
 MUX2_X1 _10118_ (.A(\registers[8][24] ),
    .B(\registers[10][24] ),
    .S(_03398_),
    .Z(_03860_));
 MUX2_X1 _10119_ (.A(\registers[9][24] ),
    .B(\registers[11][24] ),
    .S(_03400_),
    .Z(_03861_));
 MUX2_X1 _10120_ (.A(_03860_),
    .B(_03861_),
    .S(_03203_),
    .Z(_03862_));
 MUX2_X2 _10121_ (.A(_03859_),
    .B(_03862_),
    .S(_03208_),
    .Z(_03863_));
 OAI221_X2 _10122_ (.A(_03622_),
    .B1(_03183_),
    .B2(_03856_),
    .C1(_03863_),
    .C2(_03211_),
    .ZN(_03864_));
 OAI22_X1 _10123_ (.A1(_03828_),
    .A2(_03642_),
    .B1(_03847_),
    .B2(_03864_),
    .ZN(_00377_));
 INV_X1 _10124_ (.A(net54),
    .ZN(_03865_));
 BUF_X4 _10125_ (.A(_03139_),
    .Z(_03866_));
 MUX2_X1 _10126_ (.A(\registers[0][25] ),
    .B(\registers[1][25] ),
    .S(_03866_),
    .Z(_03867_));
 MUX2_X1 _10127_ (.A(\registers[6][25] ),
    .B(\registers[7][25] ),
    .S(_03791_),
    .Z(_03868_));
 OAI22_X1 _10128_ (.A1(_03789_),
    .A2(_03867_),
    .B1(_03868_),
    .B2(_03793_),
    .ZN(_03869_));
 MUX2_X1 _10129_ (.A(\registers[2][25] ),
    .B(\registers[3][25] ),
    .S(_03795_),
    .Z(_03870_));
 INV_X1 _10130_ (.A(_03870_),
    .ZN(_03871_));
 AOI21_X1 _10131_ (.A(_03869_),
    .B1(_03871_),
    .B2(_03607_),
    .ZN(_03872_));
 MUX2_X1 _10132_ (.A(\registers[4][25] ),
    .B(\registers[5][25] ),
    .S(_03529_),
    .Z(_03873_));
 INV_X1 _10133_ (.A(_03873_),
    .ZN(_03874_));
 AOI21_X1 _10134_ (.A(_03721_),
    .B1(_03609_),
    .B2(_03874_),
    .ZN(_03875_));
 MUX2_X1 _10135_ (.A(\registers[12][25] ),
    .B(\registers[14][25] ),
    .S(_03762_),
    .Z(_03876_));
 MUX2_X1 _10136_ (.A(\registers[13][25] ),
    .B(\registers[15][25] ),
    .S(_03803_),
    .Z(_03877_));
 MUX2_X1 _10137_ (.A(_03876_),
    .B(_03877_),
    .S(_03535_),
    .Z(_03878_));
 MUX2_X1 _10138_ (.A(\registers[8][25] ),
    .B(\registers[10][25] ),
    .S(_03841_),
    .Z(_03879_));
 BUF_X4 _10139_ (.A(_03231_),
    .Z(_03880_));
 MUX2_X1 _10140_ (.A(\registers[9][25] ),
    .B(\registers[11][25] ),
    .S(_03880_),
    .Z(_03881_));
 MUX2_X1 _10141_ (.A(_03879_),
    .B(_03881_),
    .S(_03579_),
    .Z(_03882_));
 MUX2_X2 _10142_ (.A(_03878_),
    .B(_03882_),
    .S(_03845_),
    .Z(_03883_));
 AOI221_X2 _10143_ (.A(_03714_),
    .B1(_03872_),
    .B2(_03875_),
    .C1(_03883_),
    .C2(_03620_),
    .ZN(_03884_));
 MUX2_X1 _10144_ (.A(\registers[28][25] ),
    .B(\registers[30][25] ),
    .S(_03542_),
    .Z(_03885_));
 MUX2_X1 _10145_ (.A(\registers[29][25] ),
    .B(\registers[31][25] ),
    .S(_03544_),
    .Z(_03886_));
 MUX2_X1 _10146_ (.A(_03885_),
    .B(_03886_),
    .S(_03504_),
    .Z(_03887_));
 MUX2_X1 _10147_ (.A(\registers[24][25] ),
    .B(\registers[26][25] ),
    .S(_03547_),
    .Z(_03888_));
 MUX2_X1 _10148_ (.A(\registers[25][25] ),
    .B(\registers[27][25] ),
    .S(_03549_),
    .Z(_03889_));
 MUX2_X1 _10149_ (.A(_03888_),
    .B(_03889_),
    .S(_03508_),
    .Z(_03890_));
 MUX2_X1 _10150_ (.A(_03887_),
    .B(_03890_),
    .S(_03629_),
    .Z(_03891_));
 MUX2_X1 _10151_ (.A(\registers[16][25] ),
    .B(\registers[17][25] ),
    .S(_03590_),
    .Z(_03892_));
 NOR2_X1 _10152_ (.A1(_03264_),
    .A2(_03892_),
    .ZN(_03893_));
 MUX2_X1 _10153_ (.A(\registers[18][25] ),
    .B(\registers[19][25] ),
    .S(_03555_),
    .Z(_03894_));
 NOR3_X1 _10154_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_03894_),
    .ZN(_03895_));
 MUX2_X1 _10155_ (.A(\registers[20][25] ),
    .B(\registers[21][25] ),
    .S(_03354_),
    .Z(_03896_));
 NOR3_X1 _10156_ (.A1(_03271_),
    .A2(_03706_),
    .A3(_03896_),
    .ZN(_03897_));
 MUX2_X1 _10157_ (.A(\registers[22][25] ),
    .B(\registers[23][25] ),
    .S(_03517_),
    .Z(_03898_));
 NOR2_X1 _10158_ (.A1(_03275_),
    .A2(_03898_),
    .ZN(_03899_));
 NOR4_X1 _10159_ (.A1(_03893_),
    .A2(_03895_),
    .A3(_03897_),
    .A4(_03899_),
    .ZN(_03900_));
 OAI221_X1 _10160_ (.A(_03622_),
    .B1(_03733_),
    .B2(_03891_),
    .C1(_03900_),
    .C2(_03750_),
    .ZN(_03901_));
 OAI22_X1 _10161_ (.A1(_03865_),
    .A2(_03642_),
    .B1(_03884_),
    .B2(_03901_),
    .ZN(_00378_));
 INV_X1 _10162_ (.A(net55),
    .ZN(_03902_));
 MUX2_X1 _10163_ (.A(\registers[16][26] ),
    .B(\registers[17][26] ),
    .S(_03866_),
    .Z(_03903_));
 MUX2_X1 _10164_ (.A(\registers[22][26] ),
    .B(\registers[23][26] ),
    .S(_03791_),
    .Z(_03904_));
 OAI22_X1 _10165_ (.A1(_03789_),
    .A2(_03903_),
    .B1(_03904_),
    .B2(_03793_),
    .ZN(_03905_));
 MUX2_X1 _10166_ (.A(\registers[18][26] ),
    .B(\registers[19][26] ),
    .S(_03795_),
    .Z(_03906_));
 INV_X1 _10167_ (.A(_03906_),
    .ZN(_03907_));
 AOI21_X1 _10168_ (.A(_03905_),
    .B1(_03907_),
    .B2(_03607_),
    .ZN(_03908_));
 BUF_X4 _10169_ (.A(_03139_),
    .Z(_03909_));
 MUX2_X1 _10170_ (.A(\registers[20][26] ),
    .B(\registers[21][26] ),
    .S(_03909_),
    .Z(_03910_));
 INV_X1 _10171_ (.A(_03910_),
    .ZN(_03911_));
 AOI21_X1 _10172_ (.A(_03721_),
    .B1(_03609_),
    .B2(_03911_),
    .ZN(_03912_));
 MUX2_X1 _10173_ (.A(\registers[28][26] ),
    .B(\registers[30][26] ),
    .S(_03762_),
    .Z(_03913_));
 MUX2_X1 _10174_ (.A(\registers[29][26] ),
    .B(\registers[31][26] ),
    .S(_03803_),
    .Z(_03914_));
 BUF_X4 _10175_ (.A(_03148_),
    .Z(_03915_));
 MUX2_X1 _10176_ (.A(_03913_),
    .B(_03914_),
    .S(_03915_),
    .Z(_03916_));
 MUX2_X1 _10177_ (.A(\registers[24][26] ),
    .B(\registers[26][26] ),
    .S(_03841_),
    .Z(_03917_));
 MUX2_X1 _10178_ (.A(\registers[25][26] ),
    .B(\registers[27][26] ),
    .S(_03880_),
    .Z(_03918_));
 MUX2_X1 _10179_ (.A(_03917_),
    .B(_03918_),
    .S(_03579_),
    .Z(_03919_));
 MUX2_X1 _10180_ (.A(_03916_),
    .B(_03919_),
    .S(_03845_),
    .Z(_03920_));
 AOI221_X1 _10181_ (.A(_03131_),
    .B1(_03908_),
    .B2(_03912_),
    .C1(_03920_),
    .C2(_03620_),
    .ZN(_03921_));
 MUX2_X1 _10182_ (.A(\registers[0][26] ),
    .B(\registers[1][26] ),
    .S(_03319_),
    .Z(_03922_));
 NOR2_X1 _10183_ (.A1(_03184_),
    .A2(_03922_),
    .ZN(_03923_));
 MUX2_X1 _10184_ (.A(\registers[2][26] ),
    .B(\registers[3][26] ),
    .S(_03163_),
    .Z(_03924_));
 NOR3_X1 _10185_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_03924_),
    .ZN(_03925_));
 MUX2_X1 _10186_ (.A(\registers[4][26] ),
    .B(\registers[5][26] ),
    .S(_03386_),
    .Z(_03926_));
 NOR3_X1 _10187_ (.A1(_03193_),
    .A2(_03258_),
    .A3(_03926_),
    .ZN(_03927_));
 MUX2_X1 _10188_ (.A(\registers[6][26] ),
    .B(\registers[7][26] ),
    .S(_03223_),
    .Z(_03928_));
 NOR2_X1 _10189_ (.A1(_03197_),
    .A2(_03928_),
    .ZN(_03929_));
 NOR4_X2 _10190_ (.A1(_03923_),
    .A2(_03925_),
    .A3(_03927_),
    .A4(_03929_),
    .ZN(_03930_));
 MUX2_X1 _10191_ (.A(\registers[12][26] ),
    .B(\registers[14][26] ),
    .S(_03392_),
    .Z(_03931_));
 MUX2_X1 _10192_ (.A(\registers[13][26] ),
    .B(\registers[15][26] ),
    .S(_03394_),
    .Z(_03932_));
 MUX2_X1 _10193_ (.A(_03931_),
    .B(_03932_),
    .S(_03396_),
    .Z(_03933_));
 MUX2_X1 _10194_ (.A(\registers[8][26] ),
    .B(\registers[10][26] ),
    .S(_03398_),
    .Z(_03934_));
 MUX2_X1 _10195_ (.A(\registers[9][26] ),
    .B(\registers[11][26] ),
    .S(_03400_),
    .Z(_03935_));
 MUX2_X1 _10196_ (.A(_03934_),
    .B(_03935_),
    .S(_03203_),
    .Z(_03936_));
 MUX2_X2 _10197_ (.A(_03933_),
    .B(_03936_),
    .S(_03208_),
    .Z(_03937_));
 OAI221_X2 _10198_ (.A(_03622_),
    .B1(_03183_),
    .B2(_03930_),
    .C1(_03937_),
    .C2(_03211_),
    .ZN(_03938_));
 OAI22_X1 _10199_ (.A1(_03902_),
    .A2(_03642_),
    .B1(_03921_),
    .B2(_03938_),
    .ZN(_00379_));
 INV_X1 _10200_ (.A(net56),
    .ZN(_03939_));
 MUX2_X1 _10201_ (.A(\registers[0][27] ),
    .B(\registers[1][27] ),
    .S(_03866_),
    .Z(_03940_));
 MUX2_X1 _10202_ (.A(\registers[6][27] ),
    .B(\registers[7][27] ),
    .S(_03791_),
    .Z(_03941_));
 OAI22_X1 _10203_ (.A1(_03789_),
    .A2(_03940_),
    .B1(_03941_),
    .B2(_03793_),
    .ZN(_03942_));
 MUX2_X1 _10204_ (.A(\registers[2][27] ),
    .B(\registers[3][27] ),
    .S(_03795_),
    .Z(_03943_));
 INV_X1 _10205_ (.A(_03943_),
    .ZN(_03944_));
 AOI21_X1 _10206_ (.A(_03942_),
    .B1(_03944_),
    .B2(_03607_),
    .ZN(_03945_));
 MUX2_X1 _10207_ (.A(\registers[4][27] ),
    .B(\registers[5][27] ),
    .S(_03909_),
    .Z(_03946_));
 INV_X1 _10208_ (.A(_03946_),
    .ZN(_03947_));
 AOI21_X1 _10209_ (.A(_03721_),
    .B1(_03609_),
    .B2(_03947_),
    .ZN(_03948_));
 MUX2_X1 _10210_ (.A(\registers[12][27] ),
    .B(\registers[14][27] ),
    .S(_03762_),
    .Z(_03949_));
 MUX2_X1 _10211_ (.A(\registers[13][27] ),
    .B(\registers[15][27] ),
    .S(_03803_),
    .Z(_03950_));
 MUX2_X1 _10212_ (.A(_03949_),
    .B(_03950_),
    .S(_03915_),
    .Z(_03951_));
 MUX2_X1 _10213_ (.A(\registers[8][27] ),
    .B(\registers[10][27] ),
    .S(_03841_),
    .Z(_03952_));
 MUX2_X1 _10214_ (.A(\registers[9][27] ),
    .B(\registers[11][27] ),
    .S(_03880_),
    .Z(_03953_));
 BUF_X4 _10215_ (.A(_03148_),
    .Z(_03954_));
 MUX2_X1 _10216_ (.A(_03952_),
    .B(_03953_),
    .S(_03954_),
    .Z(_03955_));
 MUX2_X2 _10217_ (.A(_03951_),
    .B(_03955_),
    .S(_03845_),
    .Z(_03956_));
 AOI221_X2 _10218_ (.A(_03714_),
    .B1(_03945_),
    .B2(_03948_),
    .C1(_03956_),
    .C2(_03620_),
    .ZN(_03957_));
 MUX2_X1 _10219_ (.A(\registers[28][27] ),
    .B(\registers[30][27] ),
    .S(_03542_),
    .Z(_03958_));
 MUX2_X1 _10220_ (.A(\registers[29][27] ),
    .B(\registers[31][27] ),
    .S(_03544_),
    .Z(_03959_));
 MUX2_X1 _10221_ (.A(_03958_),
    .B(_03959_),
    .S(_03504_),
    .Z(_03960_));
 MUX2_X1 _10222_ (.A(\registers[24][27] ),
    .B(\registers[26][27] ),
    .S(_03547_),
    .Z(_03961_));
 MUX2_X1 _10223_ (.A(\registers[25][27] ),
    .B(\registers[27][27] ),
    .S(_03549_),
    .Z(_03962_));
 MUX2_X1 _10224_ (.A(_03961_),
    .B(_03962_),
    .S(_03508_),
    .Z(_03963_));
 MUX2_X1 _10225_ (.A(_03960_),
    .B(_03963_),
    .S(_03629_),
    .Z(_03964_));
 MUX2_X1 _10226_ (.A(\registers[16][27] ),
    .B(\registers[17][27] ),
    .S(_03590_),
    .Z(_03965_));
 NOR2_X1 _10227_ (.A1(_03264_),
    .A2(_03965_),
    .ZN(_03966_));
 MUX2_X1 _10228_ (.A(\registers[18][27] ),
    .B(\registers[19][27] ),
    .S(_03555_),
    .Z(_03967_));
 NOR3_X1 _10229_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_03967_),
    .ZN(_03968_));
 MUX2_X1 _10230_ (.A(\registers[20][27] ),
    .B(\registers[21][27] ),
    .S(_03149_),
    .Z(_03969_));
 NOR3_X1 _10231_ (.A1(_03271_),
    .A2(_03706_),
    .A3(_03969_),
    .ZN(_03970_));
 MUX2_X1 _10232_ (.A(\registers[22][27] ),
    .B(\registers[23][27] ),
    .S(_03517_),
    .Z(_03971_));
 NOR2_X1 _10233_ (.A1(_03275_),
    .A2(_03971_),
    .ZN(_03972_));
 NOR4_X2 _10234_ (.A1(_03966_),
    .A2(_03968_),
    .A3(_03970_),
    .A4(_03972_),
    .ZN(_03973_));
 OAI221_X1 _10235_ (.A(_03622_),
    .B1(_03733_),
    .B2(_03964_),
    .C1(_03973_),
    .C2(_03750_),
    .ZN(_03974_));
 OAI22_X1 _10236_ (.A1(_03939_),
    .A2(_03642_),
    .B1(_03957_),
    .B2(_03974_),
    .ZN(_00380_));
 INV_X1 _10237_ (.A(net57),
    .ZN(_03975_));
 MUX2_X1 _10238_ (.A(\registers[16][28] ),
    .B(\registers[17][28] ),
    .S(_03866_),
    .Z(_03976_));
 MUX2_X1 _10239_ (.A(\registers[22][28] ),
    .B(\registers[23][28] ),
    .S(_03791_),
    .Z(_03977_));
 OAI22_X2 _10240_ (.A1(_03789_),
    .A2(_03976_),
    .B1(_03977_),
    .B2(_03793_),
    .ZN(_03978_));
 MUX2_X1 _10241_ (.A(\registers[18][28] ),
    .B(\registers[19][28] ),
    .S(_03795_),
    .Z(_03979_));
 INV_X1 _10242_ (.A(_03979_),
    .ZN(_03980_));
 BUF_X4 _10243_ (.A(_03154_),
    .Z(_03981_));
 AOI21_X2 _10244_ (.A(_03978_),
    .B1(_03980_),
    .B2(_03981_),
    .ZN(_03982_));
 CLKBUF_X3 _10245_ (.A(_03161_),
    .Z(_03983_));
 MUX2_X1 _10246_ (.A(\registers[20][28] ),
    .B(\registers[21][28] ),
    .S(_03909_),
    .Z(_03984_));
 INV_X1 _10247_ (.A(_03984_),
    .ZN(_03985_));
 AOI21_X1 _10248_ (.A(_03721_),
    .B1(_03983_),
    .B2(_03985_),
    .ZN(_03986_));
 MUX2_X1 _10249_ (.A(\registers[28][28] ),
    .B(\registers[30][28] ),
    .S(_03762_),
    .Z(_03987_));
 MUX2_X1 _10250_ (.A(\registers[29][28] ),
    .B(\registers[31][28] ),
    .S(_03803_),
    .Z(_03988_));
 MUX2_X1 _10251_ (.A(_03987_),
    .B(_03988_),
    .S(_03915_),
    .Z(_03989_));
 MUX2_X1 _10252_ (.A(\registers[24][28] ),
    .B(\registers[26][28] ),
    .S(_03841_),
    .Z(_03990_));
 MUX2_X1 _10253_ (.A(\registers[25][28] ),
    .B(\registers[27][28] ),
    .S(_03880_),
    .Z(_03991_));
 MUX2_X1 _10254_ (.A(_03990_),
    .B(_03991_),
    .S(_03954_),
    .Z(_03992_));
 MUX2_X1 _10255_ (.A(_03989_),
    .B(_03992_),
    .S(_03845_),
    .Z(_03993_));
 BUF_X4 _10256_ (.A(_03158_),
    .Z(_03994_));
 AOI221_X2 _10257_ (.A(_03131_),
    .B1(_03982_),
    .B2(_03986_),
    .C1(_03993_),
    .C2(_03994_),
    .ZN(_03995_));
 BUF_X4 _10258_ (.A(_03180_),
    .Z(_03996_));
 MUX2_X1 _10259_ (.A(\registers[0][28] ),
    .B(\registers[1][28] ),
    .S(_03319_),
    .Z(_03997_));
 NOR2_X1 _10260_ (.A1(_03184_),
    .A2(_03997_),
    .ZN(_03998_));
 MUX2_X1 _10261_ (.A(\registers[2][28] ),
    .B(\registers[3][28] ),
    .S(_03163_),
    .Z(_03999_));
 NOR3_X1 _10262_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_03999_),
    .ZN(_04000_));
 MUX2_X1 _10263_ (.A(\registers[4][28] ),
    .B(\registers[5][28] ),
    .S(_03386_),
    .Z(_04001_));
 NOR3_X1 _10264_ (.A1(_03193_),
    .A2(_03258_),
    .A3(_04001_),
    .ZN(_04002_));
 MUX2_X1 _10265_ (.A(\registers[6][28] ),
    .B(\registers[7][28] ),
    .S(_03223_),
    .Z(_04003_));
 NOR2_X1 _10266_ (.A1(_03197_),
    .A2(_04003_),
    .ZN(_04004_));
 NOR4_X2 _10267_ (.A1(_03998_),
    .A2(_04000_),
    .A3(_04002_),
    .A4(_04004_),
    .ZN(_04005_));
 MUX2_X1 _10268_ (.A(\registers[12][28] ),
    .B(\registers[14][28] ),
    .S(_03392_),
    .Z(_04006_));
 MUX2_X1 _10269_ (.A(\registers[13][28] ),
    .B(\registers[15][28] ),
    .S(_03394_),
    .Z(_04007_));
 MUX2_X1 _10270_ (.A(_04006_),
    .B(_04007_),
    .S(_03396_),
    .Z(_04008_));
 MUX2_X1 _10271_ (.A(\registers[8][28] ),
    .B(\registers[10][28] ),
    .S(_03398_),
    .Z(_04009_));
 MUX2_X1 _10272_ (.A(\registers[9][28] ),
    .B(\registers[11][28] ),
    .S(_03400_),
    .Z(_04010_));
 MUX2_X1 _10273_ (.A(_04009_),
    .B(_04010_),
    .S(_03203_),
    .Z(_04011_));
 MUX2_X2 _10274_ (.A(_04008_),
    .B(_04011_),
    .S(_03208_),
    .Z(_04012_));
 OAI221_X2 _10275_ (.A(_03996_),
    .B1(_03183_),
    .B2(_04005_),
    .C1(_04012_),
    .C2(_03211_),
    .ZN(_04013_));
 OAI22_X1 _10276_ (.A1(_03975_),
    .A2(_03642_),
    .B1(_03995_),
    .B2(_04013_),
    .ZN(_00381_));
 INV_X1 _10277_ (.A(net58),
    .ZN(_04014_));
 CLKBUF_X3 _10278_ (.A(_03214_),
    .Z(_04015_));
 MUX2_X1 _10279_ (.A(\registers[0][29] ),
    .B(\registers[1][29] ),
    .S(_03866_),
    .Z(_04016_));
 MUX2_X1 _10280_ (.A(\registers[6][29] ),
    .B(\registers[7][29] ),
    .S(_03791_),
    .Z(_04017_));
 OAI22_X1 _10281_ (.A1(_03789_),
    .A2(_04016_),
    .B1(_04017_),
    .B2(_03793_),
    .ZN(_04018_));
 MUX2_X1 _10282_ (.A(\registers[2][29] ),
    .B(\registers[3][29] ),
    .S(_03795_),
    .Z(_04019_));
 INV_X1 _10283_ (.A(_04019_),
    .ZN(_04020_));
 AOI21_X1 _10284_ (.A(_04018_),
    .B1(_04020_),
    .B2(_03981_),
    .ZN(_04021_));
 MUX2_X1 _10285_ (.A(\registers[4][29] ),
    .B(\registers[5][29] ),
    .S(_03909_),
    .Z(_04022_));
 INV_X1 _10286_ (.A(_04022_),
    .ZN(_04023_));
 AOI21_X1 _10287_ (.A(_03721_),
    .B1(_03983_),
    .B2(_04023_),
    .ZN(_04024_));
 MUX2_X1 _10288_ (.A(\registers[12][29] ),
    .B(\registers[14][29] ),
    .S(_03762_),
    .Z(_04025_));
 MUX2_X1 _10289_ (.A(\registers[13][29] ),
    .B(\registers[15][29] ),
    .S(_03803_),
    .Z(_04026_));
 MUX2_X1 _10290_ (.A(_04025_),
    .B(_04026_),
    .S(_03915_),
    .Z(_04027_));
 MUX2_X1 _10291_ (.A(\registers[8][29] ),
    .B(\registers[10][29] ),
    .S(_03841_),
    .Z(_04028_));
 MUX2_X1 _10292_ (.A(\registers[9][29] ),
    .B(\registers[11][29] ),
    .S(_03880_),
    .Z(_04029_));
 MUX2_X1 _10293_ (.A(_04028_),
    .B(_04029_),
    .S(_03954_),
    .Z(_04030_));
 MUX2_X2 _10294_ (.A(_04027_),
    .B(_04030_),
    .S(_03845_),
    .Z(_04031_));
 AOI221_X2 _10295_ (.A(_03714_),
    .B1(_04021_),
    .B2(_04024_),
    .C1(_04031_),
    .C2(_03994_),
    .ZN(_04032_));
 MUX2_X1 _10296_ (.A(\registers[28][29] ),
    .B(\registers[30][29] ),
    .S(_03542_),
    .Z(_04033_));
 MUX2_X1 _10297_ (.A(\registers[29][29] ),
    .B(\registers[31][29] ),
    .S(_03544_),
    .Z(_04034_));
 MUX2_X1 _10298_ (.A(_04033_),
    .B(_04034_),
    .S(_03504_),
    .Z(_04035_));
 MUX2_X1 _10299_ (.A(\registers[24][29] ),
    .B(\registers[26][29] ),
    .S(_03547_),
    .Z(_04036_));
 MUX2_X1 _10300_ (.A(\registers[25][29] ),
    .B(\registers[27][29] ),
    .S(_03549_),
    .Z(_04037_));
 MUX2_X1 _10301_ (.A(_04036_),
    .B(_04037_),
    .S(_03508_),
    .Z(_04038_));
 MUX2_X1 _10302_ (.A(_04035_),
    .B(_04038_),
    .S(_03629_),
    .Z(_04039_));
 MUX2_X1 _10303_ (.A(\registers[16][29] ),
    .B(\registers[17][29] ),
    .S(_03590_),
    .Z(_04040_));
 NOR2_X1 _10304_ (.A1(_03264_),
    .A2(_04040_),
    .ZN(_04041_));
 MUX2_X1 _10305_ (.A(\registers[18][29] ),
    .B(\registers[19][29] ),
    .S(_03555_),
    .Z(_04042_));
 NOR3_X1 _10306_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_04042_),
    .ZN(_04043_));
 MUX2_X1 _10307_ (.A(\registers[20][29] ),
    .B(\registers[21][29] ),
    .S(_03149_),
    .Z(_04044_));
 NOR3_X1 _10308_ (.A1(_03271_),
    .A2(_03706_),
    .A3(_04044_),
    .ZN(_04045_));
 MUX2_X1 _10309_ (.A(\registers[22][29] ),
    .B(\registers[23][29] ),
    .S(_03517_),
    .Z(_04046_));
 NOR2_X1 _10310_ (.A1(_03275_),
    .A2(_04046_),
    .ZN(_04047_));
 NOR4_X1 _10311_ (.A1(_04041_),
    .A2(_04043_),
    .A3(_04045_),
    .A4(_04047_),
    .ZN(_04048_));
 OAI221_X1 _10312_ (.A(_03996_),
    .B1(_03733_),
    .B2(_04039_),
    .C1(_04048_),
    .C2(_03750_),
    .ZN(_04049_));
 OAI22_X1 _10313_ (.A1(_04014_),
    .A2(_04015_),
    .B1(_04032_),
    .B2(_04049_),
    .ZN(_00382_));
 INV_X1 _10314_ (.A(net59),
    .ZN(_04050_));
 MUX2_X1 _10315_ (.A(\registers[16][2] ),
    .B(\registers[17][2] ),
    .S(_03866_),
    .Z(_04051_));
 MUX2_X1 _10316_ (.A(\registers[22][2] ),
    .B(\registers[23][2] ),
    .S(_03791_),
    .Z(_04052_));
 OAI22_X2 _10317_ (.A1(_03789_),
    .A2(_04051_),
    .B1(_04052_),
    .B2(_03793_),
    .ZN(_04053_));
 MUX2_X1 _10318_ (.A(\registers[18][2] ),
    .B(\registers[19][2] ),
    .S(_03795_),
    .Z(_04054_));
 INV_X1 _10319_ (.A(_04054_),
    .ZN(_04055_));
 AOI21_X2 _10320_ (.A(_04053_),
    .B1(_04055_),
    .B2(_03981_),
    .ZN(_04056_));
 MUX2_X1 _10321_ (.A(\registers[20][2] ),
    .B(\registers[21][2] ),
    .S(_03909_),
    .Z(_04057_));
 INV_X1 _10322_ (.A(_04057_),
    .ZN(_04058_));
 AOI21_X1 _10323_ (.A(_03721_),
    .B1(_03983_),
    .B2(_04058_),
    .ZN(_04059_));
 MUX2_X1 _10324_ (.A(\registers[28][2] ),
    .B(\registers[30][2] ),
    .S(_03762_),
    .Z(_04060_));
 MUX2_X1 _10325_ (.A(\registers[29][2] ),
    .B(\registers[31][2] ),
    .S(_03803_),
    .Z(_04061_));
 MUX2_X1 _10326_ (.A(_04060_),
    .B(_04061_),
    .S(_03915_),
    .Z(_04062_));
 MUX2_X1 _10327_ (.A(\registers[24][2] ),
    .B(\registers[26][2] ),
    .S(_03841_),
    .Z(_04063_));
 MUX2_X1 _10328_ (.A(\registers[25][2] ),
    .B(\registers[27][2] ),
    .S(_03880_),
    .Z(_04064_));
 MUX2_X1 _10329_ (.A(_04063_),
    .B(_04064_),
    .S(_03954_),
    .Z(_04065_));
 MUX2_X2 _10330_ (.A(_04062_),
    .B(_04065_),
    .S(_03845_),
    .Z(_04066_));
 AOI221_X2 _10331_ (.A(_03131_),
    .B1(_04056_),
    .B2(_04059_),
    .C1(_04066_),
    .C2(_03994_),
    .ZN(_04067_));
 MUX2_X1 _10332_ (.A(\registers[0][2] ),
    .B(\registers[1][2] ),
    .S(_03319_),
    .Z(_04068_));
 NOR2_X1 _10333_ (.A1(_03184_),
    .A2(_04068_),
    .ZN(_04069_));
 MUX2_X1 _10334_ (.A(\registers[2][2] ),
    .B(\registers[3][2] ),
    .S(_03163_),
    .Z(_04070_));
 NOR3_X1 _10335_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_04070_),
    .ZN(_04071_));
 MUX2_X1 _10336_ (.A(\registers[4][2] ),
    .B(\registers[5][2] ),
    .S(_03386_),
    .Z(_04072_));
 NOR3_X1 _10337_ (.A1(_03193_),
    .A2(_03258_),
    .A3(_04072_),
    .ZN(_04073_));
 MUX2_X1 _10338_ (.A(\registers[6][2] ),
    .B(\registers[7][2] ),
    .S(_03223_),
    .Z(_04074_));
 NOR2_X1 _10339_ (.A1(_03197_),
    .A2(_04074_),
    .ZN(_04075_));
 NOR4_X2 _10340_ (.A1(_04069_),
    .A2(_04071_),
    .A3(_04073_),
    .A4(_04075_),
    .ZN(_04076_));
 MUX2_X1 _10341_ (.A(\registers[12][2] ),
    .B(\registers[14][2] ),
    .S(_03255_),
    .Z(_04077_));
 MUX2_X1 _10342_ (.A(\registers[13][2] ),
    .B(\registers[15][2] ),
    .S(_03394_),
    .Z(_04078_));
 MUX2_X1 _10343_ (.A(_04077_),
    .B(_04078_),
    .S(_03306_),
    .Z(_04079_));
 MUX2_X1 _10344_ (.A(\registers[8][2] ),
    .B(\registers[10][2] ),
    .S(_03398_),
    .Z(_04080_));
 MUX2_X1 _10345_ (.A(\registers[9][2] ),
    .B(\registers[11][2] ),
    .S(_03400_),
    .Z(_04081_));
 MUX2_X1 _10346_ (.A(_04080_),
    .B(_04081_),
    .S(_03203_),
    .Z(_04082_));
 MUX2_X2 _10347_ (.A(_04079_),
    .B(_04082_),
    .S(_03208_),
    .Z(_04083_));
 OAI221_X2 _10348_ (.A(_03996_),
    .B1(_03183_),
    .B2(_04076_),
    .C1(_04083_),
    .C2(_03211_),
    .ZN(_04084_));
 OAI22_X1 _10349_ (.A1(_04050_),
    .A2(_04015_),
    .B1(_04067_),
    .B2(_04084_),
    .ZN(_00383_));
 INV_X1 _10350_ (.A(net60),
    .ZN(_04085_));
 MUX2_X1 _10351_ (.A(\registers[0][30] ),
    .B(\registers[1][30] ),
    .S(_03866_),
    .Z(_04086_));
 MUX2_X1 _10352_ (.A(\registers[6][30] ),
    .B(\registers[7][30] ),
    .S(_03791_),
    .Z(_04087_));
 OAI22_X1 _10353_ (.A1(_03789_),
    .A2(_04086_),
    .B1(_04087_),
    .B2(_03793_),
    .ZN(_04088_));
 MUX2_X1 _10354_ (.A(\registers[2][30] ),
    .B(\registers[3][30] ),
    .S(_03795_),
    .Z(_04089_));
 INV_X1 _10355_ (.A(_04089_),
    .ZN(_04090_));
 AOI21_X1 _10356_ (.A(_04088_),
    .B1(_04090_),
    .B2(_03981_),
    .ZN(_04091_));
 MUX2_X1 _10357_ (.A(\registers[4][30] ),
    .B(\registers[5][30] ),
    .S(_03909_),
    .Z(_04092_));
 INV_X1 _10358_ (.A(_04092_),
    .ZN(_04093_));
 AOI21_X1 _10359_ (.A(_03261_),
    .B1(_03983_),
    .B2(_04093_),
    .ZN(_04094_));
 MUX2_X1 _10360_ (.A(\registers[12][30] ),
    .B(\registers[14][30] ),
    .S(_03762_),
    .Z(_04095_));
 MUX2_X1 _10361_ (.A(\registers[13][30] ),
    .B(\registers[15][30] ),
    .S(_03803_),
    .Z(_04096_));
 MUX2_X1 _10362_ (.A(_04095_),
    .B(_04096_),
    .S(_03915_),
    .Z(_04097_));
 MUX2_X1 _10363_ (.A(\registers[8][30] ),
    .B(\registers[10][30] ),
    .S(_03841_),
    .Z(_04098_));
 MUX2_X1 _10364_ (.A(\registers[9][30] ),
    .B(\registers[11][30] ),
    .S(_03880_),
    .Z(_04099_));
 MUX2_X1 _10365_ (.A(_04098_),
    .B(_04099_),
    .S(_03954_),
    .Z(_04100_));
 MUX2_X2 _10366_ (.A(_04097_),
    .B(_04100_),
    .S(_03845_),
    .Z(_04101_));
 AOI221_X2 _10367_ (.A(_03714_),
    .B1(_04091_),
    .B2(_04094_),
    .C1(_04101_),
    .C2(_03994_),
    .ZN(_04102_));
 MUX2_X1 _10368_ (.A(\registers[28][30] ),
    .B(\registers[30][30] ),
    .S(_03542_),
    .Z(_04103_));
 MUX2_X1 _10369_ (.A(\registers[29][30] ),
    .B(\registers[31][30] ),
    .S(_03544_),
    .Z(_04104_));
 MUX2_X1 _10370_ (.A(_04103_),
    .B(_04104_),
    .S(_03504_),
    .Z(_04105_));
 MUX2_X1 _10371_ (.A(\registers[24][30] ),
    .B(\registers[26][30] ),
    .S(_03547_),
    .Z(_04106_));
 MUX2_X1 _10372_ (.A(\registers[25][30] ),
    .B(\registers[27][30] ),
    .S(_03549_),
    .Z(_04107_));
 MUX2_X1 _10373_ (.A(_04106_),
    .B(_04107_),
    .S(_03508_),
    .Z(_04108_));
 MUX2_X1 _10374_ (.A(_04105_),
    .B(_04108_),
    .S(_03629_),
    .Z(_04109_));
 MUX2_X1 _10375_ (.A(\registers[16][30] ),
    .B(\registers[17][30] ),
    .S(_03590_),
    .Z(_04110_));
 NOR2_X1 _10376_ (.A1(_03264_),
    .A2(_04110_),
    .ZN(_04111_));
 MUX2_X1 _10377_ (.A(\registers[18][30] ),
    .B(\registers[19][30] ),
    .S(_03555_),
    .Z(_04112_));
 NOR3_X1 _10378_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_04112_),
    .ZN(_04113_));
 MUX2_X1 _10379_ (.A(\registers[20][30] ),
    .B(\registers[21][30] ),
    .S(_03149_),
    .Z(_04114_));
 NOR3_X1 _10380_ (.A1(_03271_),
    .A2(_03706_),
    .A3(_04114_),
    .ZN(_04115_));
 MUX2_X1 _10381_ (.A(\registers[22][30] ),
    .B(\registers[23][30] ),
    .S(_03517_),
    .Z(_04116_));
 NOR2_X1 _10382_ (.A1(_03275_),
    .A2(_04116_),
    .ZN(_04117_));
 NOR4_X2 _10383_ (.A1(_04111_),
    .A2(_04113_),
    .A3(_04115_),
    .A4(_04117_),
    .ZN(_04118_));
 OAI221_X1 _10384_ (.A(_03996_),
    .B1(_03733_),
    .B2(_04109_),
    .C1(_04118_),
    .C2(_03750_),
    .ZN(_04119_));
 OAI22_X1 _10385_ (.A1(_04085_),
    .A2(_04015_),
    .B1(_04102_),
    .B2(_04119_),
    .ZN(_00384_));
 INV_X1 _10386_ (.A(net61),
    .ZN(_04120_));
 MUX2_X1 _10387_ (.A(\registers[16][31] ),
    .B(\registers[17][31] ),
    .S(_03866_),
    .Z(_04121_));
 MUX2_X1 _10388_ (.A(\registers[22][31] ),
    .B(\registers[23][31] ),
    .S(_03791_),
    .Z(_04122_));
 OAI22_X2 _10389_ (.A1(_03789_),
    .A2(_04121_),
    .B1(_04122_),
    .B2(_03793_),
    .ZN(_04123_));
 MUX2_X1 _10390_ (.A(\registers[18][31] ),
    .B(\registers[19][31] ),
    .S(_03795_),
    .Z(_04124_));
 INV_X1 _10391_ (.A(_04124_),
    .ZN(_04125_));
 AOI21_X2 _10392_ (.A(_04123_),
    .B1(_04125_),
    .B2(_03981_),
    .ZN(_04126_));
 MUX2_X1 _10393_ (.A(\registers[20][31] ),
    .B(\registers[21][31] ),
    .S(_03909_),
    .Z(_04127_));
 INV_X1 _10394_ (.A(_04127_),
    .ZN(_04128_));
 AOI21_X1 _10395_ (.A(_03261_),
    .B1(_03983_),
    .B2(_04128_),
    .ZN(_04129_));
 MUX2_X1 _10396_ (.A(\registers[28][31] ),
    .B(\registers[30][31] ),
    .S(_03142_),
    .Z(_04130_));
 MUX2_X1 _10397_ (.A(\registers[29][31] ),
    .B(\registers[31][31] ),
    .S(_03803_),
    .Z(_04131_));
 MUX2_X1 _10398_ (.A(_04130_),
    .B(_04131_),
    .S(_03915_),
    .Z(_04132_));
 MUX2_X1 _10399_ (.A(\registers[24][31] ),
    .B(\registers[26][31] ),
    .S(_03841_),
    .Z(_04133_));
 MUX2_X1 _10400_ (.A(\registers[25][31] ),
    .B(\registers[27][31] ),
    .S(_03880_),
    .Z(_04134_));
 MUX2_X1 _10401_ (.A(_04133_),
    .B(_04134_),
    .S(_03954_),
    .Z(_04135_));
 MUX2_X1 _10402_ (.A(_04132_),
    .B(_04135_),
    .S(_03845_),
    .Z(_04136_));
 AOI221_X2 _10403_ (.A(_03131_),
    .B1(_04126_),
    .B2(_04129_),
    .C1(_04136_),
    .C2(_03994_),
    .ZN(_04137_));
 MUX2_X1 _10404_ (.A(\registers[0][31] ),
    .B(\registers[1][31] ),
    .S(_03319_),
    .Z(_04138_));
 NOR2_X1 _10405_ (.A1(_03184_),
    .A2(_04138_),
    .ZN(_04139_));
 MUX2_X1 _10406_ (.A(\registers[2][31] ),
    .B(\registers[3][31] ),
    .S(_03163_),
    .Z(_04140_));
 NOR3_X1 _10407_ (.A1(_03188_),
    .A2(_03189_),
    .A3(_04140_),
    .ZN(_04141_));
 MUX2_X1 _10408_ (.A(\registers[4][31] ),
    .B(\registers[5][31] ),
    .S(_03227_),
    .Z(_04142_));
 NOR3_X1 _10409_ (.A1(_03193_),
    .A2(_03258_),
    .A3(_04142_),
    .ZN(_04143_));
 MUX2_X1 _10410_ (.A(\registers[6][31] ),
    .B(\registers[7][31] ),
    .S(_03223_),
    .Z(_04144_));
 NOR2_X1 _10411_ (.A1(_03197_),
    .A2(_04144_),
    .ZN(_04145_));
 NOR4_X2 _10412_ (.A1(_04139_),
    .A2(_04141_),
    .A3(_04143_),
    .A4(_04145_),
    .ZN(_04146_));
 MUX2_X1 _10413_ (.A(\registers[12][31] ),
    .B(\registers[14][31] ),
    .S(_03255_),
    .Z(_04147_));
 MUX2_X1 _10414_ (.A(\registers[13][31] ),
    .B(\registers[15][31] ),
    .S(_03392_),
    .Z(_04148_));
 MUX2_X1 _10415_ (.A(_04147_),
    .B(_04148_),
    .S(_03306_),
    .Z(_04149_));
 MUX2_X1 _10416_ (.A(\registers[8][31] ),
    .B(\registers[10][31] ),
    .S(_03398_),
    .Z(_04150_));
 MUX2_X1 _10417_ (.A(\registers[9][31] ),
    .B(\registers[11][31] ),
    .S(_03400_),
    .Z(_04151_));
 MUX2_X1 _10418_ (.A(_04150_),
    .B(_04151_),
    .S(_03396_),
    .Z(_04152_));
 MUX2_X1 _10419_ (.A(_04149_),
    .B(_04152_),
    .S(_03208_),
    .Z(_04153_));
 OAI221_X2 _10420_ (.A(_03996_),
    .B1(_03183_),
    .B2(_04146_),
    .C1(_04153_),
    .C2(_03211_),
    .ZN(_04154_));
 OAI22_X1 _10421_ (.A1(_04120_),
    .A2(_04015_),
    .B1(_04137_),
    .B2(_04154_),
    .ZN(_00385_));
 INV_X1 _10422_ (.A(net62),
    .ZN(_04155_));
 MUX2_X1 _10423_ (.A(\registers[0][3] ),
    .B(\registers[1][3] ),
    .S(_03866_),
    .Z(_04156_));
 MUX2_X1 _10424_ (.A(\registers[6][3] ),
    .B(\registers[7][3] ),
    .S(_03169_),
    .Z(_04157_));
 OAI22_X1 _10425_ (.A1(_03136_),
    .A2(_04156_),
    .B1(_04157_),
    .B2(_03143_),
    .ZN(_04158_));
 MUX2_X1 _10426_ (.A(\registers[2][3] ),
    .B(\registers[3][3] ),
    .S(_03194_),
    .Z(_04159_));
 INV_X1 _10427_ (.A(_04159_),
    .ZN(_04160_));
 AOI21_X1 _10428_ (.A(_04158_),
    .B1(_04160_),
    .B2(_03981_),
    .ZN(_04161_));
 MUX2_X1 _10429_ (.A(\registers[4][3] ),
    .B(\registers[5][3] ),
    .S(_03909_),
    .Z(_04162_));
 INV_X1 _10430_ (.A(_04162_),
    .ZN(_04163_));
 AOI21_X1 _10431_ (.A(_03261_),
    .B1(_03983_),
    .B2(_04163_),
    .ZN(_04164_));
 MUX2_X1 _10432_ (.A(\registers[12][3] ),
    .B(\registers[14][3] ),
    .S(_03142_),
    .Z(_04165_));
 MUX2_X1 _10433_ (.A(\registers[13][3] ),
    .B(\registers[15][3] ),
    .S(_03232_),
    .Z(_04166_));
 MUX2_X1 _10434_ (.A(_04165_),
    .B(_04166_),
    .S(_03915_),
    .Z(_04167_));
 MUX2_X1 _10435_ (.A(\registers[8][3] ),
    .B(\registers[10][3] ),
    .S(_03841_),
    .Z(_04168_));
 MUX2_X1 _10436_ (.A(\registers[9][3] ),
    .B(\registers[11][3] ),
    .S(_03880_),
    .Z(_04169_));
 MUX2_X1 _10437_ (.A(_04168_),
    .B(_04169_),
    .S(_03954_),
    .Z(_04170_));
 MUX2_X2 _10438_ (.A(_04167_),
    .B(_04170_),
    .S(_03845_),
    .Z(_04171_));
 AOI221_X2 _10439_ (.A(_03714_),
    .B1(_04161_),
    .B2(_04164_),
    .C1(_04171_),
    .C2(_03994_),
    .ZN(_04172_));
 MUX2_X1 _10440_ (.A(\registers[28][3] ),
    .B(\registers[30][3] ),
    .S(_03542_),
    .Z(_04173_));
 MUX2_X1 _10441_ (.A(\registers[29][3] ),
    .B(\registers[31][3] ),
    .S(_03544_),
    .Z(_04174_));
 MUX2_X1 _10442_ (.A(_04173_),
    .B(_04174_),
    .S(_03380_),
    .Z(_04175_));
 MUX2_X1 _10443_ (.A(\registers[24][3] ),
    .B(\registers[26][3] ),
    .S(_03547_),
    .Z(_04176_));
 MUX2_X1 _10444_ (.A(\registers[25][3] ),
    .B(\registers[27][3] ),
    .S(_03549_),
    .Z(_04177_));
 MUX2_X1 _10445_ (.A(_04176_),
    .B(_04177_),
    .S(_03251_),
    .Z(_04178_));
 MUX2_X1 _10446_ (.A(_04175_),
    .B(_04178_),
    .S(_03629_),
    .Z(_04179_));
 MUX2_X1 _10447_ (.A(\registers[16][3] ),
    .B(\registers[17][3] ),
    .S(_03590_),
    .Z(_04180_));
 NOR2_X1 _10448_ (.A1(_03264_),
    .A2(_04180_),
    .ZN(_04181_));
 MUX2_X1 _10449_ (.A(\registers[18][3] ),
    .B(\registers[19][3] ),
    .S(_03555_),
    .Z(_04182_));
 NOR3_X1 _10450_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_04182_),
    .ZN(_04183_));
 MUX2_X1 _10451_ (.A(\registers[20][3] ),
    .B(\registers[21][3] ),
    .S(_03149_),
    .Z(_04184_));
 NOR3_X1 _10452_ (.A1(_03271_),
    .A2(_03706_),
    .A3(_04184_),
    .ZN(_04185_));
 MUX2_X1 _10453_ (.A(\registers[22][3] ),
    .B(\registers[23][3] ),
    .S(_03311_),
    .Z(_04186_));
 NOR2_X1 _10454_ (.A1(_03275_),
    .A2(_04186_),
    .ZN(_04187_));
 NOR4_X2 _10455_ (.A1(_04181_),
    .A2(_04183_),
    .A3(_04185_),
    .A4(_04187_),
    .ZN(_04188_));
 OAI221_X1 _10456_ (.A(_03996_),
    .B1(_03733_),
    .B2(_04179_),
    .C1(_04188_),
    .C2(_03750_),
    .ZN(_04189_));
 OAI22_X1 _10457_ (.A1(_04155_),
    .A2(_04015_),
    .B1(_04172_),
    .B2(_04189_),
    .ZN(_00386_));
 INV_X1 _10458_ (.A(net63),
    .ZN(_04190_));
 MUX2_X1 _10459_ (.A(\registers[16][4] ),
    .B(\registers[17][4] ),
    .S(_03866_),
    .Z(_04191_));
 MUX2_X1 _10460_ (.A(\registers[22][4] ),
    .B(\registers[23][4] ),
    .S(_03169_),
    .Z(_04192_));
 OAI22_X1 _10461_ (.A1(_03136_),
    .A2(_04191_),
    .B1(_04192_),
    .B2(_03143_),
    .ZN(_04193_));
 MUX2_X1 _10462_ (.A(\registers[18][4] ),
    .B(\registers[19][4] ),
    .S(_03194_),
    .Z(_04194_));
 INV_X1 _10463_ (.A(_04194_),
    .ZN(_04195_));
 AOI21_X2 _10464_ (.A(_04193_),
    .B1(_04195_),
    .B2(_03981_),
    .ZN(_04196_));
 MUX2_X1 _10465_ (.A(\registers[20][4] ),
    .B(\registers[21][4] ),
    .S(_03909_),
    .Z(_04197_));
 INV_X1 _10466_ (.A(_04197_),
    .ZN(_04198_));
 AOI21_X1 _10467_ (.A(_03261_),
    .B1(_03983_),
    .B2(_04198_),
    .ZN(_04199_));
 MUX2_X1 _10468_ (.A(\registers[28][4] ),
    .B(\registers[30][4] ),
    .S(_03142_),
    .Z(_04200_));
 MUX2_X1 _10469_ (.A(\registers[29][4] ),
    .B(\registers[31][4] ),
    .S(_03232_),
    .Z(_04201_));
 MUX2_X1 _10470_ (.A(_04200_),
    .B(_04201_),
    .S(_03915_),
    .Z(_04202_));
 MUX2_X1 _10471_ (.A(\registers[24][4] ),
    .B(\registers[26][4] ),
    .S(_03234_),
    .Z(_04203_));
 MUX2_X1 _10472_ (.A(\registers[25][4] ),
    .B(\registers[27][4] ),
    .S(_03880_),
    .Z(_04204_));
 MUX2_X1 _10473_ (.A(_04203_),
    .B(_04204_),
    .S(_03954_),
    .Z(_04205_));
 MUX2_X1 _10474_ (.A(_04202_),
    .B(_04205_),
    .S(_03385_),
    .Z(_04206_));
 AOI221_X2 _10475_ (.A(_03130_),
    .B1(_04196_),
    .B2(_04199_),
    .C1(_04206_),
    .C2(_03994_),
    .ZN(_04207_));
 MUX2_X1 _10476_ (.A(\registers[0][4] ),
    .B(\registers[1][4] ),
    .S(_03319_),
    .Z(_04208_));
 NOR2_X1 _10477_ (.A1(_03137_),
    .A2(_04208_),
    .ZN(_04209_));
 MUX2_X1 _10478_ (.A(\registers[2][4] ),
    .B(\registers[3][4] ),
    .S(_03386_),
    .Z(_04210_));
 NOR3_X1 _10479_ (.A1(_03153_),
    .A2(_03134_),
    .A3(_04210_),
    .ZN(_04211_));
 MUX2_X1 _10480_ (.A(\registers[4][4] ),
    .B(\registers[5][4] ),
    .S(_03227_),
    .Z(_04212_));
 NOR3_X1 _10481_ (.A1(_03159_),
    .A2(_03258_),
    .A3(_04212_),
    .ZN(_04213_));
 MUX2_X1 _10482_ (.A(\registers[6][4] ),
    .B(\registers[7][4] ),
    .S(_03223_),
    .Z(_04214_));
 NOR2_X1 _10483_ (.A1(_03144_),
    .A2(_04214_),
    .ZN(_04215_));
 NOR4_X1 _10484_ (.A1(_04209_),
    .A2(_04211_),
    .A3(_04213_),
    .A4(_04215_),
    .ZN(_04216_));
 MUX2_X1 _10485_ (.A(\registers[12][4] ),
    .B(\registers[14][4] ),
    .S(_03255_),
    .Z(_04217_));
 MUX2_X1 _10486_ (.A(\registers[13][4] ),
    .B(\registers[15][4] ),
    .S(_03392_),
    .Z(_04218_));
 MUX2_X1 _10487_ (.A(_04217_),
    .B(_04218_),
    .S(_03306_),
    .Z(_04219_));
 MUX2_X1 _10488_ (.A(\registers[8][4] ),
    .B(\registers[10][4] ),
    .S(_03394_),
    .Z(_04220_));
 MUX2_X1 _10489_ (.A(\registers[9][4] ),
    .B(\registers[11][4] ),
    .S(_03400_),
    .Z(_04221_));
 MUX2_X1 _10490_ (.A(_04220_),
    .B(_04221_),
    .S(_03396_),
    .Z(_04222_));
 MUX2_X2 _10491_ (.A(_04219_),
    .B(_04222_),
    .S(_03259_),
    .Z(_04223_));
 OAI221_X2 _10492_ (.A(_03996_),
    .B1(_03182_),
    .B2(_04216_),
    .C1(_04223_),
    .C2(_03210_),
    .ZN(_04224_));
 OAI22_X1 _10493_ (.A1(_04190_),
    .A2(_04015_),
    .B1(_04207_),
    .B2(_04224_),
    .ZN(_00387_));
 INV_X1 _10494_ (.A(net64),
    .ZN(_04225_));
 MUX2_X1 _10495_ (.A(\registers[0][5] ),
    .B(\registers[1][5] ),
    .S(_03145_),
    .Z(_04226_));
 MUX2_X1 _10496_ (.A(\registers[6][5] ),
    .B(\registers[7][5] ),
    .S(_03169_),
    .Z(_04227_));
 OAI22_X1 _10497_ (.A1(_03136_),
    .A2(_04226_),
    .B1(_04227_),
    .B2(_03143_),
    .ZN(_04228_));
 MUX2_X1 _10498_ (.A(\registers[2][5] ),
    .B(\registers[3][5] ),
    .S(_03194_),
    .Z(_04229_));
 INV_X1 _10499_ (.A(_04229_),
    .ZN(_04230_));
 AOI21_X1 _10500_ (.A(_04228_),
    .B1(_04230_),
    .B2(_03981_),
    .ZN(_04231_));
 MUX2_X1 _10501_ (.A(\registers[4][5] ),
    .B(\registers[5][5] ),
    .S(_03909_),
    .Z(_04232_));
 INV_X1 _10502_ (.A(_04232_),
    .ZN(_04233_));
 AOI21_X1 _10503_ (.A(_03261_),
    .B1(_03983_),
    .B2(_04233_),
    .ZN(_04234_));
 MUX2_X1 _10504_ (.A(\registers[12][5] ),
    .B(\registers[14][5] ),
    .S(_03142_),
    .Z(_04235_));
 MUX2_X1 _10505_ (.A(\registers[13][5] ),
    .B(\registers[15][5] ),
    .S(_03232_),
    .Z(_04236_));
 MUX2_X1 _10506_ (.A(_04235_),
    .B(_04236_),
    .S(_03915_),
    .Z(_04237_));
 MUX2_X1 _10507_ (.A(\registers[8][5] ),
    .B(\registers[10][5] ),
    .S(_03234_),
    .Z(_04238_));
 MUX2_X1 _10508_ (.A(\registers[9][5] ),
    .B(\registers[11][5] ),
    .S(_03238_),
    .Z(_04239_));
 MUX2_X1 _10509_ (.A(_04238_),
    .B(_04239_),
    .S(_03954_),
    .Z(_04240_));
 MUX2_X2 _10510_ (.A(_04237_),
    .B(_04240_),
    .S(_03385_),
    .Z(_04241_));
 AOI221_X2 _10511_ (.A(_03714_),
    .B1(_04231_),
    .B2(_04234_),
    .C1(_04241_),
    .C2(_03994_),
    .ZN(_04242_));
 MUX2_X1 _10512_ (.A(\registers[28][5] ),
    .B(\registers[30][5] ),
    .S(_03152_),
    .Z(_04243_));
 MUX2_X1 _10513_ (.A(\registers[29][5] ),
    .B(\registers[31][5] ),
    .S(_03247_),
    .Z(_04244_));
 MUX2_X1 _10514_ (.A(_04243_),
    .B(_04244_),
    .S(_03380_),
    .Z(_04245_));
 MUX2_X1 _10515_ (.A(\registers[24][5] ),
    .B(\registers[26][5] ),
    .S(_03249_),
    .Z(_04246_));
 MUX2_X1 _10516_ (.A(\registers[25][5] ),
    .B(\registers[27][5] ),
    .S(_03253_),
    .Z(_04247_));
 MUX2_X1 _10517_ (.A(_04246_),
    .B(_04247_),
    .S(_03251_),
    .Z(_04248_));
 MUX2_X1 _10518_ (.A(_04245_),
    .B(_04248_),
    .S(_03629_),
    .Z(_04249_));
 MUX2_X1 _10519_ (.A(\registers[16][5] ),
    .B(\registers[17][5] ),
    .S(_03590_),
    .Z(_04250_));
 NOR2_X1 _10520_ (.A1(_03264_),
    .A2(_04250_),
    .ZN(_04251_));
 MUX2_X1 _10521_ (.A(\registers[18][5] ),
    .B(\registers[19][5] ),
    .S(_03170_),
    .Z(_04252_));
 NOR3_X1 _10522_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_04252_),
    .ZN(_04253_));
 MUX2_X1 _10523_ (.A(\registers[20][5] ),
    .B(\registers[21][5] ),
    .S(_03149_),
    .Z(_04254_));
 NOR3_X1 _10524_ (.A1(_03271_),
    .A2(_03706_),
    .A3(_04254_),
    .ZN(_04255_));
 MUX2_X1 _10525_ (.A(\registers[22][5] ),
    .B(\registers[23][5] ),
    .S(_03311_),
    .Z(_04256_));
 NOR2_X1 _10526_ (.A1(_03275_),
    .A2(_04256_),
    .ZN(_04257_));
 NOR4_X1 _10527_ (.A1(_04251_),
    .A2(_04253_),
    .A3(_04255_),
    .A4(_04257_),
    .ZN(_04258_));
 OAI221_X1 _10528_ (.A(_03996_),
    .B1(_03733_),
    .B2(_04249_),
    .C1(_04258_),
    .C2(_03750_),
    .ZN(_04259_));
 OAI22_X1 _10529_ (.A1(_04225_),
    .A2(_04015_),
    .B1(_04242_),
    .B2(_04259_),
    .ZN(_00388_));
 INV_X1 _10530_ (.A(net65),
    .ZN(_04260_));
 MUX2_X1 _10531_ (.A(\registers[16][6] ),
    .B(\registers[17][6] ),
    .S(_03145_),
    .Z(_04261_));
 MUX2_X1 _10532_ (.A(\registers[22][6] ),
    .B(\registers[23][6] ),
    .S(_03169_),
    .Z(_04262_));
 OAI22_X1 _10533_ (.A1(_03136_),
    .A2(_04261_),
    .B1(_04262_),
    .B2(_03143_),
    .ZN(_04263_));
 MUX2_X1 _10534_ (.A(\registers[18][6] ),
    .B(\registers[19][6] ),
    .S(_03194_),
    .Z(_04264_));
 INV_X1 _10535_ (.A(_04264_),
    .ZN(_04265_));
 AOI21_X1 _10536_ (.A(_04263_),
    .B1(_04265_),
    .B2(_03981_),
    .ZN(_04266_));
 MUX2_X1 _10537_ (.A(\registers[20][6] ),
    .B(\registers[21][6] ),
    .S(_03140_),
    .Z(_04267_));
 INV_X1 _10538_ (.A(_04267_),
    .ZN(_04268_));
 AOI21_X1 _10539_ (.A(_03261_),
    .B1(_03983_),
    .B2(_04268_),
    .ZN(_04269_));
 MUX2_X1 _10540_ (.A(\registers[28][6] ),
    .B(\registers[30][6] ),
    .S(_03142_),
    .Z(_04270_));
 MUX2_X1 _10541_ (.A(\registers[29][6] ),
    .B(\registers[31][6] ),
    .S(_03232_),
    .Z(_04271_));
 MUX2_X1 _10542_ (.A(_04270_),
    .B(_04271_),
    .S(_03272_),
    .Z(_04272_));
 MUX2_X1 _10543_ (.A(\registers[24][6] ),
    .B(\registers[26][6] ),
    .S(_03234_),
    .Z(_04273_));
 MUX2_X1 _10544_ (.A(\registers[25][6] ),
    .B(\registers[27][6] ),
    .S(_03238_),
    .Z(_04274_));
 MUX2_X1 _10545_ (.A(_04273_),
    .B(_04274_),
    .S(_03954_),
    .Z(_04275_));
 MUX2_X1 _10546_ (.A(_04272_),
    .B(_04275_),
    .S(_03385_),
    .Z(_04276_));
 AOI221_X1 _10547_ (.A(_03130_),
    .B1(_04266_),
    .B2(_04269_),
    .C1(_04276_),
    .C2(_03994_),
    .ZN(_04277_));
 MUX2_X1 _10548_ (.A(\registers[0][6] ),
    .B(\registers[1][6] ),
    .S(_03319_),
    .Z(_04278_));
 NOR2_X1 _10549_ (.A1(_03137_),
    .A2(_04278_),
    .ZN(_04279_));
 MUX2_X1 _10550_ (.A(\registers[2][6] ),
    .B(\registers[3][6] ),
    .S(_03386_),
    .Z(_04280_));
 NOR3_X1 _10551_ (.A1(_03153_),
    .A2(_03134_),
    .A3(_04280_),
    .ZN(_04281_));
 MUX2_X1 _10552_ (.A(\registers[4][6] ),
    .B(\registers[5][6] ),
    .S(_03227_),
    .Z(_04282_));
 NOR3_X1 _10553_ (.A1(_03159_),
    .A2(_03258_),
    .A3(_04282_),
    .ZN(_04283_));
 MUX2_X1 _10554_ (.A(\registers[6][6] ),
    .B(\registers[7][6] ),
    .S(_03223_),
    .Z(_04284_));
 NOR2_X1 _10555_ (.A1(_03144_),
    .A2(_04284_),
    .ZN(_04285_));
 NOR4_X1 _10556_ (.A1(_04279_),
    .A2(_04281_),
    .A3(_04283_),
    .A4(_04285_),
    .ZN(_04286_));
 MUX2_X1 _10557_ (.A(\registers[12][6] ),
    .B(\registers[14][6] ),
    .S(_03255_),
    .Z(_04287_));
 MUX2_X1 _10558_ (.A(\registers[13][6] ),
    .B(\registers[15][6] ),
    .S(_03392_),
    .Z(_04288_));
 MUX2_X1 _10559_ (.A(_04287_),
    .B(_04288_),
    .S(_03306_),
    .Z(_04289_));
 MUX2_X1 _10560_ (.A(\registers[8][6] ),
    .B(\registers[10][6] ),
    .S(_03394_),
    .Z(_04290_));
 MUX2_X1 _10561_ (.A(\registers[9][6] ),
    .B(\registers[11][6] ),
    .S(_03398_),
    .Z(_04291_));
 MUX2_X1 _10562_ (.A(_04290_),
    .B(_04291_),
    .S(_03396_),
    .Z(_04292_));
 MUX2_X2 _10563_ (.A(_04289_),
    .B(_04292_),
    .S(_03259_),
    .Z(_04293_));
 OAI221_X2 _10564_ (.A(_03996_),
    .B1(_03182_),
    .B2(_04286_),
    .C1(_04293_),
    .C2(_03210_),
    .ZN(_04294_));
 OAI22_X1 _10565_ (.A1(_04260_),
    .A2(_04015_),
    .B1(_04277_),
    .B2(_04294_),
    .ZN(_00389_));
 INV_X1 _10566_ (.A(net66),
    .ZN(_04295_));
 MUX2_X1 _10567_ (.A(\registers[0][7] ),
    .B(\registers[1][7] ),
    .S(_03145_),
    .Z(_04296_));
 MUX2_X1 _10568_ (.A(\registers[6][7] ),
    .B(\registers[7][7] ),
    .S(_03169_),
    .Z(_04297_));
 OAI22_X1 _10569_ (.A1(_03136_),
    .A2(_04296_),
    .B1(_04297_),
    .B2(_03143_),
    .ZN(_04298_));
 MUX2_X1 _10570_ (.A(\registers[2][7] ),
    .B(\registers[3][7] ),
    .S(_03194_),
    .Z(_04299_));
 INV_X1 _10571_ (.A(_04299_),
    .ZN(_04300_));
 AOI21_X1 _10572_ (.A(_04298_),
    .B1(_04300_),
    .B2(_03981_),
    .ZN(_04301_));
 MUX2_X1 _10573_ (.A(\registers[4][7] ),
    .B(\registers[5][7] ),
    .S(_03140_),
    .Z(_04302_));
 INV_X1 _10574_ (.A(_04302_),
    .ZN(_04303_));
 AOI21_X1 _10575_ (.A(_03261_),
    .B1(_03983_),
    .B2(_04303_),
    .ZN(_04304_));
 MUX2_X1 _10576_ (.A(\registers[12][7] ),
    .B(\registers[14][7] ),
    .S(_03142_),
    .Z(_04305_));
 MUX2_X1 _10577_ (.A(\registers[13][7] ),
    .B(\registers[15][7] ),
    .S(_03232_),
    .Z(_04306_));
 MUX2_X1 _10578_ (.A(_04305_),
    .B(_04306_),
    .S(_03272_),
    .Z(_04307_));
 MUX2_X1 _10579_ (.A(\registers[8][7] ),
    .B(\registers[10][7] ),
    .S(_03234_),
    .Z(_04308_));
 MUX2_X1 _10580_ (.A(\registers[9][7] ),
    .B(\registers[11][7] ),
    .S(_03238_),
    .Z(_04309_));
 MUX2_X1 _10581_ (.A(_04308_),
    .B(_04309_),
    .S(_03236_),
    .Z(_04310_));
 MUX2_X2 _10582_ (.A(_04307_),
    .B(_04310_),
    .S(_03385_),
    .Z(_04311_));
 AOI221_X2 _10583_ (.A(_03714_),
    .B1(_04301_),
    .B2(_04304_),
    .C1(_04311_),
    .C2(_03994_),
    .ZN(_04312_));
 MUX2_X1 _10584_ (.A(\registers[28][7] ),
    .B(\registers[30][7] ),
    .S(_03152_),
    .Z(_04313_));
 MUX2_X1 _10585_ (.A(\registers[29][7] ),
    .B(\registers[31][7] ),
    .S(_03247_),
    .Z(_04314_));
 MUX2_X1 _10586_ (.A(_04313_),
    .B(_04314_),
    .S(_03380_),
    .Z(_04315_));
 MUX2_X1 _10587_ (.A(\registers[24][7] ),
    .B(\registers[26][7] ),
    .S(_03249_),
    .Z(_04316_));
 MUX2_X1 _10588_ (.A(\registers[25][7] ),
    .B(\registers[27][7] ),
    .S(_03253_),
    .Z(_04317_));
 MUX2_X1 _10589_ (.A(_04316_),
    .B(_04317_),
    .S(_03251_),
    .Z(_04318_));
 MUX2_X1 _10590_ (.A(_04315_),
    .B(_04318_),
    .S(_03629_),
    .Z(_04319_));
 MUX2_X1 _10591_ (.A(\registers[16][7] ),
    .B(\registers[17][7] ),
    .S(_03185_),
    .Z(_04320_));
 NOR2_X1 _10592_ (.A1(_03264_),
    .A2(_04320_),
    .ZN(_04321_));
 MUX2_X1 _10593_ (.A(\registers[18][7] ),
    .B(\registers[19][7] ),
    .S(_03170_),
    .Z(_04322_));
 NOR3_X1 _10594_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_04322_),
    .ZN(_04323_));
 MUX2_X1 _10595_ (.A(\registers[20][7] ),
    .B(\registers[21][7] ),
    .S(_03149_),
    .Z(_04324_));
 NOR3_X1 _10596_ (.A1(_03271_),
    .A2(_03706_),
    .A3(_04324_),
    .ZN(_04325_));
 MUX2_X1 _10597_ (.A(\registers[22][7] ),
    .B(\registers[23][7] ),
    .S(_03311_),
    .Z(_04326_));
 NOR2_X1 _10598_ (.A1(_03275_),
    .A2(_04326_),
    .ZN(_04327_));
 NOR4_X2 _10599_ (.A1(_04321_),
    .A2(_04323_),
    .A3(_04325_),
    .A4(_04327_),
    .ZN(_04328_));
 OAI221_X1 _10600_ (.A(_03996_),
    .B1(_03733_),
    .B2(_04319_),
    .C1(_04328_),
    .C2(_03750_),
    .ZN(_04329_));
 OAI22_X1 _10601_ (.A1(_04295_),
    .A2(_04015_),
    .B1(_04312_),
    .B2(_04329_),
    .ZN(_00390_));
 INV_X1 _10602_ (.A(net67),
    .ZN(_04330_));
 MUX2_X1 _10603_ (.A(\registers[0][8] ),
    .B(\registers[1][8] ),
    .S(_03145_),
    .Z(_04331_));
 MUX2_X1 _10604_ (.A(\registers[6][8] ),
    .B(\registers[7][8] ),
    .S(_03169_),
    .Z(_04332_));
 OAI22_X1 _10605_ (.A1(_03136_),
    .A2(_04331_),
    .B1(_04332_),
    .B2(_03143_),
    .ZN(_04333_));
 MUX2_X1 _10606_ (.A(\registers[2][8] ),
    .B(\registers[3][8] ),
    .S(_03194_),
    .Z(_04334_));
 INV_X1 _10607_ (.A(_04334_),
    .ZN(_04335_));
 AOI21_X1 _10608_ (.A(_04333_),
    .B1(_04335_),
    .B2(_03154_),
    .ZN(_04336_));
 MUX2_X1 _10609_ (.A(\registers[4][8] ),
    .B(\registers[5][8] ),
    .S(_03140_),
    .Z(_04337_));
 INV_X1 _10610_ (.A(_04337_),
    .ZN(_04338_));
 AOI21_X1 _10611_ (.A(_03261_),
    .B1(_03161_),
    .B2(_04338_),
    .ZN(_04339_));
 MUX2_X1 _10612_ (.A(\registers[12][8] ),
    .B(\registers[14][8] ),
    .S(_03142_),
    .Z(_04340_));
 MUX2_X1 _10613_ (.A(\registers[13][8] ),
    .B(\registers[15][8] ),
    .S(_03232_),
    .Z(_04341_));
 MUX2_X1 _10614_ (.A(_04340_),
    .B(_04341_),
    .S(_03272_),
    .Z(_04342_));
 MUX2_X1 _10615_ (.A(\registers[8][8] ),
    .B(\registers[10][8] ),
    .S(_03234_),
    .Z(_04343_));
 MUX2_X1 _10616_ (.A(\registers[9][8] ),
    .B(\registers[11][8] ),
    .S(_03238_),
    .Z(_04344_));
 MUX2_X1 _10617_ (.A(_04343_),
    .B(_04344_),
    .S(_03236_),
    .Z(_04345_));
 MUX2_X2 _10618_ (.A(_04342_),
    .B(_04345_),
    .S(_03385_),
    .Z(_04346_));
 AOI221_X2 _10619_ (.A(_03714_),
    .B1(_04336_),
    .B2(_04339_),
    .C1(_04346_),
    .C2(_03158_),
    .ZN(_04347_));
 MUX2_X1 _10620_ (.A(\registers[28][8] ),
    .B(\registers[30][8] ),
    .S(_03152_),
    .Z(_04348_));
 MUX2_X1 _10621_ (.A(\registers[29][8] ),
    .B(\registers[31][8] ),
    .S(_03247_),
    .Z(_04349_));
 MUX2_X1 _10622_ (.A(_04348_),
    .B(_04349_),
    .S(_03380_),
    .Z(_04350_));
 MUX2_X1 _10623_ (.A(\registers[24][8] ),
    .B(\registers[26][8] ),
    .S(_03249_),
    .Z(_04351_));
 MUX2_X1 _10624_ (.A(\registers[25][8] ),
    .B(\registers[27][8] ),
    .S(_03253_),
    .Z(_04352_));
 MUX2_X1 _10625_ (.A(_04351_),
    .B(_04352_),
    .S(_03251_),
    .Z(_04353_));
 MUX2_X1 _10626_ (.A(_04350_),
    .B(_04353_),
    .S(_03315_),
    .Z(_04354_));
 MUX2_X1 _10627_ (.A(\registers[16][8] ),
    .B(\registers[17][8] ),
    .S(_03185_),
    .Z(_04355_));
 NOR2_X1 _10628_ (.A1(_03264_),
    .A2(_04355_),
    .ZN(_04356_));
 MUX2_X1 _10629_ (.A(\registers[18][8] ),
    .B(\registers[19][8] ),
    .S(_03170_),
    .Z(_04357_));
 NOR3_X1 _10630_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_04357_),
    .ZN(_04358_));
 MUX2_X1 _10631_ (.A(\registers[20][8] ),
    .B(\registers[21][8] ),
    .S(_03149_),
    .Z(_04359_));
 NOR3_X1 _10632_ (.A1(_03271_),
    .A2(_03706_),
    .A3(_04359_),
    .ZN(_04360_));
 MUX2_X1 _10633_ (.A(\registers[22][8] ),
    .B(\registers[23][8] ),
    .S(_03311_),
    .Z(_04361_));
 NOR2_X1 _10634_ (.A1(_03275_),
    .A2(_04361_),
    .ZN(_04362_));
 NOR4_X2 _10635_ (.A1(_04356_),
    .A2(_04358_),
    .A3(_04360_),
    .A4(_04362_),
    .ZN(_04363_));
 OAI221_X1 _10636_ (.A(_03180_),
    .B1(_03733_),
    .B2(_04354_),
    .C1(_04363_),
    .C2(_03750_),
    .ZN(_04364_));
 OAI22_X1 _10637_ (.A1(_04330_),
    .A2(_04015_),
    .B1(_04347_),
    .B2(_04364_),
    .ZN(_00391_));
 INV_X1 _10638_ (.A(net68),
    .ZN(_04365_));
 MUX2_X1 _10639_ (.A(\registers[0][9] ),
    .B(\registers[1][9] ),
    .S(_03145_),
    .Z(_04366_));
 MUX2_X1 _10640_ (.A(\registers[6][9] ),
    .B(\registers[7][9] ),
    .S(_03169_),
    .Z(_04367_));
 OAI22_X1 _10641_ (.A1(_03136_),
    .A2(_04366_),
    .B1(_04367_),
    .B2(_03143_),
    .ZN(_04368_));
 MUX2_X1 _10642_ (.A(\registers[2][9] ),
    .B(\registers[3][9] ),
    .S(_03194_),
    .Z(_04369_));
 INV_X1 _10643_ (.A(_04369_),
    .ZN(_04370_));
 AOI21_X1 _10644_ (.A(_04368_),
    .B1(_04370_),
    .B2(_03154_),
    .ZN(_04371_));
 MUX2_X1 _10645_ (.A(\registers[4][9] ),
    .B(\registers[5][9] ),
    .S(_03140_),
    .Z(_04372_));
 INV_X1 _10646_ (.A(_04372_),
    .ZN(_04373_));
 AOI21_X1 _10647_ (.A(_03261_),
    .B1(_03161_),
    .B2(_04373_),
    .ZN(_04374_));
 MUX2_X1 _10648_ (.A(\registers[12][9] ),
    .B(\registers[14][9] ),
    .S(_03142_),
    .Z(_04375_));
 MUX2_X1 _10649_ (.A(\registers[13][9] ),
    .B(\registers[15][9] ),
    .S(_03232_),
    .Z(_04376_));
 MUX2_X1 _10650_ (.A(_04375_),
    .B(_04376_),
    .S(_03272_),
    .Z(_04377_));
 MUX2_X1 _10651_ (.A(\registers[8][9] ),
    .B(\registers[10][9] ),
    .S(_03234_),
    .Z(_04378_));
 MUX2_X1 _10652_ (.A(\registers[9][9] ),
    .B(\registers[11][9] ),
    .S(_03238_),
    .Z(_04379_));
 MUX2_X1 _10653_ (.A(_04378_),
    .B(_04379_),
    .S(_03236_),
    .Z(_04380_));
 MUX2_X2 _10654_ (.A(_04377_),
    .B(_04380_),
    .S(_03385_),
    .Z(_04381_));
 AOI221_X2 _10655_ (.A(_03714_),
    .B1(_04371_),
    .B2(_04374_),
    .C1(_04381_),
    .C2(_03158_),
    .ZN(_04382_));
 MUX2_X1 _10656_ (.A(\registers[28][9] ),
    .B(\registers[30][9] ),
    .S(_03152_),
    .Z(_04383_));
 MUX2_X1 _10657_ (.A(\registers[29][9] ),
    .B(\registers[31][9] ),
    .S(_03247_),
    .Z(_04384_));
 MUX2_X1 _10658_ (.A(_04383_),
    .B(_04384_),
    .S(_03380_),
    .Z(_04385_));
 MUX2_X1 _10659_ (.A(\registers[24][9] ),
    .B(\registers[26][9] ),
    .S(_03249_),
    .Z(_04386_));
 MUX2_X1 _10660_ (.A(\registers[25][9] ),
    .B(\registers[27][9] ),
    .S(_03253_),
    .Z(_04387_));
 MUX2_X1 _10661_ (.A(_04386_),
    .B(_04387_),
    .S(_03251_),
    .Z(_04388_));
 MUX2_X1 _10662_ (.A(_04385_),
    .B(_04388_),
    .S(_03315_),
    .Z(_04389_));
 MUX2_X1 _10663_ (.A(\registers[16][9] ),
    .B(\registers[17][9] ),
    .S(_03185_),
    .Z(_04390_));
 NOR2_X1 _10664_ (.A1(_03264_),
    .A2(_04390_),
    .ZN(_04391_));
 MUX2_X1 _10665_ (.A(\registers[18][9] ),
    .B(\registers[19][9] ),
    .S(_03170_),
    .Z(_04392_));
 NOR3_X1 _10666_ (.A1(_03267_),
    .A2(_03268_),
    .A3(_04392_),
    .ZN(_04393_));
 MUX2_X1 _10667_ (.A(\registers[20][9] ),
    .B(\registers[21][9] ),
    .S(_03149_),
    .Z(_04394_));
 NOR3_X1 _10668_ (.A1(_03271_),
    .A2(_03175_),
    .A3(_04394_),
    .ZN(_04395_));
 MUX2_X1 _10669_ (.A(\registers[22][9] ),
    .B(\registers[23][9] ),
    .S(_03311_),
    .Z(_04396_));
 NOR2_X1 _10670_ (.A1(_03275_),
    .A2(_04396_),
    .ZN(_04397_));
 NOR4_X1 _10671_ (.A1(_04391_),
    .A2(_04393_),
    .A3(_04395_),
    .A4(_04397_),
    .ZN(_04398_));
 OAI221_X1 _10672_ (.A(_03180_),
    .B1(_03733_),
    .B2(_04389_),
    .C1(_04398_),
    .C2(_03750_),
    .ZN(_04399_));
 OAI22_X1 _10673_ (.A1(_04365_),
    .A2(_03214_),
    .B1(_04382_),
    .B2(_04399_),
    .ZN(_00392_));
 NOR2_X1 _10674_ (.A1(_01138_),
    .A2(_01737_),
    .ZN(_04400_));
 CLKBUF_X3 _10675_ (.A(_04400_),
    .Z(_04401_));
 CLKBUF_X3 _10676_ (.A(_04401_),
    .Z(_04402_));
 NAND2_X1 _10677_ (.A1(_01137_),
    .A2(_04402_),
    .ZN(_04403_));
 CLKBUF_X3 _10678_ (.A(_01674_),
    .Z(_04404_));
 NAND2_X1 _10679_ (.A1(_04404_),
    .A2(\registers[0][0] ),
    .ZN(_04405_));
 CLKBUF_X3 _10680_ (.A(_04401_),
    .Z(_04406_));
 OAI21_X1 _10681_ (.A(_04403_),
    .B1(_04405_),
    .B2(_04406_),
    .ZN(_00393_));
 NAND2_X1 _10682_ (.A1(_01149_),
    .A2(_04402_),
    .ZN(_04407_));
 NAND2_X1 _10683_ (.A1(_04404_),
    .A2(\registers[0][10] ),
    .ZN(_04408_));
 OAI21_X1 _10684_ (.A(_04407_),
    .B1(_04408_),
    .B2(_04406_),
    .ZN(_00394_));
 NAND2_X1 _10685_ (.A1(_01153_),
    .A2(_04402_),
    .ZN(_04409_));
 NAND2_X1 _10686_ (.A1(_04404_),
    .A2(\registers[0][11] ),
    .ZN(_04410_));
 OAI21_X1 _10687_ (.A(_04409_),
    .B1(_04410_),
    .B2(_04406_),
    .ZN(_00395_));
 NAND2_X1 _10688_ (.A1(_01158_),
    .A2(_04402_),
    .ZN(_04411_));
 NAND2_X1 _10689_ (.A1(_04404_),
    .A2(\registers[0][12] ),
    .ZN(_04412_));
 OAI21_X1 _10690_ (.A(_04411_),
    .B1(_04412_),
    .B2(_04406_),
    .ZN(_00396_));
 NAND2_X1 _10691_ (.A1(_01162_),
    .A2(_04402_),
    .ZN(_04413_));
 NAND2_X1 _10692_ (.A1(_04404_),
    .A2(\registers[0][13] ),
    .ZN(_04414_));
 OAI21_X1 _10693_ (.A(_04413_),
    .B1(_04414_),
    .B2(_04406_),
    .ZN(_00397_));
 NAND2_X1 _10694_ (.A1(_01166_),
    .A2(_04402_),
    .ZN(_04415_));
 NAND2_X1 _10695_ (.A1(_04404_),
    .A2(\registers[0][14] ),
    .ZN(_04416_));
 OAI21_X1 _10696_ (.A(_04415_),
    .B1(_04416_),
    .B2(_04406_),
    .ZN(_00398_));
 NAND2_X1 _10697_ (.A1(_01170_),
    .A2(_04402_),
    .ZN(_04417_));
 NAND2_X1 _10698_ (.A1(_04404_),
    .A2(\registers[0][15] ),
    .ZN(_04418_));
 OAI21_X1 _10699_ (.A(_04417_),
    .B1(_04418_),
    .B2(_04406_),
    .ZN(_00399_));
 NAND2_X1 _10700_ (.A1(_01174_),
    .A2(_04402_),
    .ZN(_04419_));
 NAND2_X1 _10701_ (.A1(_04404_),
    .A2(\registers[0][16] ),
    .ZN(_04420_));
 OAI21_X1 _10702_ (.A(_04419_),
    .B1(_04420_),
    .B2(_04406_),
    .ZN(_00400_));
 CLKBUF_X3 _10703_ (.A(_04401_),
    .Z(_04421_));
 NAND2_X1 _10704_ (.A1(_01178_),
    .A2(_04421_),
    .ZN(_04422_));
 NAND2_X1 _10705_ (.A1(_04404_),
    .A2(\registers[0][17] ),
    .ZN(_04423_));
 OAI21_X1 _10706_ (.A(_04422_),
    .B1(_04423_),
    .B2(_04406_),
    .ZN(_00401_));
 NAND2_X1 _10707_ (.A1(_01183_),
    .A2(_04421_),
    .ZN(_04424_));
 NAND2_X1 _10708_ (.A1(_04404_),
    .A2(\registers[0][18] ),
    .ZN(_04425_));
 OAI21_X1 _10709_ (.A(_04424_),
    .B1(_04425_),
    .B2(_04406_),
    .ZN(_00402_));
 NAND2_X1 _10710_ (.A1(_01187_),
    .A2(_04421_),
    .ZN(_04426_));
 CLKBUF_X3 _10711_ (.A(_01674_),
    .Z(_04427_));
 NAND2_X1 _10712_ (.A1(_04427_),
    .A2(\registers[0][19] ),
    .ZN(_04428_));
 CLKBUF_X3 _10713_ (.A(_04401_),
    .Z(_04429_));
 OAI21_X1 _10714_ (.A(_04426_),
    .B1(_04428_),
    .B2(_04429_),
    .ZN(_00403_));
 NAND2_X1 _10715_ (.A1(_01192_),
    .A2(_04421_),
    .ZN(_04430_));
 NAND2_X1 _10716_ (.A1(_04427_),
    .A2(\registers[0][1] ),
    .ZN(_04431_));
 OAI21_X1 _10717_ (.A(_04430_),
    .B1(_04431_),
    .B2(_04429_),
    .ZN(_00404_));
 NAND2_X1 _10718_ (.A1(_01196_),
    .A2(_04421_),
    .ZN(_04432_));
 NAND2_X1 _10719_ (.A1(_04427_),
    .A2(\registers[0][20] ),
    .ZN(_04433_));
 OAI21_X1 _10720_ (.A(_04432_),
    .B1(_04433_),
    .B2(_04429_),
    .ZN(_00405_));
 NAND2_X1 _10721_ (.A1(_01201_),
    .A2(_04421_),
    .ZN(_04434_));
 NAND2_X1 _10722_ (.A1(_04427_),
    .A2(\registers[0][21] ),
    .ZN(_04435_));
 OAI21_X1 _10723_ (.A(_04434_),
    .B1(_04435_),
    .B2(_04429_),
    .ZN(_00406_));
 NAND2_X1 _10724_ (.A1(_01205_),
    .A2(_04421_),
    .ZN(_04436_));
 NAND2_X1 _10725_ (.A1(_04427_),
    .A2(\registers[0][22] ),
    .ZN(_04437_));
 OAI21_X1 _10726_ (.A(_04436_),
    .B1(_04437_),
    .B2(_04429_),
    .ZN(_00407_));
 NAND2_X1 _10727_ (.A1(_01209_),
    .A2(_04421_),
    .ZN(_04438_));
 NAND2_X1 _10728_ (.A1(_04427_),
    .A2(\registers[0][23] ),
    .ZN(_04439_));
 OAI21_X1 _10729_ (.A(_04438_),
    .B1(_04439_),
    .B2(_04429_),
    .ZN(_00408_));
 NAND2_X1 _10730_ (.A1(_01213_),
    .A2(_04421_),
    .ZN(_04440_));
 NAND2_X1 _10731_ (.A1(_04427_),
    .A2(\registers[0][24] ),
    .ZN(_04441_));
 OAI21_X1 _10732_ (.A(_04440_),
    .B1(_04441_),
    .B2(_04429_),
    .ZN(_00409_));
 NAND2_X1 _10733_ (.A1(_01217_),
    .A2(_04421_),
    .ZN(_04442_));
 NAND2_X1 _10734_ (.A1(_04427_),
    .A2(\registers[0][25] ),
    .ZN(_04443_));
 OAI21_X1 _10735_ (.A(_04442_),
    .B1(_04443_),
    .B2(_04429_),
    .ZN(_00410_));
 CLKBUF_X3 _10736_ (.A(_04401_),
    .Z(_04444_));
 NAND2_X1 _10737_ (.A1(_01221_),
    .A2(_04444_),
    .ZN(_04445_));
 NAND2_X1 _10738_ (.A1(_04427_),
    .A2(\registers[0][26] ),
    .ZN(_04446_));
 OAI21_X1 _10739_ (.A(_04445_),
    .B1(_04446_),
    .B2(_04429_),
    .ZN(_00411_));
 NAND2_X1 _10740_ (.A1(_01226_),
    .A2(_04444_),
    .ZN(_04447_));
 NAND2_X1 _10741_ (.A1(_04427_),
    .A2(\registers[0][27] ),
    .ZN(_04448_));
 OAI21_X1 _10742_ (.A(_04447_),
    .B1(_04448_),
    .B2(_04429_),
    .ZN(_00412_));
 NAND2_X1 _10743_ (.A1(_01230_),
    .A2(_04444_),
    .ZN(_04449_));
 CLKBUF_X3 _10744_ (.A(_01674_),
    .Z(_04450_));
 NAND2_X1 _10745_ (.A1(_04450_),
    .A2(\registers[0][28] ),
    .ZN(_04451_));
 CLKBUF_X3 _10746_ (.A(_04401_),
    .Z(_04452_));
 OAI21_X1 _10747_ (.A(_04449_),
    .B1(_04451_),
    .B2(_04452_),
    .ZN(_00413_));
 NAND2_X1 _10748_ (.A1(_01235_),
    .A2(_04444_),
    .ZN(_04453_));
 NAND2_X1 _10749_ (.A1(_04450_),
    .A2(\registers[0][29] ),
    .ZN(_04454_));
 OAI21_X1 _10750_ (.A(_04453_),
    .B1(_04454_),
    .B2(_04452_),
    .ZN(_00414_));
 NAND2_X1 _10751_ (.A1(_01239_),
    .A2(_04444_),
    .ZN(_04455_));
 NAND2_X1 _10752_ (.A1(_04450_),
    .A2(\registers[0][2] ),
    .ZN(_04456_));
 OAI21_X1 _10753_ (.A(_04455_),
    .B1(_04456_),
    .B2(_04452_),
    .ZN(_00415_));
 NAND2_X1 _10754_ (.A1(_01244_),
    .A2(_04444_),
    .ZN(_04457_));
 NAND2_X1 _10755_ (.A1(_04450_),
    .A2(\registers[0][30] ),
    .ZN(_04458_));
 OAI21_X1 _10756_ (.A(_04457_),
    .B1(_04458_),
    .B2(_04452_),
    .ZN(_00416_));
 NAND2_X1 _10757_ (.A1(_01089_),
    .A2(_04444_),
    .ZN(_04459_));
 NAND2_X1 _10758_ (.A1(_04450_),
    .A2(\registers[0][31] ),
    .ZN(_04460_));
 OAI21_X1 _10759_ (.A(_04459_),
    .B1(_04460_),
    .B2(_04452_),
    .ZN(_00417_));
 NAND2_X1 _10760_ (.A1(_01109_),
    .A2(_04444_),
    .ZN(_04461_));
 NAND2_X1 _10761_ (.A1(_04450_),
    .A2(\registers[0][3] ),
    .ZN(_04462_));
 OAI21_X1 _10762_ (.A(_04461_),
    .B1(_04462_),
    .B2(_04452_),
    .ZN(_00418_));
 NAND2_X1 _10763_ (.A1(_01113_),
    .A2(_04444_),
    .ZN(_04463_));
 NAND2_X1 _10764_ (.A1(_04450_),
    .A2(\registers[0][4] ),
    .ZN(_04464_));
 OAI21_X1 _10765_ (.A(_04463_),
    .B1(_04464_),
    .B2(_04452_),
    .ZN(_00419_));
 NAND2_X1 _10766_ (.A1(_01117_),
    .A2(_04444_),
    .ZN(_04465_));
 NAND2_X1 _10767_ (.A1(_04450_),
    .A2(\registers[0][5] ),
    .ZN(_04466_));
 OAI21_X1 _10768_ (.A(_04465_),
    .B1(_04466_),
    .B2(_04452_),
    .ZN(_00420_));
 NAND2_X1 _10769_ (.A1(_01121_),
    .A2(_04401_),
    .ZN(_04467_));
 NAND2_X1 _10770_ (.A1(_04450_),
    .A2(\registers[0][6] ),
    .ZN(_04468_));
 OAI21_X1 _10771_ (.A(_04467_),
    .B1(_04468_),
    .B2(_04452_),
    .ZN(_00421_));
 NAND2_X1 _10772_ (.A1(_01125_),
    .A2(_04401_),
    .ZN(_04469_));
 NAND2_X1 _10773_ (.A1(_04450_),
    .A2(\registers[0][7] ),
    .ZN(_04470_));
 OAI21_X1 _10774_ (.A(_04469_),
    .B1(_04470_),
    .B2(_04452_),
    .ZN(_00422_));
 NAND2_X1 _10775_ (.A1(_01129_),
    .A2(_04401_),
    .ZN(_04471_));
 BUF_X4 _10776_ (.A(_01674_),
    .Z(_04472_));
 NAND2_X1 _10777_ (.A1(_04472_),
    .A2(\registers[0][8] ),
    .ZN(_04473_));
 OAI21_X1 _10778_ (.A(_04471_),
    .B1(_04473_),
    .B2(_04402_),
    .ZN(_00423_));
 NAND2_X1 _10779_ (.A1(_01133_),
    .A2(_04401_),
    .ZN(_04474_));
 NAND2_X1 _10780_ (.A1(_04472_),
    .A2(\registers[0][9] ),
    .ZN(_04475_));
 OAI21_X1 _10781_ (.A(_04474_),
    .B1(_04475_),
    .B2(_04402_),
    .ZN(_00424_));
 NOR2_X1 _10782_ (.A1(_01141_),
    .A2(_01739_),
    .ZN(_04476_));
 BUF_X4 _10783_ (.A(_04476_),
    .Z(_04477_));
 BUF_X4 _10784_ (.A(_04477_),
    .Z(_04478_));
 NAND2_X1 _10785_ (.A1(_01137_),
    .A2(_04478_),
    .ZN(_04479_));
 NAND2_X1 _10786_ (.A1(_04472_),
    .A2(\registers[10][0] ),
    .ZN(_04480_));
 CLKBUF_X3 _10787_ (.A(_04477_),
    .Z(_04481_));
 OAI21_X1 _10788_ (.A(_04479_),
    .B1(_04480_),
    .B2(_04481_),
    .ZN(_00425_));
 NAND2_X1 _10789_ (.A1(_01149_),
    .A2(_04478_),
    .ZN(_04482_));
 NAND2_X1 _10790_ (.A1(_04472_),
    .A2(\registers[10][10] ),
    .ZN(_04483_));
 OAI21_X1 _10791_ (.A(_04482_),
    .B1(_04483_),
    .B2(_04481_),
    .ZN(_00426_));
 NAND2_X1 _10792_ (.A1(_01153_),
    .A2(_04478_),
    .ZN(_04484_));
 NAND2_X1 _10793_ (.A1(_04472_),
    .A2(\registers[10][11] ),
    .ZN(_04485_));
 OAI21_X1 _10794_ (.A(_04484_),
    .B1(_04485_),
    .B2(_04481_),
    .ZN(_00427_));
 NAND2_X1 _10795_ (.A1(_01158_),
    .A2(_04478_),
    .ZN(_04486_));
 NAND2_X1 _10796_ (.A1(_04472_),
    .A2(\registers[10][12] ),
    .ZN(_04487_));
 OAI21_X1 _10797_ (.A(_04486_),
    .B1(_04487_),
    .B2(_04481_),
    .ZN(_00428_));
 NAND2_X1 _10798_ (.A1(_01162_),
    .A2(_04478_),
    .ZN(_04488_));
 NAND2_X1 _10799_ (.A1(_04472_),
    .A2(\registers[10][13] ),
    .ZN(_04489_));
 OAI21_X1 _10800_ (.A(_04488_),
    .B1(_04489_),
    .B2(_04481_),
    .ZN(_00429_));
 NAND2_X1 _10801_ (.A1(_01166_),
    .A2(_04478_),
    .ZN(_04490_));
 NAND2_X1 _10802_ (.A1(_04472_),
    .A2(\registers[10][14] ),
    .ZN(_04491_));
 OAI21_X1 _10803_ (.A(_04490_),
    .B1(_04491_),
    .B2(_04481_),
    .ZN(_00430_));
 NAND2_X1 _10804_ (.A1(_01170_),
    .A2(_04478_),
    .ZN(_04492_));
 NAND2_X1 _10805_ (.A1(_04472_),
    .A2(\registers[10][15] ),
    .ZN(_04493_));
 OAI21_X1 _10806_ (.A(_04492_),
    .B1(_04493_),
    .B2(_04481_),
    .ZN(_00431_));
 NAND2_X1 _10807_ (.A1(_01174_),
    .A2(_04478_),
    .ZN(_04494_));
 NAND2_X1 _10808_ (.A1(_04472_),
    .A2(\registers[10][16] ),
    .ZN(_04495_));
 OAI21_X1 _10809_ (.A(_04494_),
    .B1(_04495_),
    .B2(_04481_),
    .ZN(_00432_));
 CLKBUF_X3 _10810_ (.A(_04477_),
    .Z(_04496_));
 NAND2_X1 _10811_ (.A1(_01178_),
    .A2(_04496_),
    .ZN(_04497_));
 BUF_X4 _10812_ (.A(_01103_),
    .Z(_04498_));
 CLKBUF_X3 _10813_ (.A(_04498_),
    .Z(_04499_));
 NAND2_X1 _10814_ (.A1(_04499_),
    .A2(\registers[10][17] ),
    .ZN(_04500_));
 OAI21_X1 _10815_ (.A(_04497_),
    .B1(_04500_),
    .B2(_04481_),
    .ZN(_00433_));
 NAND2_X1 _10816_ (.A1(_01183_),
    .A2(_04496_),
    .ZN(_04501_));
 NAND2_X1 _10817_ (.A1(_04499_),
    .A2(\registers[10][18] ),
    .ZN(_04502_));
 OAI21_X1 _10818_ (.A(_04501_),
    .B1(_04502_),
    .B2(_04481_),
    .ZN(_00434_));
 NAND2_X1 _10819_ (.A1(_01187_),
    .A2(_04496_),
    .ZN(_04503_));
 NAND2_X1 _10820_ (.A1(_04499_),
    .A2(\registers[10][19] ),
    .ZN(_04504_));
 CLKBUF_X3 _10821_ (.A(_04477_),
    .Z(_04505_));
 OAI21_X1 _10822_ (.A(_04503_),
    .B1(_04504_),
    .B2(_04505_),
    .ZN(_00435_));
 NAND2_X1 _10823_ (.A1(_01192_),
    .A2(_04496_),
    .ZN(_04506_));
 NAND2_X1 _10824_ (.A1(_04499_),
    .A2(\registers[10][1] ),
    .ZN(_04507_));
 OAI21_X1 _10825_ (.A(_04506_),
    .B1(_04507_),
    .B2(_04505_),
    .ZN(_00436_));
 NAND2_X1 _10826_ (.A1(_01196_),
    .A2(_04496_),
    .ZN(_04508_));
 NAND2_X1 _10827_ (.A1(_04499_),
    .A2(\registers[10][20] ),
    .ZN(_04509_));
 OAI21_X1 _10828_ (.A(_04508_),
    .B1(_04509_),
    .B2(_04505_),
    .ZN(_00437_));
 NAND2_X1 _10829_ (.A1(_01201_),
    .A2(_04496_),
    .ZN(_04510_));
 NAND2_X1 _10830_ (.A1(_04499_),
    .A2(\registers[10][21] ),
    .ZN(_04511_));
 OAI21_X1 _10831_ (.A(_04510_),
    .B1(_04511_),
    .B2(_04505_),
    .ZN(_00438_));
 NAND2_X1 _10832_ (.A1(_01205_),
    .A2(_04496_),
    .ZN(_04512_));
 NAND2_X1 _10833_ (.A1(_04499_),
    .A2(\registers[10][22] ),
    .ZN(_04513_));
 OAI21_X1 _10834_ (.A(_04512_),
    .B1(_04513_),
    .B2(_04505_),
    .ZN(_00439_));
 NAND2_X1 _10835_ (.A1(_01209_),
    .A2(_04496_),
    .ZN(_04514_));
 NAND2_X1 _10836_ (.A1(_04499_),
    .A2(\registers[10][23] ),
    .ZN(_04515_));
 OAI21_X1 _10837_ (.A(_04514_),
    .B1(_04515_),
    .B2(_04505_),
    .ZN(_00440_));
 NAND2_X1 _10838_ (.A1(_01213_),
    .A2(_04496_),
    .ZN(_04516_));
 NAND2_X1 _10839_ (.A1(_04499_),
    .A2(\registers[10][24] ),
    .ZN(_04517_));
 OAI21_X1 _10840_ (.A(_04516_),
    .B1(_04517_),
    .B2(_04505_),
    .ZN(_00441_));
 NAND2_X1 _10841_ (.A1(_01217_),
    .A2(_04496_),
    .ZN(_04518_));
 NAND2_X1 _10842_ (.A1(_04499_),
    .A2(\registers[10][25] ),
    .ZN(_04519_));
 OAI21_X1 _10843_ (.A(_04518_),
    .B1(_04519_),
    .B2(_04505_),
    .ZN(_00442_));
 CLKBUF_X3 _10844_ (.A(_04477_),
    .Z(_04520_));
 NAND2_X1 _10845_ (.A1(_01221_),
    .A2(_04520_),
    .ZN(_04521_));
 CLKBUF_X3 _10846_ (.A(_04498_),
    .Z(_04522_));
 NAND2_X1 _10847_ (.A1(_04522_),
    .A2(\registers[10][26] ),
    .ZN(_04523_));
 OAI21_X1 _10848_ (.A(_04521_),
    .B1(_04523_),
    .B2(_04505_),
    .ZN(_00443_));
 NAND2_X1 _10849_ (.A1(_01226_),
    .A2(_04520_),
    .ZN(_04524_));
 NAND2_X1 _10850_ (.A1(_04522_),
    .A2(\registers[10][27] ),
    .ZN(_04525_));
 OAI21_X1 _10851_ (.A(_04524_),
    .B1(_04525_),
    .B2(_04505_),
    .ZN(_00444_));
 NAND2_X1 _10852_ (.A1(_01230_),
    .A2(_04520_),
    .ZN(_04526_));
 NAND2_X1 _10853_ (.A1(_04522_),
    .A2(\registers[10][28] ),
    .ZN(_04527_));
 CLKBUF_X3 _10854_ (.A(_04477_),
    .Z(_04528_));
 OAI21_X1 _10855_ (.A(_04526_),
    .B1(_04527_),
    .B2(_04528_),
    .ZN(_00445_));
 NAND2_X1 _10856_ (.A1(_01235_),
    .A2(_04520_),
    .ZN(_04529_));
 NAND2_X1 _10857_ (.A1(_04522_),
    .A2(\registers[10][29] ),
    .ZN(_04530_));
 OAI21_X1 _10858_ (.A(_04529_),
    .B1(_04530_),
    .B2(_04528_),
    .ZN(_00446_));
 NAND2_X1 _10859_ (.A1(_01239_),
    .A2(_04520_),
    .ZN(_04531_));
 NAND2_X1 _10860_ (.A1(_04522_),
    .A2(\registers[10][2] ),
    .ZN(_04532_));
 OAI21_X1 _10861_ (.A(_04531_),
    .B1(_04532_),
    .B2(_04528_),
    .ZN(_00447_));
 NAND2_X1 _10862_ (.A1(_01244_),
    .A2(_04520_),
    .ZN(_04533_));
 NAND2_X1 _10863_ (.A1(_04522_),
    .A2(\registers[10][30] ),
    .ZN(_04534_));
 OAI21_X1 _10864_ (.A(_04533_),
    .B1(_04534_),
    .B2(_04528_),
    .ZN(_00448_));
 NAND2_X1 _10865_ (.A1(_01089_),
    .A2(_04520_),
    .ZN(_04535_));
 NAND2_X1 _10866_ (.A1(_04522_),
    .A2(\registers[10][31] ),
    .ZN(_04536_));
 OAI21_X1 _10867_ (.A(_04535_),
    .B1(_04536_),
    .B2(_04528_),
    .ZN(_00449_));
 NAND2_X1 _10868_ (.A1(_01109_),
    .A2(_04520_),
    .ZN(_04537_));
 NAND2_X1 _10869_ (.A1(_04522_),
    .A2(\registers[10][3] ),
    .ZN(_04538_));
 OAI21_X1 _10870_ (.A(_04537_),
    .B1(_04538_),
    .B2(_04528_),
    .ZN(_00450_));
 NAND2_X1 _10871_ (.A1(_01113_),
    .A2(_04520_),
    .ZN(_04539_));
 NAND2_X1 _10872_ (.A1(_04522_),
    .A2(\registers[10][4] ),
    .ZN(_04540_));
 OAI21_X1 _10873_ (.A(_04539_),
    .B1(_04540_),
    .B2(_04528_),
    .ZN(_00451_));
 NAND2_X1 _10874_ (.A1(_01117_),
    .A2(_04520_),
    .ZN(_04541_));
 NAND2_X1 _10875_ (.A1(_04522_),
    .A2(\registers[10][5] ),
    .ZN(_04542_));
 OAI21_X1 _10876_ (.A(_04541_),
    .B1(_04542_),
    .B2(_04528_),
    .ZN(_00452_));
 NAND2_X1 _10877_ (.A1(_01121_),
    .A2(_04477_),
    .ZN(_04543_));
 BUF_X4 _10878_ (.A(_04498_),
    .Z(_04544_));
 NAND2_X1 _10879_ (.A1(_04544_),
    .A2(\registers[10][6] ),
    .ZN(_04545_));
 OAI21_X1 _10880_ (.A(_04543_),
    .B1(_04545_),
    .B2(_04528_),
    .ZN(_00453_));
 NAND2_X1 _10881_ (.A1(_01125_),
    .A2(_04477_),
    .ZN(_04546_));
 NAND2_X1 _10882_ (.A1(_04544_),
    .A2(\registers[10][7] ),
    .ZN(_04547_));
 OAI21_X1 _10883_ (.A(_04546_),
    .B1(_04547_),
    .B2(_04528_),
    .ZN(_00454_));
 NAND2_X1 _10884_ (.A1(_01129_),
    .A2(_04477_),
    .ZN(_04548_));
 NAND2_X1 _10885_ (.A1(_04544_),
    .A2(\registers[10][8] ),
    .ZN(_04549_));
 OAI21_X1 _10886_ (.A(_04548_),
    .B1(_04549_),
    .B2(_04478_),
    .ZN(_00455_));
 NAND2_X1 _10887_ (.A1(_01133_),
    .A2(_04477_),
    .ZN(_04550_));
 NAND2_X1 _10888_ (.A1(_04544_),
    .A2(\registers[10][9] ),
    .ZN(_04551_));
 OAI21_X1 _10889_ (.A(_04550_),
    .B1(_04551_),
    .B2(_04478_),
    .ZN(_00456_));
 OR2_X1 _10890_ (.A1(_01340_),
    .A2(_01739_),
    .ZN(_04552_));
 BUF_X4 _10891_ (.A(_04552_),
    .Z(_04553_));
 BUF_X4 _10892_ (.A(_04553_),
    .Z(_04554_));
 NAND3_X1 _10893_ (.A1(_01774_),
    .A2(\registers[11][0] ),
    .A3(_04554_),
    .ZN(_04555_));
 CLKBUF_X3 _10894_ (.A(_04553_),
    .Z(_04556_));
 OAI21_X1 _10895_ (.A(_04555_),
    .B1(_04556_),
    .B2(_01424_),
    .ZN(_00457_));
 NAND3_X1 _10896_ (.A1(_01774_),
    .A2(\registers[11][10] ),
    .A3(_04554_),
    .ZN(_04557_));
 OAI21_X1 _10897_ (.A(_04557_),
    .B1(_04556_),
    .B2(_01426_),
    .ZN(_00458_));
 CLKBUF_X3 _10898_ (.A(_01536_),
    .Z(_04558_));
 NAND3_X1 _10899_ (.A1(_04558_),
    .A2(\registers[11][11] ),
    .A3(_04554_),
    .ZN(_04559_));
 OAI21_X1 _10900_ (.A(_04559_),
    .B1(_04556_),
    .B2(_01428_),
    .ZN(_00459_));
 NAND3_X1 _10901_ (.A1(_04558_),
    .A2(\registers[11][12] ),
    .A3(_04554_),
    .ZN(_04560_));
 OAI21_X1 _10902_ (.A(_04560_),
    .B1(_04556_),
    .B2(_01430_),
    .ZN(_00460_));
 NAND3_X1 _10903_ (.A1(_04558_),
    .A2(\registers[11][13] ),
    .A3(_04554_),
    .ZN(_04561_));
 OAI21_X1 _10904_ (.A(_04561_),
    .B1(_04556_),
    .B2(_01432_),
    .ZN(_00461_));
 NAND3_X1 _10905_ (.A1(_04558_),
    .A2(\registers[11][14] ),
    .A3(_04554_),
    .ZN(_04562_));
 OAI21_X1 _10906_ (.A(_04562_),
    .B1(_04556_),
    .B2(_01434_),
    .ZN(_00462_));
 NAND3_X1 _10907_ (.A1(_04558_),
    .A2(\registers[11][15] ),
    .A3(_04554_),
    .ZN(_04563_));
 OAI21_X1 _10908_ (.A(_04563_),
    .B1(_04556_),
    .B2(_01436_),
    .ZN(_00463_));
 NAND3_X1 _10909_ (.A1(_04558_),
    .A2(\registers[11][16] ),
    .A3(_04554_),
    .ZN(_04564_));
 OAI21_X1 _10910_ (.A(_04564_),
    .B1(_04556_),
    .B2(_01438_),
    .ZN(_00464_));
 CLKBUF_X3 _10911_ (.A(_04553_),
    .Z(_04565_));
 NAND3_X1 _10912_ (.A1(_04558_),
    .A2(\registers[11][17] ),
    .A3(_04565_),
    .ZN(_04566_));
 OAI21_X1 _10913_ (.A(_04566_),
    .B1(_04556_),
    .B2(_01441_),
    .ZN(_00465_));
 NAND3_X1 _10914_ (.A1(_04558_),
    .A2(\registers[11][18] ),
    .A3(_04565_),
    .ZN(_04567_));
 OAI21_X1 _10915_ (.A(_04567_),
    .B1(_04556_),
    .B2(_01443_),
    .ZN(_00466_));
 NAND3_X1 _10916_ (.A1(_04558_),
    .A2(\registers[11][19] ),
    .A3(_04565_),
    .ZN(_04568_));
 CLKBUF_X3 _10917_ (.A(_04553_),
    .Z(_04569_));
 OAI21_X1 _10918_ (.A(_04568_),
    .B1(_04569_),
    .B2(_01447_),
    .ZN(_00467_));
 NAND3_X1 _10919_ (.A1(_04558_),
    .A2(\registers[11][1] ),
    .A3(_04565_),
    .ZN(_04570_));
 OAI21_X1 _10920_ (.A(_04570_),
    .B1(_04569_),
    .B2(_01449_),
    .ZN(_00468_));
 CLKBUF_X3 _10921_ (.A(_01536_),
    .Z(_04571_));
 NAND3_X1 _10922_ (.A1(_04571_),
    .A2(\registers[11][20] ),
    .A3(_04565_),
    .ZN(_04572_));
 OAI21_X1 _10923_ (.A(_04572_),
    .B1(_04569_),
    .B2(_01451_),
    .ZN(_00469_));
 NAND3_X1 _10924_ (.A1(_04571_),
    .A2(\registers[11][21] ),
    .A3(_04565_),
    .ZN(_04573_));
 OAI21_X1 _10925_ (.A(_04573_),
    .B1(_04569_),
    .B2(_01453_),
    .ZN(_00470_));
 NAND3_X1 _10926_ (.A1(_04571_),
    .A2(\registers[11][22] ),
    .A3(_04565_),
    .ZN(_04574_));
 OAI21_X1 _10927_ (.A(_04574_),
    .B1(_04569_),
    .B2(_01455_),
    .ZN(_00471_));
 NAND3_X1 _10928_ (.A1(_04571_),
    .A2(\registers[11][23] ),
    .A3(_04565_),
    .ZN(_04575_));
 OAI21_X1 _10929_ (.A(_04575_),
    .B1(_04569_),
    .B2(_01457_),
    .ZN(_00472_));
 NAND3_X1 _10930_ (.A1(_04571_),
    .A2(\registers[11][24] ),
    .A3(_04565_),
    .ZN(_04576_));
 OAI21_X1 _10931_ (.A(_04576_),
    .B1(_04569_),
    .B2(_01459_),
    .ZN(_00473_));
 NAND3_X1 _10932_ (.A1(_04571_),
    .A2(\registers[11][25] ),
    .A3(_04565_),
    .ZN(_04577_));
 OAI21_X1 _10933_ (.A(_04577_),
    .B1(_04569_),
    .B2(_01461_),
    .ZN(_00474_));
 CLKBUF_X3 _10934_ (.A(_04553_),
    .Z(_04578_));
 NAND3_X1 _10935_ (.A1(_04571_),
    .A2(\registers[11][26] ),
    .A3(_04578_),
    .ZN(_04579_));
 OAI21_X1 _10936_ (.A(_04579_),
    .B1(_04569_),
    .B2(_01464_),
    .ZN(_00475_));
 NAND3_X1 _10937_ (.A1(_04571_),
    .A2(\registers[11][27] ),
    .A3(_04578_),
    .ZN(_04580_));
 OAI21_X1 _10938_ (.A(_04580_),
    .B1(_04569_),
    .B2(_01466_),
    .ZN(_00476_));
 NAND3_X1 _10939_ (.A1(_04571_),
    .A2(\registers[11][28] ),
    .A3(_04578_),
    .ZN(_04581_));
 CLKBUF_X3 _10940_ (.A(_04553_),
    .Z(_04582_));
 OAI21_X1 _10941_ (.A(_04581_),
    .B1(_04582_),
    .B2(_01470_),
    .ZN(_00477_));
 NAND3_X1 _10942_ (.A1(_04571_),
    .A2(\registers[11][29] ),
    .A3(_04578_),
    .ZN(_04583_));
 OAI21_X1 _10943_ (.A(_04583_),
    .B1(_04582_),
    .B2(_01472_),
    .ZN(_00478_));
 BUF_X4 _10944_ (.A(_01536_),
    .Z(_04584_));
 NAND3_X1 _10945_ (.A1(_04584_),
    .A2(\registers[11][2] ),
    .A3(_04578_),
    .ZN(_04585_));
 OAI21_X1 _10946_ (.A(_04585_),
    .B1(_04582_),
    .B2(_01474_),
    .ZN(_00479_));
 NAND3_X1 _10947_ (.A1(_04584_),
    .A2(\registers[11][30] ),
    .A3(_04578_),
    .ZN(_04586_));
 OAI21_X1 _10948_ (.A(_04586_),
    .B1(_04582_),
    .B2(_01476_),
    .ZN(_00480_));
 NAND3_X1 _10949_ (.A1(_04584_),
    .A2(\registers[11][31] ),
    .A3(_04578_),
    .ZN(_04587_));
 OAI21_X1 _10950_ (.A(_04587_),
    .B1(_04582_),
    .B2(_01478_),
    .ZN(_00481_));
 NAND3_X1 _10951_ (.A1(_04584_),
    .A2(\registers[11][3] ),
    .A3(_04578_),
    .ZN(_04588_));
 OAI21_X1 _10952_ (.A(_04588_),
    .B1(_04582_),
    .B2(_01480_),
    .ZN(_00482_));
 NAND3_X1 _10953_ (.A1(_04584_),
    .A2(\registers[11][4] ),
    .A3(_04578_),
    .ZN(_04589_));
 OAI21_X1 _10954_ (.A(_04589_),
    .B1(_04582_),
    .B2(_01482_),
    .ZN(_00483_));
 NAND3_X1 _10955_ (.A1(_04584_),
    .A2(\registers[11][5] ),
    .A3(_04578_),
    .ZN(_04590_));
 OAI21_X1 _10956_ (.A(_04590_),
    .B1(_04582_),
    .B2(_01484_),
    .ZN(_00484_));
 NAND3_X1 _10957_ (.A1(_04584_),
    .A2(\registers[11][6] ),
    .A3(_04553_),
    .ZN(_04591_));
 OAI21_X1 _10958_ (.A(_04591_),
    .B1(_04582_),
    .B2(_01486_),
    .ZN(_00485_));
 NAND3_X1 _10959_ (.A1(_04584_),
    .A2(\registers[11][7] ),
    .A3(_04553_),
    .ZN(_04592_));
 OAI21_X1 _10960_ (.A(_04592_),
    .B1(_04582_),
    .B2(_01488_),
    .ZN(_00486_));
 NAND3_X1 _10961_ (.A1(_04584_),
    .A2(\registers[11][8] ),
    .A3(_04553_),
    .ZN(_04593_));
 OAI21_X1 _10962_ (.A(_04593_),
    .B1(_04554_),
    .B2(_01491_),
    .ZN(_00487_));
 NAND3_X1 _10963_ (.A1(_04584_),
    .A2(\registers[11][9] ),
    .A3(_04553_),
    .ZN(_04594_));
 OAI21_X1 _10964_ (.A(_04594_),
    .B1(_04554_),
    .B2(_01493_),
    .ZN(_00488_));
 BUF_X4 _10965_ (.A(_01103_),
    .Z(_04595_));
 CLKBUF_X3 _10966_ (.A(_04595_),
    .Z(_04596_));
 NAND3_X2 _10967_ (.A1(_01090_),
    .A2(_01738_),
    .A3(_01092_),
    .ZN(_04597_));
 OR2_X1 _10968_ (.A1(_01737_),
    .A2(_04597_),
    .ZN(_04598_));
 BUF_X4 _10969_ (.A(_04598_),
    .Z(_04599_));
 CLKBUF_X3 _10970_ (.A(_04599_),
    .Z(_04600_));
 NAND3_X1 _10971_ (.A1(_04596_),
    .A2(\registers[12][0] ),
    .A3(_04600_),
    .ZN(_04601_));
 CLKBUF_X3 _10972_ (.A(_04599_),
    .Z(_04602_));
 OAI21_X1 _10973_ (.A(_04601_),
    .B1(_04602_),
    .B2(_01424_),
    .ZN(_00489_));
 NAND3_X1 _10974_ (.A1(_04596_),
    .A2(\registers[12][10] ),
    .A3(_04600_),
    .ZN(_04603_));
 OAI21_X1 _10975_ (.A(_04603_),
    .B1(_04602_),
    .B2(_01426_),
    .ZN(_00490_));
 NAND3_X1 _10976_ (.A1(_04596_),
    .A2(\registers[12][11] ),
    .A3(_04600_),
    .ZN(_04604_));
 OAI21_X1 _10977_ (.A(_04604_),
    .B1(_04602_),
    .B2(_01428_),
    .ZN(_00491_));
 NAND3_X1 _10978_ (.A1(_04596_),
    .A2(\registers[12][12] ),
    .A3(_04600_),
    .ZN(_04605_));
 OAI21_X1 _10979_ (.A(_04605_),
    .B1(_04602_),
    .B2(_01430_),
    .ZN(_00492_));
 NAND3_X1 _10980_ (.A1(_04596_),
    .A2(\registers[12][13] ),
    .A3(_04600_),
    .ZN(_04606_));
 OAI21_X1 _10981_ (.A(_04606_),
    .B1(_04602_),
    .B2(_01432_),
    .ZN(_00493_));
 NAND3_X1 _10982_ (.A1(_04596_),
    .A2(\registers[12][14] ),
    .A3(_04600_),
    .ZN(_04607_));
 OAI21_X1 _10983_ (.A(_04607_),
    .B1(_04602_),
    .B2(_01434_),
    .ZN(_00494_));
 NAND3_X1 _10984_ (.A1(_04596_),
    .A2(\registers[12][15] ),
    .A3(_04600_),
    .ZN(_04608_));
 OAI21_X1 _10985_ (.A(_04608_),
    .B1(_04602_),
    .B2(_01436_),
    .ZN(_00495_));
 NAND3_X1 _10986_ (.A1(_04596_),
    .A2(\registers[12][16] ),
    .A3(_04600_),
    .ZN(_04609_));
 OAI21_X1 _10987_ (.A(_04609_),
    .B1(_04602_),
    .B2(_01438_),
    .ZN(_00496_));
 CLKBUF_X3 _10988_ (.A(_04599_),
    .Z(_04610_));
 NAND3_X1 _10989_ (.A1(_04596_),
    .A2(\registers[12][17] ),
    .A3(_04610_),
    .ZN(_04611_));
 OAI21_X1 _10990_ (.A(_04611_),
    .B1(_04602_),
    .B2(_01441_),
    .ZN(_00497_));
 NAND3_X1 _10991_ (.A1(_04596_),
    .A2(\registers[12][18] ),
    .A3(_04610_),
    .ZN(_04612_));
 OAI21_X1 _10992_ (.A(_04612_),
    .B1(_04602_),
    .B2(_01443_),
    .ZN(_00498_));
 CLKBUF_X3 _10993_ (.A(_04595_),
    .Z(_04613_));
 NAND3_X1 _10994_ (.A1(_04613_),
    .A2(\registers[12][19] ),
    .A3(_04610_),
    .ZN(_04614_));
 CLKBUF_X3 _10995_ (.A(_04599_),
    .Z(_04615_));
 OAI21_X1 _10996_ (.A(_04614_),
    .B1(_04615_),
    .B2(_01447_),
    .ZN(_00499_));
 NAND3_X1 _10997_ (.A1(_04613_),
    .A2(\registers[12][1] ),
    .A3(_04610_),
    .ZN(_04616_));
 OAI21_X1 _10998_ (.A(_04616_),
    .B1(_04615_),
    .B2(_01449_),
    .ZN(_00500_));
 NAND3_X1 _10999_ (.A1(_04613_),
    .A2(\registers[12][20] ),
    .A3(_04610_),
    .ZN(_04617_));
 OAI21_X1 _11000_ (.A(_04617_),
    .B1(_04615_),
    .B2(_01451_),
    .ZN(_00501_));
 NAND3_X1 _11001_ (.A1(_04613_),
    .A2(\registers[12][21] ),
    .A3(_04610_),
    .ZN(_04618_));
 OAI21_X1 _11002_ (.A(_04618_),
    .B1(_04615_),
    .B2(_01453_),
    .ZN(_00502_));
 NAND3_X1 _11003_ (.A1(_04613_),
    .A2(\registers[12][22] ),
    .A3(_04610_),
    .ZN(_04619_));
 OAI21_X1 _11004_ (.A(_04619_),
    .B1(_04615_),
    .B2(_01455_),
    .ZN(_00503_));
 NAND3_X1 _11005_ (.A1(_04613_),
    .A2(\registers[12][23] ),
    .A3(_04610_),
    .ZN(_04620_));
 OAI21_X1 _11006_ (.A(_04620_),
    .B1(_04615_),
    .B2(_01457_),
    .ZN(_00504_));
 NAND3_X1 _11007_ (.A1(_04613_),
    .A2(\registers[12][24] ),
    .A3(_04610_),
    .ZN(_04621_));
 OAI21_X1 _11008_ (.A(_04621_),
    .B1(_04615_),
    .B2(_01459_),
    .ZN(_00505_));
 NAND3_X1 _11009_ (.A1(_04613_),
    .A2(\registers[12][25] ),
    .A3(_04610_),
    .ZN(_04622_));
 OAI21_X1 _11010_ (.A(_04622_),
    .B1(_04615_),
    .B2(_01461_),
    .ZN(_00506_));
 CLKBUF_X3 _11011_ (.A(_04599_),
    .Z(_04623_));
 NAND3_X1 _11012_ (.A1(_04613_),
    .A2(\registers[12][26] ),
    .A3(_04623_),
    .ZN(_04624_));
 OAI21_X1 _11013_ (.A(_04624_),
    .B1(_04615_),
    .B2(_01464_),
    .ZN(_00507_));
 NAND3_X1 _11014_ (.A1(_04613_),
    .A2(\registers[12][27] ),
    .A3(_04623_),
    .ZN(_04625_));
 OAI21_X1 _11015_ (.A(_04625_),
    .B1(_04615_),
    .B2(_01466_),
    .ZN(_00508_));
 CLKBUF_X3 _11016_ (.A(_04595_),
    .Z(_04626_));
 NAND3_X1 _11017_ (.A1(_04626_),
    .A2(\registers[12][28] ),
    .A3(_04623_),
    .ZN(_04627_));
 CLKBUF_X3 _11018_ (.A(_04599_),
    .Z(_04628_));
 OAI21_X1 _11019_ (.A(_04627_),
    .B1(_04628_),
    .B2(_01470_),
    .ZN(_00509_));
 NAND3_X1 _11020_ (.A1(_04626_),
    .A2(\registers[12][29] ),
    .A3(_04623_),
    .ZN(_04629_));
 OAI21_X1 _11021_ (.A(_04629_),
    .B1(_04628_),
    .B2(_01472_),
    .ZN(_00510_));
 NAND3_X1 _11022_ (.A1(_04626_),
    .A2(\registers[12][2] ),
    .A3(_04623_),
    .ZN(_04630_));
 OAI21_X1 _11023_ (.A(_04630_),
    .B1(_04628_),
    .B2(_01474_),
    .ZN(_00511_));
 NAND3_X1 _11024_ (.A1(_04626_),
    .A2(\registers[12][30] ),
    .A3(_04623_),
    .ZN(_04631_));
 OAI21_X1 _11025_ (.A(_04631_),
    .B1(_04628_),
    .B2(_01476_),
    .ZN(_00512_));
 NAND3_X1 _11026_ (.A1(_04626_),
    .A2(\registers[12][31] ),
    .A3(_04623_),
    .ZN(_04632_));
 OAI21_X1 _11027_ (.A(_04632_),
    .B1(_04628_),
    .B2(_01478_),
    .ZN(_00513_));
 NAND3_X1 _11028_ (.A1(_04626_),
    .A2(\registers[12][3] ),
    .A3(_04623_),
    .ZN(_04633_));
 OAI21_X1 _11029_ (.A(_04633_),
    .B1(_04628_),
    .B2(_01480_),
    .ZN(_00514_));
 NAND3_X1 _11030_ (.A1(_04626_),
    .A2(\registers[12][4] ),
    .A3(_04623_),
    .ZN(_04634_));
 OAI21_X1 _11031_ (.A(_04634_),
    .B1(_04628_),
    .B2(_01482_),
    .ZN(_00515_));
 NAND3_X1 _11032_ (.A1(_04626_),
    .A2(\registers[12][5] ),
    .A3(_04623_),
    .ZN(_04635_));
 OAI21_X1 _11033_ (.A(_04635_),
    .B1(_04628_),
    .B2(_01484_),
    .ZN(_00516_));
 NAND3_X1 _11034_ (.A1(_04626_),
    .A2(\registers[12][6] ),
    .A3(_04599_),
    .ZN(_04636_));
 OAI21_X1 _11035_ (.A(_04636_),
    .B1(_04628_),
    .B2(_01486_),
    .ZN(_00517_));
 NAND3_X1 _11036_ (.A1(_04626_),
    .A2(\registers[12][7] ),
    .A3(_04599_),
    .ZN(_04637_));
 OAI21_X1 _11037_ (.A(_04637_),
    .B1(_04628_),
    .B2(_01488_),
    .ZN(_00518_));
 BUF_X4 _11038_ (.A(_04595_),
    .Z(_04638_));
 NAND3_X1 _11039_ (.A1(_04638_),
    .A2(\registers[12][8] ),
    .A3(_04599_),
    .ZN(_04639_));
 OAI21_X1 _11040_ (.A(_04639_),
    .B1(_04600_),
    .B2(_01491_),
    .ZN(_00519_));
 NAND3_X1 _11041_ (.A1(_04638_),
    .A2(\registers[12][9] ),
    .A3(_04599_),
    .ZN(_04640_));
 OAI21_X1 _11042_ (.A(_04640_),
    .B1(_04600_),
    .B2(_01493_),
    .ZN(_00520_));
 NOR2_X1 _11043_ (.A1(_01098_),
    .A2(_04597_),
    .ZN(_04641_));
 CLKBUF_X3 _11044_ (.A(_04641_),
    .Z(_04642_));
 CLKBUF_X3 _11045_ (.A(_04642_),
    .Z(_04643_));
 NAND2_X1 _11046_ (.A1(_01137_),
    .A2(_04643_),
    .ZN(_04644_));
 NAND2_X1 _11047_ (.A1(_04544_),
    .A2(\registers[13][0] ),
    .ZN(_04645_));
 CLKBUF_X3 _11048_ (.A(_04642_),
    .Z(_04646_));
 OAI21_X1 _11049_ (.A(_04644_),
    .B1(_04645_),
    .B2(_04646_),
    .ZN(_00521_));
 NAND2_X1 _11050_ (.A1(_01149_),
    .A2(_04643_),
    .ZN(_04647_));
 NAND2_X1 _11051_ (.A1(_04544_),
    .A2(\registers[13][10] ),
    .ZN(_04648_));
 OAI21_X1 _11052_ (.A(_04647_),
    .B1(_04648_),
    .B2(_04646_),
    .ZN(_00522_));
 NAND2_X1 _11053_ (.A1(_01153_),
    .A2(_04643_),
    .ZN(_04649_));
 NAND2_X1 _11054_ (.A1(_04544_),
    .A2(\registers[13][11] ),
    .ZN(_04650_));
 OAI21_X1 _11055_ (.A(_04649_),
    .B1(_04650_),
    .B2(_04646_),
    .ZN(_00523_));
 NAND2_X1 _11056_ (.A1(_01158_),
    .A2(_04643_),
    .ZN(_04651_));
 NAND2_X1 _11057_ (.A1(_04544_),
    .A2(\registers[13][12] ),
    .ZN(_04652_));
 OAI21_X1 _11058_ (.A(_04651_),
    .B1(_04652_),
    .B2(_04646_),
    .ZN(_00524_));
 NAND2_X1 _11059_ (.A1(_01162_),
    .A2(_04643_),
    .ZN(_04653_));
 NAND2_X1 _11060_ (.A1(_04544_),
    .A2(\registers[13][13] ),
    .ZN(_04654_));
 OAI21_X1 _11061_ (.A(_04653_),
    .B1(_04654_),
    .B2(_04646_),
    .ZN(_00525_));
 NAND2_X1 _11062_ (.A1(_01166_),
    .A2(_04643_),
    .ZN(_04655_));
 NAND2_X1 _11063_ (.A1(_04544_),
    .A2(\registers[13][14] ),
    .ZN(_04656_));
 OAI21_X1 _11064_ (.A(_04655_),
    .B1(_04656_),
    .B2(_04646_),
    .ZN(_00526_));
 NAND2_X1 _11065_ (.A1(_01170_),
    .A2(_04643_),
    .ZN(_04657_));
 CLKBUF_X3 _11066_ (.A(_04498_),
    .Z(_04658_));
 NAND2_X1 _11067_ (.A1(_04658_),
    .A2(\registers[13][15] ),
    .ZN(_04659_));
 OAI21_X1 _11068_ (.A(_04657_),
    .B1(_04659_),
    .B2(_04646_),
    .ZN(_00527_));
 NAND2_X1 _11069_ (.A1(_01174_),
    .A2(_04643_),
    .ZN(_04660_));
 NAND2_X1 _11070_ (.A1(_04658_),
    .A2(\registers[13][16] ),
    .ZN(_04661_));
 OAI21_X1 _11071_ (.A(_04660_),
    .B1(_04661_),
    .B2(_04646_),
    .ZN(_00528_));
 CLKBUF_X3 _11072_ (.A(_04642_),
    .Z(_04662_));
 NAND2_X1 _11073_ (.A1(_01178_),
    .A2(_04662_),
    .ZN(_04663_));
 NAND2_X1 _11074_ (.A1(_04658_),
    .A2(\registers[13][17] ),
    .ZN(_04664_));
 OAI21_X1 _11075_ (.A(_04663_),
    .B1(_04664_),
    .B2(_04646_),
    .ZN(_00529_));
 NAND2_X1 _11076_ (.A1(_01183_),
    .A2(_04662_),
    .ZN(_04665_));
 NAND2_X1 _11077_ (.A1(_04658_),
    .A2(\registers[13][18] ),
    .ZN(_04666_));
 OAI21_X1 _11078_ (.A(_04665_),
    .B1(_04666_),
    .B2(_04646_),
    .ZN(_00530_));
 NAND2_X1 _11079_ (.A1(_01187_),
    .A2(_04662_),
    .ZN(_04667_));
 NAND2_X1 _11080_ (.A1(_04658_),
    .A2(\registers[13][19] ),
    .ZN(_04668_));
 CLKBUF_X3 _11081_ (.A(_04642_),
    .Z(_04669_));
 OAI21_X1 _11082_ (.A(_04667_),
    .B1(_04668_),
    .B2(_04669_),
    .ZN(_00531_));
 NAND2_X1 _11083_ (.A1(_01192_),
    .A2(_04662_),
    .ZN(_04670_));
 NAND2_X1 _11084_ (.A1(_04658_),
    .A2(\registers[13][1] ),
    .ZN(_04671_));
 OAI21_X1 _11085_ (.A(_04670_),
    .B1(_04671_),
    .B2(_04669_),
    .ZN(_00532_));
 NAND2_X1 _11086_ (.A1(_01196_),
    .A2(_04662_),
    .ZN(_04672_));
 NAND2_X1 _11087_ (.A1(_04658_),
    .A2(\registers[13][20] ),
    .ZN(_04673_));
 OAI21_X1 _11088_ (.A(_04672_),
    .B1(_04673_),
    .B2(_04669_),
    .ZN(_00533_));
 NAND2_X1 _11089_ (.A1(_01201_),
    .A2(_04662_),
    .ZN(_04674_));
 NAND2_X1 _11090_ (.A1(_04658_),
    .A2(\registers[13][21] ),
    .ZN(_04675_));
 OAI21_X1 _11091_ (.A(_04674_),
    .B1(_04675_),
    .B2(_04669_),
    .ZN(_00534_));
 NAND2_X1 _11092_ (.A1(_01205_),
    .A2(_04662_),
    .ZN(_04676_));
 NAND2_X1 _11093_ (.A1(_04658_),
    .A2(\registers[13][22] ),
    .ZN(_04677_));
 OAI21_X1 _11094_ (.A(_04676_),
    .B1(_04677_),
    .B2(_04669_),
    .ZN(_00535_));
 NAND2_X1 _11095_ (.A1(_01209_),
    .A2(_04662_),
    .ZN(_04678_));
 NAND2_X1 _11096_ (.A1(_04658_),
    .A2(\registers[13][23] ),
    .ZN(_04679_));
 OAI21_X1 _11097_ (.A(_04678_),
    .B1(_04679_),
    .B2(_04669_),
    .ZN(_00536_));
 NAND2_X1 _11098_ (.A1(_01213_),
    .A2(_04662_),
    .ZN(_04680_));
 CLKBUF_X3 _11099_ (.A(_04498_),
    .Z(_04681_));
 NAND2_X1 _11100_ (.A1(_04681_),
    .A2(\registers[13][24] ),
    .ZN(_04682_));
 OAI21_X1 _11101_ (.A(_04680_),
    .B1(_04682_),
    .B2(_04669_),
    .ZN(_00537_));
 NAND2_X1 _11102_ (.A1(_01217_),
    .A2(_04662_),
    .ZN(_04683_));
 NAND2_X1 _11103_ (.A1(_04681_),
    .A2(\registers[13][25] ),
    .ZN(_04684_));
 OAI21_X1 _11104_ (.A(_04683_),
    .B1(_04684_),
    .B2(_04669_),
    .ZN(_00538_));
 CLKBUF_X3 _11105_ (.A(_04642_),
    .Z(_04685_));
 NAND2_X1 _11106_ (.A1(_01221_),
    .A2(_04685_),
    .ZN(_04686_));
 NAND2_X1 _11107_ (.A1(_04681_),
    .A2(\registers[13][26] ),
    .ZN(_04687_));
 OAI21_X1 _11108_ (.A(_04686_),
    .B1(_04687_),
    .B2(_04669_),
    .ZN(_00539_));
 NAND2_X1 _11109_ (.A1(_01226_),
    .A2(_04685_),
    .ZN(_04688_));
 NAND2_X1 _11110_ (.A1(_04681_),
    .A2(\registers[13][27] ),
    .ZN(_04689_));
 OAI21_X1 _11111_ (.A(_04688_),
    .B1(_04689_),
    .B2(_04669_),
    .ZN(_00540_));
 NAND2_X1 _11112_ (.A1(_01230_),
    .A2(_04685_),
    .ZN(_04690_));
 NAND2_X1 _11113_ (.A1(_04681_),
    .A2(\registers[13][28] ),
    .ZN(_04691_));
 CLKBUF_X3 _11114_ (.A(_04642_),
    .Z(_04692_));
 OAI21_X1 _11115_ (.A(_04690_),
    .B1(_04691_),
    .B2(_04692_),
    .ZN(_00541_));
 NAND2_X1 _11116_ (.A1(_01235_),
    .A2(_04685_),
    .ZN(_04693_));
 NAND2_X1 _11117_ (.A1(_04681_),
    .A2(\registers[13][29] ),
    .ZN(_04694_));
 OAI21_X1 _11118_ (.A(_04693_),
    .B1(_04694_),
    .B2(_04692_),
    .ZN(_00542_));
 NAND2_X1 _11119_ (.A1(_01239_),
    .A2(_04685_),
    .ZN(_04695_));
 NAND2_X1 _11120_ (.A1(_04681_),
    .A2(\registers[13][2] ),
    .ZN(_04696_));
 OAI21_X1 _11121_ (.A(_04695_),
    .B1(_04696_),
    .B2(_04692_),
    .ZN(_00543_));
 NAND2_X1 _11122_ (.A1(_01244_),
    .A2(_04685_),
    .ZN(_04697_));
 NAND2_X1 _11123_ (.A1(_04681_),
    .A2(\registers[13][30] ),
    .ZN(_04698_));
 OAI21_X1 _11124_ (.A(_04697_),
    .B1(_04698_),
    .B2(_04692_),
    .ZN(_00544_));
 NAND2_X1 _11125_ (.A1(_01089_),
    .A2(_04685_),
    .ZN(_04699_));
 NAND2_X1 _11126_ (.A1(_04681_),
    .A2(\registers[13][31] ),
    .ZN(_04700_));
 OAI21_X1 _11127_ (.A(_04699_),
    .B1(_04700_),
    .B2(_04692_),
    .ZN(_00545_));
 NAND2_X1 _11128_ (.A1(_01109_),
    .A2(_04685_),
    .ZN(_04701_));
 NAND2_X1 _11129_ (.A1(_04681_),
    .A2(\registers[13][3] ),
    .ZN(_04702_));
 OAI21_X1 _11130_ (.A(_04701_),
    .B1(_04702_),
    .B2(_04692_),
    .ZN(_00546_));
 NAND2_X1 _11131_ (.A1(_01113_),
    .A2(_04685_),
    .ZN(_04703_));
 BUF_X4 _11132_ (.A(_04498_),
    .Z(_04704_));
 NAND2_X1 _11133_ (.A1(_04704_),
    .A2(\registers[13][4] ),
    .ZN(_04705_));
 OAI21_X1 _11134_ (.A(_04703_),
    .B1(_04705_),
    .B2(_04692_),
    .ZN(_00547_));
 NAND2_X1 _11135_ (.A1(_01117_),
    .A2(_04685_),
    .ZN(_04706_));
 NAND2_X1 _11136_ (.A1(_04704_),
    .A2(\registers[13][5] ),
    .ZN(_04707_));
 OAI21_X1 _11137_ (.A(_04706_),
    .B1(_04707_),
    .B2(_04692_),
    .ZN(_00548_));
 NAND2_X1 _11138_ (.A1(_01121_),
    .A2(_04642_),
    .ZN(_04708_));
 NAND2_X1 _11139_ (.A1(_04704_),
    .A2(\registers[13][6] ),
    .ZN(_04709_));
 OAI21_X1 _11140_ (.A(_04708_),
    .B1(_04709_),
    .B2(_04692_),
    .ZN(_00549_));
 NAND2_X1 _11141_ (.A1(_01125_),
    .A2(_04642_),
    .ZN(_04710_));
 NAND2_X1 _11142_ (.A1(_04704_),
    .A2(\registers[13][7] ),
    .ZN(_04711_));
 OAI21_X1 _11143_ (.A(_04710_),
    .B1(_04711_),
    .B2(_04692_),
    .ZN(_00550_));
 NAND2_X1 _11144_ (.A1(_01129_),
    .A2(_04642_),
    .ZN(_04712_));
 NAND2_X1 _11145_ (.A1(_04704_),
    .A2(\registers[13][8] ),
    .ZN(_04713_));
 OAI21_X1 _11146_ (.A(_04712_),
    .B1(_04713_),
    .B2(_04643_),
    .ZN(_00551_));
 NAND2_X1 _11147_ (.A1(_01133_),
    .A2(_04642_),
    .ZN(_04714_));
 NAND2_X1 _11148_ (.A1(_04704_),
    .A2(\registers[13][9] ),
    .ZN(_04715_));
 OAI21_X1 _11149_ (.A(_04714_),
    .B1(_04715_),
    .B2(_04643_),
    .ZN(_00552_));
 NOR2_X1 _11150_ (.A1(_01141_),
    .A2(_04597_),
    .ZN(_04716_));
 BUF_X4 _11151_ (.A(_04716_),
    .Z(_04717_));
 CLKBUF_X3 _11152_ (.A(_04717_),
    .Z(_04718_));
 NAND2_X1 _11153_ (.A1(_01137_),
    .A2(_04718_),
    .ZN(_04719_));
 NAND2_X1 _11154_ (.A1(_04704_),
    .A2(\registers[14][0] ),
    .ZN(_04720_));
 CLKBUF_X3 _11155_ (.A(_04717_),
    .Z(_04721_));
 OAI21_X1 _11156_ (.A(_04719_),
    .B1(_04720_),
    .B2(_04721_),
    .ZN(_00553_));
 NAND2_X1 _11157_ (.A1(_01149_),
    .A2(_04718_),
    .ZN(_04722_));
 NAND2_X1 _11158_ (.A1(_04704_),
    .A2(\registers[14][10] ),
    .ZN(_04723_));
 OAI21_X1 _11159_ (.A(_04722_),
    .B1(_04723_),
    .B2(_04721_),
    .ZN(_00554_));
 NAND2_X1 _11160_ (.A1(_01153_),
    .A2(_04718_),
    .ZN(_04724_));
 NAND2_X1 _11161_ (.A1(_04704_),
    .A2(\registers[14][11] ),
    .ZN(_04725_));
 OAI21_X1 _11162_ (.A(_04724_),
    .B1(_04725_),
    .B2(_04721_),
    .ZN(_00555_));
 NAND2_X1 _11163_ (.A1(_01158_),
    .A2(_04718_),
    .ZN(_04726_));
 NAND2_X1 _11164_ (.A1(_04704_),
    .A2(\registers[14][12] ),
    .ZN(_04727_));
 OAI21_X1 _11165_ (.A(_04726_),
    .B1(_04727_),
    .B2(_04721_),
    .ZN(_00556_));
 NAND2_X1 _11166_ (.A1(_01162_),
    .A2(_04718_),
    .ZN(_04728_));
 CLKBUF_X3 _11167_ (.A(_04498_),
    .Z(_04729_));
 NAND2_X1 _11168_ (.A1(_04729_),
    .A2(\registers[14][13] ),
    .ZN(_04730_));
 OAI21_X1 _11169_ (.A(_04728_),
    .B1(_04730_),
    .B2(_04721_),
    .ZN(_00557_));
 NAND2_X1 _11170_ (.A1(_01166_),
    .A2(_04718_),
    .ZN(_04731_));
 NAND2_X1 _11171_ (.A1(_04729_),
    .A2(\registers[14][14] ),
    .ZN(_04732_));
 OAI21_X1 _11172_ (.A(_04731_),
    .B1(_04732_),
    .B2(_04721_),
    .ZN(_00558_));
 NAND2_X1 _11173_ (.A1(_01170_),
    .A2(_04718_),
    .ZN(_04733_));
 NAND2_X1 _11174_ (.A1(_04729_),
    .A2(\registers[14][15] ),
    .ZN(_04734_));
 OAI21_X1 _11175_ (.A(_04733_),
    .B1(_04734_),
    .B2(_04721_),
    .ZN(_00559_));
 NAND2_X1 _11176_ (.A1(_01174_),
    .A2(_04718_),
    .ZN(_04735_));
 NAND2_X1 _11177_ (.A1(_04729_),
    .A2(\registers[14][16] ),
    .ZN(_04736_));
 OAI21_X1 _11178_ (.A(_04735_),
    .B1(_04736_),
    .B2(_04721_),
    .ZN(_00560_));
 CLKBUF_X3 _11179_ (.A(_04717_),
    .Z(_04737_));
 NAND2_X1 _11180_ (.A1(_01178_),
    .A2(_04737_),
    .ZN(_04738_));
 NAND2_X1 _11181_ (.A1(_04729_),
    .A2(\registers[14][17] ),
    .ZN(_04739_));
 OAI21_X1 _11182_ (.A(_04738_),
    .B1(_04739_),
    .B2(_04721_),
    .ZN(_00561_));
 NAND2_X1 _11183_ (.A1(_01183_),
    .A2(_04737_),
    .ZN(_04740_));
 NAND2_X1 _11184_ (.A1(_04729_),
    .A2(\registers[14][18] ),
    .ZN(_04741_));
 OAI21_X1 _11185_ (.A(_04740_),
    .B1(_04741_),
    .B2(_04721_),
    .ZN(_00562_));
 NAND2_X1 _11186_ (.A1(_01187_),
    .A2(_04737_),
    .ZN(_04742_));
 NAND2_X1 _11187_ (.A1(_04729_),
    .A2(\registers[14][19] ),
    .ZN(_04743_));
 CLKBUF_X3 _11188_ (.A(_04717_),
    .Z(_04744_));
 OAI21_X1 _11189_ (.A(_04742_),
    .B1(_04743_),
    .B2(_04744_),
    .ZN(_00563_));
 NAND2_X1 _11190_ (.A1(_01192_),
    .A2(_04737_),
    .ZN(_04745_));
 NAND2_X1 _11191_ (.A1(_04729_),
    .A2(\registers[14][1] ),
    .ZN(_04746_));
 OAI21_X1 _11192_ (.A(_04745_),
    .B1(_04746_),
    .B2(_04744_),
    .ZN(_00564_));
 NAND2_X1 _11193_ (.A1(_01196_),
    .A2(_04737_),
    .ZN(_04747_));
 NAND2_X1 _11194_ (.A1(_04729_),
    .A2(\registers[14][20] ),
    .ZN(_04748_));
 OAI21_X1 _11195_ (.A(_04747_),
    .B1(_04748_),
    .B2(_04744_),
    .ZN(_00565_));
 NAND2_X1 _11196_ (.A1(_01201_),
    .A2(_04737_),
    .ZN(_04749_));
 NAND2_X1 _11197_ (.A1(_04729_),
    .A2(\registers[14][21] ),
    .ZN(_04750_));
 OAI21_X1 _11198_ (.A(_04749_),
    .B1(_04750_),
    .B2(_04744_),
    .ZN(_00566_));
 NAND2_X1 _11199_ (.A1(_01205_),
    .A2(_04737_),
    .ZN(_04751_));
 CLKBUF_X3 _11200_ (.A(_04498_),
    .Z(_04752_));
 NAND2_X1 _11201_ (.A1(_04752_),
    .A2(\registers[14][22] ),
    .ZN(_04753_));
 OAI21_X1 _11202_ (.A(_04751_),
    .B1(_04753_),
    .B2(_04744_),
    .ZN(_00567_));
 NAND2_X1 _11203_ (.A1(_01209_),
    .A2(_04737_),
    .ZN(_04754_));
 NAND2_X1 _11204_ (.A1(_04752_),
    .A2(\registers[14][23] ),
    .ZN(_04755_));
 OAI21_X1 _11205_ (.A(_04754_),
    .B1(_04755_),
    .B2(_04744_),
    .ZN(_00568_));
 NAND2_X1 _11206_ (.A1(_01213_),
    .A2(_04737_),
    .ZN(_04756_));
 NAND2_X1 _11207_ (.A1(_04752_),
    .A2(\registers[14][24] ),
    .ZN(_04757_));
 OAI21_X1 _11208_ (.A(_04756_),
    .B1(_04757_),
    .B2(_04744_),
    .ZN(_00569_));
 NAND2_X1 _11209_ (.A1(_01217_),
    .A2(_04737_),
    .ZN(_04758_));
 NAND2_X1 _11210_ (.A1(_04752_),
    .A2(\registers[14][25] ),
    .ZN(_04759_));
 OAI21_X1 _11211_ (.A(_04758_),
    .B1(_04759_),
    .B2(_04744_),
    .ZN(_00570_));
 CLKBUF_X3 _11212_ (.A(_04717_),
    .Z(_04760_));
 NAND2_X1 _11213_ (.A1(_01221_),
    .A2(_04760_),
    .ZN(_04761_));
 NAND2_X1 _11214_ (.A1(_04752_),
    .A2(\registers[14][26] ),
    .ZN(_04762_));
 OAI21_X1 _11215_ (.A(_04761_),
    .B1(_04762_),
    .B2(_04744_),
    .ZN(_00571_));
 NAND2_X1 _11216_ (.A1(_01226_),
    .A2(_04760_),
    .ZN(_04763_));
 NAND2_X1 _11217_ (.A1(_04752_),
    .A2(\registers[14][27] ),
    .ZN(_04764_));
 OAI21_X1 _11218_ (.A(_04763_),
    .B1(_04764_),
    .B2(_04744_),
    .ZN(_00572_));
 NAND2_X1 _11219_ (.A1(_01230_),
    .A2(_04760_),
    .ZN(_04765_));
 NAND2_X1 _11220_ (.A1(_04752_),
    .A2(\registers[14][28] ),
    .ZN(_04766_));
 CLKBUF_X3 _11221_ (.A(_04717_),
    .Z(_04767_));
 OAI21_X1 _11222_ (.A(_04765_),
    .B1(_04766_),
    .B2(_04767_),
    .ZN(_00573_));
 NAND2_X1 _11223_ (.A1(_01235_),
    .A2(_04760_),
    .ZN(_04768_));
 NAND2_X1 _11224_ (.A1(_04752_),
    .A2(\registers[14][29] ),
    .ZN(_04769_));
 OAI21_X1 _11225_ (.A(_04768_),
    .B1(_04769_),
    .B2(_04767_),
    .ZN(_00574_));
 NAND2_X1 _11226_ (.A1(_01239_),
    .A2(_04760_),
    .ZN(_04770_));
 NAND2_X1 _11227_ (.A1(_04752_),
    .A2(\registers[14][2] ),
    .ZN(_04771_));
 OAI21_X1 _11228_ (.A(_04770_),
    .B1(_04771_),
    .B2(_04767_),
    .ZN(_00575_));
 NAND2_X1 _11229_ (.A1(_01244_),
    .A2(_04760_),
    .ZN(_04772_));
 NAND2_X1 _11230_ (.A1(_04752_),
    .A2(\registers[14][30] ),
    .ZN(_04773_));
 OAI21_X1 _11231_ (.A(_04772_),
    .B1(_04773_),
    .B2(_04767_),
    .ZN(_00576_));
 BUF_X4 _11232_ (.A(_01088_),
    .Z(_04774_));
 NAND2_X1 _11233_ (.A1(_04774_),
    .A2(_04760_),
    .ZN(_04775_));
 BUF_X4 _11234_ (.A(_04498_),
    .Z(_04776_));
 NAND2_X1 _11235_ (.A1(_04776_),
    .A2(\registers[14][31] ),
    .ZN(_04777_));
 OAI21_X1 _11236_ (.A(_04775_),
    .B1(_04777_),
    .B2(_04767_),
    .ZN(_00577_));
 BUF_X4 _11237_ (.A(_01108_),
    .Z(_04778_));
 NAND2_X1 _11238_ (.A1(_04778_),
    .A2(_04760_),
    .ZN(_04779_));
 NAND2_X1 _11239_ (.A1(_04776_),
    .A2(\registers[14][3] ),
    .ZN(_04780_));
 OAI21_X1 _11240_ (.A(_04779_),
    .B1(_04780_),
    .B2(_04767_),
    .ZN(_00578_));
 BUF_X4 _11241_ (.A(_01112_),
    .Z(_04781_));
 NAND2_X1 _11242_ (.A1(_04781_),
    .A2(_04760_),
    .ZN(_04782_));
 NAND2_X1 _11243_ (.A1(_04776_),
    .A2(\registers[14][4] ),
    .ZN(_04783_));
 OAI21_X1 _11244_ (.A(_04782_),
    .B1(_04783_),
    .B2(_04767_),
    .ZN(_00579_));
 BUF_X4 _11245_ (.A(_01116_),
    .Z(_04784_));
 NAND2_X1 _11246_ (.A1(_04784_),
    .A2(_04760_),
    .ZN(_04785_));
 NAND2_X1 _11247_ (.A1(_04776_),
    .A2(\registers[14][5] ),
    .ZN(_04786_));
 OAI21_X1 _11248_ (.A(_04785_),
    .B1(_04786_),
    .B2(_04767_),
    .ZN(_00580_));
 BUF_X4 _11249_ (.A(_01120_),
    .Z(_04787_));
 NAND2_X1 _11250_ (.A1(_04787_),
    .A2(_04717_),
    .ZN(_04788_));
 NAND2_X1 _11251_ (.A1(_04776_),
    .A2(\registers[14][6] ),
    .ZN(_04789_));
 OAI21_X1 _11252_ (.A(_04788_),
    .B1(_04789_),
    .B2(_04767_),
    .ZN(_00581_));
 BUF_X4 _11253_ (.A(_01124_),
    .Z(_04790_));
 NAND2_X1 _11254_ (.A1(_04790_),
    .A2(_04717_),
    .ZN(_04791_));
 NAND2_X1 _11255_ (.A1(_04776_),
    .A2(\registers[14][7] ),
    .ZN(_04792_));
 OAI21_X1 _11256_ (.A(_04791_),
    .B1(_04792_),
    .B2(_04767_),
    .ZN(_00582_));
 BUF_X4 _11257_ (.A(_01128_),
    .Z(_04793_));
 NAND2_X1 _11258_ (.A1(_04793_),
    .A2(_04717_),
    .ZN(_04794_));
 NAND2_X1 _11259_ (.A1(_04776_),
    .A2(\registers[14][8] ),
    .ZN(_04795_));
 OAI21_X1 _11260_ (.A(_04794_),
    .B1(_04795_),
    .B2(_04718_),
    .ZN(_00583_));
 BUF_X4 _11261_ (.A(_01132_),
    .Z(_04796_));
 NAND2_X1 _11262_ (.A1(_04796_),
    .A2(_04717_),
    .ZN(_04797_));
 NAND2_X1 _11263_ (.A1(_04776_),
    .A2(\registers[14][9] ),
    .ZN(_04798_));
 OAI21_X1 _11264_ (.A(_04797_),
    .B1(_04798_),
    .B2(_04718_),
    .ZN(_00584_));
 BUF_X4 _11265_ (.A(_01136_),
    .Z(_04799_));
 NOR2_X1 _11266_ (.A1(_01340_),
    .A2(_04597_),
    .ZN(_04800_));
 CLKBUF_X3 _11267_ (.A(_04800_),
    .Z(_04801_));
 CLKBUF_X3 _11268_ (.A(_04801_),
    .Z(_04802_));
 NAND2_X1 _11269_ (.A1(_04799_),
    .A2(_04802_),
    .ZN(_04803_));
 NAND2_X1 _11270_ (.A1(_04776_),
    .A2(\registers[15][0] ),
    .ZN(_04804_));
 CLKBUF_X3 _11271_ (.A(_04801_),
    .Z(_04805_));
 OAI21_X1 _11272_ (.A(_04803_),
    .B1(_04804_),
    .B2(_04805_),
    .ZN(_00585_));
 BUF_X4 _11273_ (.A(_01148_),
    .Z(_04806_));
 NAND2_X1 _11274_ (.A1(_04806_),
    .A2(_04802_),
    .ZN(_04807_));
 NAND2_X1 _11275_ (.A1(_04776_),
    .A2(\registers[15][10] ),
    .ZN(_04808_));
 OAI21_X1 _11276_ (.A(_04807_),
    .B1(_04808_),
    .B2(_04805_),
    .ZN(_00586_));
 BUF_X4 _11277_ (.A(_01152_),
    .Z(_04809_));
 NAND2_X1 _11278_ (.A1(_04809_),
    .A2(_04802_),
    .ZN(_04810_));
 CLKBUF_X3 _11279_ (.A(_04498_),
    .Z(_04811_));
 NAND2_X1 _11280_ (.A1(_04811_),
    .A2(\registers[15][11] ),
    .ZN(_04812_));
 OAI21_X1 _11281_ (.A(_04810_),
    .B1(_04812_),
    .B2(_04805_),
    .ZN(_00587_));
 BUF_X4 _11282_ (.A(_01157_),
    .Z(_04813_));
 NAND2_X1 _11283_ (.A1(_04813_),
    .A2(_04802_),
    .ZN(_04814_));
 NAND2_X1 _11284_ (.A1(_04811_),
    .A2(\registers[15][12] ),
    .ZN(_04815_));
 OAI21_X1 _11285_ (.A(_04814_),
    .B1(_04815_),
    .B2(_04805_),
    .ZN(_00588_));
 BUF_X4 _11286_ (.A(_01161_),
    .Z(_04816_));
 NAND2_X1 _11287_ (.A1(_04816_),
    .A2(_04802_),
    .ZN(_04817_));
 NAND2_X1 _11288_ (.A1(_04811_),
    .A2(\registers[15][13] ),
    .ZN(_04818_));
 OAI21_X1 _11289_ (.A(_04817_),
    .B1(_04818_),
    .B2(_04805_),
    .ZN(_00589_));
 BUF_X4 _11290_ (.A(_01165_),
    .Z(_04819_));
 NAND2_X1 _11291_ (.A1(_04819_),
    .A2(_04802_),
    .ZN(_04820_));
 NAND2_X1 _11292_ (.A1(_04811_),
    .A2(\registers[15][14] ),
    .ZN(_04821_));
 OAI21_X1 _11293_ (.A(_04820_),
    .B1(_04821_),
    .B2(_04805_),
    .ZN(_00590_));
 BUF_X4 _11294_ (.A(_01169_),
    .Z(_04822_));
 NAND2_X1 _11295_ (.A1(_04822_),
    .A2(_04802_),
    .ZN(_04823_));
 NAND2_X1 _11296_ (.A1(_04811_),
    .A2(\registers[15][15] ),
    .ZN(_04824_));
 OAI21_X1 _11297_ (.A(_04823_),
    .B1(_04824_),
    .B2(_04805_),
    .ZN(_00591_));
 BUF_X4 _11298_ (.A(_01173_),
    .Z(_04825_));
 NAND2_X1 _11299_ (.A1(_04825_),
    .A2(_04802_),
    .ZN(_04826_));
 NAND2_X1 _11300_ (.A1(_04811_),
    .A2(\registers[15][16] ),
    .ZN(_04827_));
 OAI21_X1 _11301_ (.A(_04826_),
    .B1(_04827_),
    .B2(_04805_),
    .ZN(_00592_));
 BUF_X4 _11302_ (.A(_01177_),
    .Z(_04828_));
 CLKBUF_X3 _11303_ (.A(_04801_),
    .Z(_04829_));
 NAND2_X1 _11304_ (.A1(_04828_),
    .A2(_04829_),
    .ZN(_04830_));
 NAND2_X1 _11305_ (.A1(_04811_),
    .A2(\registers[15][17] ),
    .ZN(_04831_));
 OAI21_X1 _11306_ (.A(_04830_),
    .B1(_04831_),
    .B2(_04805_),
    .ZN(_00593_));
 BUF_X4 _11307_ (.A(_01182_),
    .Z(_04832_));
 NAND2_X1 _11308_ (.A1(_04832_),
    .A2(_04829_),
    .ZN(_04833_));
 NAND2_X1 _11309_ (.A1(_04811_),
    .A2(\registers[15][18] ),
    .ZN(_04834_));
 OAI21_X1 _11310_ (.A(_04833_),
    .B1(_04834_),
    .B2(_04805_),
    .ZN(_00594_));
 BUF_X4 _11311_ (.A(_01186_),
    .Z(_04835_));
 NAND2_X1 _11312_ (.A1(_04835_),
    .A2(_04829_),
    .ZN(_04836_));
 NAND2_X1 _11313_ (.A1(_04811_),
    .A2(\registers[15][19] ),
    .ZN(_04837_));
 CLKBUF_X3 _11314_ (.A(_04801_),
    .Z(_04838_));
 OAI21_X1 _11315_ (.A(_04836_),
    .B1(_04837_),
    .B2(_04838_),
    .ZN(_00595_));
 BUF_X4 _11316_ (.A(_01191_),
    .Z(_04839_));
 NAND2_X1 _11317_ (.A1(_04839_),
    .A2(_04829_),
    .ZN(_04840_));
 NAND2_X1 _11318_ (.A1(_04811_),
    .A2(\registers[15][1] ),
    .ZN(_04841_));
 OAI21_X1 _11319_ (.A(_04840_),
    .B1(_04841_),
    .B2(_04838_),
    .ZN(_00596_));
 BUF_X4 _11320_ (.A(_01195_),
    .Z(_04842_));
 NAND2_X1 _11321_ (.A1(_04842_),
    .A2(_04829_),
    .ZN(_04843_));
 BUF_X4 _11322_ (.A(_01103_),
    .Z(_04844_));
 CLKBUF_X3 _11323_ (.A(_04844_),
    .Z(_04845_));
 NAND2_X1 _11324_ (.A1(_04845_),
    .A2(\registers[15][20] ),
    .ZN(_04846_));
 OAI21_X1 _11325_ (.A(_04843_),
    .B1(_04846_),
    .B2(_04838_),
    .ZN(_00597_));
 BUF_X4 _11326_ (.A(_01200_),
    .Z(_04847_));
 NAND2_X1 _11327_ (.A1(_04847_),
    .A2(_04829_),
    .ZN(_04848_));
 NAND2_X1 _11328_ (.A1(_04845_),
    .A2(\registers[15][21] ),
    .ZN(_04849_));
 OAI21_X1 _11329_ (.A(_04848_),
    .B1(_04849_),
    .B2(_04838_),
    .ZN(_00598_));
 BUF_X4 _11330_ (.A(_01204_),
    .Z(_04850_));
 NAND2_X1 _11331_ (.A1(_04850_),
    .A2(_04829_),
    .ZN(_04851_));
 NAND2_X1 _11332_ (.A1(_04845_),
    .A2(\registers[15][22] ),
    .ZN(_04852_));
 OAI21_X1 _11333_ (.A(_04851_),
    .B1(_04852_),
    .B2(_04838_),
    .ZN(_00599_));
 BUF_X4 _11334_ (.A(_01208_),
    .Z(_04853_));
 NAND2_X1 _11335_ (.A1(_04853_),
    .A2(_04829_),
    .ZN(_04854_));
 NAND2_X1 _11336_ (.A1(_04845_),
    .A2(\registers[15][23] ),
    .ZN(_04855_));
 OAI21_X1 _11337_ (.A(_04854_),
    .B1(_04855_),
    .B2(_04838_),
    .ZN(_00600_));
 BUF_X4 _11338_ (.A(_01212_),
    .Z(_04856_));
 NAND2_X1 _11339_ (.A1(_04856_),
    .A2(_04829_),
    .ZN(_04857_));
 NAND2_X1 _11340_ (.A1(_04845_),
    .A2(\registers[15][24] ),
    .ZN(_04858_));
 OAI21_X1 _11341_ (.A(_04857_),
    .B1(_04858_),
    .B2(_04838_),
    .ZN(_00601_));
 BUF_X4 _11342_ (.A(_01216_),
    .Z(_04859_));
 NAND2_X1 _11343_ (.A1(_04859_),
    .A2(_04829_),
    .ZN(_04860_));
 NAND2_X1 _11344_ (.A1(_04845_),
    .A2(\registers[15][25] ),
    .ZN(_04861_));
 OAI21_X1 _11345_ (.A(_04860_),
    .B1(_04861_),
    .B2(_04838_),
    .ZN(_00602_));
 BUF_X4 _11346_ (.A(_01220_),
    .Z(_04862_));
 CLKBUF_X3 _11347_ (.A(_04801_),
    .Z(_04863_));
 NAND2_X1 _11348_ (.A1(_04862_),
    .A2(_04863_),
    .ZN(_04864_));
 NAND2_X1 _11349_ (.A1(_04845_),
    .A2(\registers[15][26] ),
    .ZN(_04865_));
 OAI21_X1 _11350_ (.A(_04864_),
    .B1(_04865_),
    .B2(_04838_),
    .ZN(_00603_));
 BUF_X4 _11351_ (.A(_01225_),
    .Z(_04866_));
 NAND2_X1 _11352_ (.A1(_04866_),
    .A2(_04863_),
    .ZN(_04867_));
 NAND2_X1 _11353_ (.A1(_04845_),
    .A2(\registers[15][27] ),
    .ZN(_04868_));
 OAI21_X1 _11354_ (.A(_04867_),
    .B1(_04868_),
    .B2(_04838_),
    .ZN(_00604_));
 BUF_X4 _11355_ (.A(_01229_),
    .Z(_04869_));
 NAND2_X1 _11356_ (.A1(_04869_),
    .A2(_04863_),
    .ZN(_04870_));
 NAND2_X1 _11357_ (.A1(_04845_),
    .A2(\registers[15][28] ),
    .ZN(_04871_));
 CLKBUF_X3 _11358_ (.A(_04801_),
    .Z(_04872_));
 OAI21_X1 _11359_ (.A(_04870_),
    .B1(_04871_),
    .B2(_04872_),
    .ZN(_00605_));
 BUF_X4 _11360_ (.A(_01234_),
    .Z(_04873_));
 NAND2_X1 _11361_ (.A1(_04873_),
    .A2(_04863_),
    .ZN(_04874_));
 NAND2_X1 _11362_ (.A1(_04845_),
    .A2(\registers[15][29] ),
    .ZN(_04875_));
 OAI21_X1 _11363_ (.A(_04874_),
    .B1(_04875_),
    .B2(_04872_),
    .ZN(_00606_));
 BUF_X4 _11364_ (.A(_01238_),
    .Z(_04876_));
 NAND2_X1 _11365_ (.A1(_04876_),
    .A2(_04863_),
    .ZN(_04877_));
 CLKBUF_X3 _11366_ (.A(_04844_),
    .Z(_04878_));
 NAND2_X1 _11367_ (.A1(_04878_),
    .A2(\registers[15][2] ),
    .ZN(_04879_));
 OAI21_X1 _11368_ (.A(_04877_),
    .B1(_04879_),
    .B2(_04872_),
    .ZN(_00607_));
 BUF_X4 _11369_ (.A(_01243_),
    .Z(_04880_));
 NAND2_X1 _11370_ (.A1(_04880_),
    .A2(_04863_),
    .ZN(_04881_));
 NAND2_X1 _11371_ (.A1(_04878_),
    .A2(\registers[15][30] ),
    .ZN(_04882_));
 OAI21_X1 _11372_ (.A(_04881_),
    .B1(_04882_),
    .B2(_04872_),
    .ZN(_00608_));
 NAND2_X1 _11373_ (.A1(_04774_),
    .A2(_04863_),
    .ZN(_04883_));
 NAND2_X1 _11374_ (.A1(_04878_),
    .A2(\registers[15][31] ),
    .ZN(_04884_));
 OAI21_X1 _11375_ (.A(_04883_),
    .B1(_04884_),
    .B2(_04872_),
    .ZN(_00609_));
 NAND2_X1 _11376_ (.A1(_04778_),
    .A2(_04863_),
    .ZN(_04885_));
 NAND2_X1 _11377_ (.A1(_04878_),
    .A2(\registers[15][3] ),
    .ZN(_04886_));
 OAI21_X1 _11378_ (.A(_04885_),
    .B1(_04886_),
    .B2(_04872_),
    .ZN(_00610_));
 NAND2_X1 _11379_ (.A1(_04781_),
    .A2(_04863_),
    .ZN(_04887_));
 NAND2_X1 _11380_ (.A1(_04878_),
    .A2(\registers[15][4] ),
    .ZN(_04888_));
 OAI21_X1 _11381_ (.A(_04887_),
    .B1(_04888_),
    .B2(_04872_),
    .ZN(_00611_));
 NAND2_X1 _11382_ (.A1(_04784_),
    .A2(_04863_),
    .ZN(_04889_));
 NAND2_X1 _11383_ (.A1(_04878_),
    .A2(\registers[15][5] ),
    .ZN(_04890_));
 OAI21_X1 _11384_ (.A(_04889_),
    .B1(_04890_),
    .B2(_04872_),
    .ZN(_00612_));
 NAND2_X1 _11385_ (.A1(_04787_),
    .A2(_04801_),
    .ZN(_04891_));
 NAND2_X1 _11386_ (.A1(_04878_),
    .A2(\registers[15][6] ),
    .ZN(_04892_));
 OAI21_X1 _11387_ (.A(_04891_),
    .B1(_04892_),
    .B2(_04872_),
    .ZN(_00613_));
 NAND2_X1 _11388_ (.A1(_04790_),
    .A2(_04801_),
    .ZN(_04893_));
 NAND2_X1 _11389_ (.A1(_04878_),
    .A2(\registers[15][7] ),
    .ZN(_04894_));
 OAI21_X1 _11390_ (.A(_04893_),
    .B1(_04894_),
    .B2(_04872_),
    .ZN(_00614_));
 NAND2_X1 _11391_ (.A1(_04793_),
    .A2(_04801_),
    .ZN(_04895_));
 NAND2_X1 _11392_ (.A1(_04878_),
    .A2(\registers[15][8] ),
    .ZN(_04896_));
 OAI21_X1 _11393_ (.A(_04895_),
    .B1(_04896_),
    .B2(_04802_),
    .ZN(_00615_));
 NAND2_X1 _11394_ (.A1(_04796_),
    .A2(_04801_),
    .ZN(_04897_));
 NAND2_X1 _11395_ (.A1(_04878_),
    .A2(\registers[15][9] ),
    .ZN(_04898_));
 OAI21_X1 _11396_ (.A(_04897_),
    .B1(_04898_),
    .B2(_04802_),
    .ZN(_00616_));
 NOR3_X1 _11397_ (.A1(_01090_),
    .A2(_01738_),
    .A3(_01092_),
    .ZN(_04899_));
 NAND2_X1 _11398_ (.A1(_01497_),
    .A2(_04899_),
    .ZN(_04900_));
 CLKBUF_X3 _11399_ (.A(_04900_),
    .Z(_04901_));
 CLKBUF_X3 _11400_ (.A(_04901_),
    .Z(_04902_));
 NAND3_X1 _11401_ (.A1(_04638_),
    .A2(\registers[16][0] ),
    .A3(_04902_),
    .ZN(_04903_));
 CLKBUF_X3 _11402_ (.A(_04901_),
    .Z(_04904_));
 OAI21_X1 _11403_ (.A(_04903_),
    .B1(_04904_),
    .B2(_01424_),
    .ZN(_00617_));
 NAND3_X1 _11404_ (.A1(_04638_),
    .A2(\registers[16][10] ),
    .A3(_04902_),
    .ZN(_04905_));
 OAI21_X1 _11405_ (.A(_04905_),
    .B1(_04904_),
    .B2(_01426_),
    .ZN(_00618_));
 NAND3_X1 _11406_ (.A1(_04638_),
    .A2(\registers[16][11] ),
    .A3(_04902_),
    .ZN(_04906_));
 OAI21_X1 _11407_ (.A(_04906_),
    .B1(_04904_),
    .B2(_01428_),
    .ZN(_00619_));
 NAND3_X1 _11408_ (.A1(_04638_),
    .A2(\registers[16][12] ),
    .A3(_04902_),
    .ZN(_04907_));
 OAI21_X1 _11409_ (.A(_04907_),
    .B1(_04904_),
    .B2(_01430_),
    .ZN(_00620_));
 NAND3_X1 _11410_ (.A1(_04638_),
    .A2(\registers[16][13] ),
    .A3(_04902_),
    .ZN(_04908_));
 OAI21_X1 _11411_ (.A(_04908_),
    .B1(_04904_),
    .B2(_01432_),
    .ZN(_00621_));
 NAND3_X1 _11412_ (.A1(_04638_),
    .A2(\registers[16][14] ),
    .A3(_04902_),
    .ZN(_04909_));
 OAI21_X1 _11413_ (.A(_04909_),
    .B1(_04904_),
    .B2(_01434_),
    .ZN(_00622_));
 NAND3_X1 _11414_ (.A1(_04638_),
    .A2(\registers[16][15] ),
    .A3(_04902_),
    .ZN(_04910_));
 OAI21_X1 _11415_ (.A(_04910_),
    .B1(_04904_),
    .B2(_01436_),
    .ZN(_00623_));
 NAND3_X1 _11416_ (.A1(_04638_),
    .A2(\registers[16][16] ),
    .A3(_04902_),
    .ZN(_04911_));
 OAI21_X1 _11417_ (.A(_04911_),
    .B1(_04904_),
    .B2(_01438_),
    .ZN(_00624_));
 CLKBUF_X3 _11418_ (.A(_04595_),
    .Z(_04912_));
 CLKBUF_X3 _11419_ (.A(_04901_),
    .Z(_04913_));
 NAND3_X1 _11420_ (.A1(_04912_),
    .A2(\registers[16][17] ),
    .A3(_04913_),
    .ZN(_04914_));
 OAI21_X1 _11421_ (.A(_04914_),
    .B1(_04904_),
    .B2(_01441_),
    .ZN(_00625_));
 NAND3_X1 _11422_ (.A1(_04912_),
    .A2(\registers[16][18] ),
    .A3(_04913_),
    .ZN(_04915_));
 OAI21_X1 _11423_ (.A(_04915_),
    .B1(_04904_),
    .B2(_01443_),
    .ZN(_00626_));
 NAND3_X1 _11424_ (.A1(_04912_),
    .A2(\registers[16][19] ),
    .A3(_04913_),
    .ZN(_04916_));
 CLKBUF_X3 _11425_ (.A(_04901_),
    .Z(_04917_));
 OAI21_X1 _11426_ (.A(_04916_),
    .B1(_04917_),
    .B2(_01447_),
    .ZN(_00627_));
 NAND3_X1 _11427_ (.A1(_04912_),
    .A2(\registers[16][1] ),
    .A3(_04913_),
    .ZN(_04918_));
 OAI21_X1 _11428_ (.A(_04918_),
    .B1(_04917_),
    .B2(_01449_),
    .ZN(_00628_));
 NAND3_X1 _11429_ (.A1(_04912_),
    .A2(\registers[16][20] ),
    .A3(_04913_),
    .ZN(_04919_));
 OAI21_X1 _11430_ (.A(_04919_),
    .B1(_04917_),
    .B2(_01451_),
    .ZN(_00629_));
 NAND3_X1 _11431_ (.A1(_04912_),
    .A2(\registers[16][21] ),
    .A3(_04913_),
    .ZN(_04920_));
 OAI21_X1 _11432_ (.A(_04920_),
    .B1(_04917_),
    .B2(_01453_),
    .ZN(_00630_));
 NAND3_X1 _11433_ (.A1(_04912_),
    .A2(\registers[16][22] ),
    .A3(_04913_),
    .ZN(_04921_));
 OAI21_X1 _11434_ (.A(_04921_),
    .B1(_04917_),
    .B2(_01455_),
    .ZN(_00631_));
 NAND3_X1 _11435_ (.A1(_04912_),
    .A2(\registers[16][23] ),
    .A3(_04913_),
    .ZN(_04922_));
 OAI21_X1 _11436_ (.A(_04922_),
    .B1(_04917_),
    .B2(_01457_),
    .ZN(_00632_));
 NAND3_X1 _11437_ (.A1(_04912_),
    .A2(\registers[16][24] ),
    .A3(_04913_),
    .ZN(_04923_));
 OAI21_X1 _11438_ (.A(_04923_),
    .B1(_04917_),
    .B2(_01459_),
    .ZN(_00633_));
 NAND3_X1 _11439_ (.A1(_04912_),
    .A2(\registers[16][25] ),
    .A3(_04913_),
    .ZN(_04924_));
 OAI21_X1 _11440_ (.A(_04924_),
    .B1(_04917_),
    .B2(_01461_),
    .ZN(_00634_));
 CLKBUF_X3 _11441_ (.A(_04595_),
    .Z(_04925_));
 CLKBUF_X3 _11442_ (.A(_04901_),
    .Z(_04926_));
 NAND3_X1 _11443_ (.A1(_04925_),
    .A2(\registers[16][26] ),
    .A3(_04926_),
    .ZN(_04927_));
 OAI21_X1 _11444_ (.A(_04927_),
    .B1(_04917_),
    .B2(_01464_),
    .ZN(_00635_));
 NAND3_X1 _11445_ (.A1(_04925_),
    .A2(\registers[16][27] ),
    .A3(_04926_),
    .ZN(_04928_));
 OAI21_X1 _11446_ (.A(_04928_),
    .B1(_04917_),
    .B2(_01466_),
    .ZN(_00636_));
 NAND3_X1 _11447_ (.A1(_04925_),
    .A2(\registers[16][28] ),
    .A3(_04926_),
    .ZN(_04929_));
 CLKBUF_X3 _11448_ (.A(_04901_),
    .Z(_04930_));
 OAI21_X1 _11449_ (.A(_04929_),
    .B1(_04930_),
    .B2(_01470_),
    .ZN(_00637_));
 NAND3_X1 _11450_ (.A1(_04925_),
    .A2(\registers[16][29] ),
    .A3(_04926_),
    .ZN(_04931_));
 OAI21_X1 _11451_ (.A(_04931_),
    .B1(_04930_),
    .B2(_01472_),
    .ZN(_00638_));
 NAND3_X1 _11452_ (.A1(_04925_),
    .A2(\registers[16][2] ),
    .A3(_04926_),
    .ZN(_04932_));
 OAI21_X1 _11453_ (.A(_04932_),
    .B1(_04930_),
    .B2(_01474_),
    .ZN(_00639_));
 NAND3_X1 _11454_ (.A1(_04925_),
    .A2(\registers[16][30] ),
    .A3(_04926_),
    .ZN(_04933_));
 OAI21_X1 _11455_ (.A(_04933_),
    .B1(_04930_),
    .B2(_01476_),
    .ZN(_00640_));
 NAND3_X1 _11456_ (.A1(_04925_),
    .A2(\registers[16][31] ),
    .A3(_04926_),
    .ZN(_04934_));
 OAI21_X1 _11457_ (.A(_04934_),
    .B1(_04930_),
    .B2(_01478_),
    .ZN(_00641_));
 NAND3_X1 _11458_ (.A1(_04925_),
    .A2(\registers[16][3] ),
    .A3(_04926_),
    .ZN(_04935_));
 OAI21_X1 _11459_ (.A(_04935_),
    .B1(_04930_),
    .B2(_01480_),
    .ZN(_00642_));
 NAND3_X1 _11460_ (.A1(_04925_),
    .A2(\registers[16][4] ),
    .A3(_04926_),
    .ZN(_04936_));
 OAI21_X1 _11461_ (.A(_04936_),
    .B1(_04930_),
    .B2(_01482_),
    .ZN(_00643_));
 NAND3_X1 _11462_ (.A1(_04925_),
    .A2(\registers[16][5] ),
    .A3(_04926_),
    .ZN(_04937_));
 OAI21_X1 _11463_ (.A(_04937_),
    .B1(_04930_),
    .B2(_01484_),
    .ZN(_00644_));
 BUF_X4 _11464_ (.A(_04595_),
    .Z(_04938_));
 NAND3_X1 _11465_ (.A1(_04938_),
    .A2(\registers[16][6] ),
    .A3(_04901_),
    .ZN(_04939_));
 OAI21_X1 _11466_ (.A(_04939_),
    .B1(_04930_),
    .B2(_01486_),
    .ZN(_00645_));
 NAND3_X1 _11467_ (.A1(_04938_),
    .A2(\registers[16][7] ),
    .A3(_04901_),
    .ZN(_04940_));
 OAI21_X1 _11468_ (.A(_04940_),
    .B1(_04930_),
    .B2(_01488_),
    .ZN(_00646_));
 NAND3_X1 _11469_ (.A1(_04938_),
    .A2(\registers[16][8] ),
    .A3(_04901_),
    .ZN(_04941_));
 OAI21_X1 _11470_ (.A(_04941_),
    .B1(_04902_),
    .B2(_01491_),
    .ZN(_00647_));
 NAND3_X1 _11471_ (.A1(_04938_),
    .A2(\registers[16][9] ),
    .A3(_04901_),
    .ZN(_04942_));
 OAI21_X1 _11472_ (.A(_04942_),
    .B1(_04902_),
    .B2(_01493_),
    .ZN(_00648_));
 NAND2_X1 _11473_ (.A1(_01542_),
    .A2(_04899_),
    .ZN(_04943_));
 CLKBUF_X3 _11474_ (.A(_04943_),
    .Z(_04944_));
 CLKBUF_X3 _11475_ (.A(_04944_),
    .Z(_04945_));
 NAND3_X1 _11476_ (.A1(_04938_),
    .A2(\registers[17][0] ),
    .A3(_04945_),
    .ZN(_04946_));
 CLKBUF_X3 _11477_ (.A(_04944_),
    .Z(_04947_));
 OAI21_X1 _11478_ (.A(_04946_),
    .B1(_04947_),
    .B2(_01424_),
    .ZN(_00649_));
 NAND3_X1 _11479_ (.A1(_04938_),
    .A2(\registers[17][10] ),
    .A3(_04945_),
    .ZN(_04948_));
 OAI21_X1 _11480_ (.A(_04948_),
    .B1(_04947_),
    .B2(_01426_),
    .ZN(_00650_));
 NAND3_X1 _11481_ (.A1(_04938_),
    .A2(\registers[17][11] ),
    .A3(_04945_),
    .ZN(_04949_));
 OAI21_X1 _11482_ (.A(_04949_),
    .B1(_04947_),
    .B2(_01428_),
    .ZN(_00651_));
 NAND3_X1 _11483_ (.A1(_04938_),
    .A2(\registers[17][12] ),
    .A3(_04945_),
    .ZN(_04950_));
 OAI21_X1 _11484_ (.A(_04950_),
    .B1(_04947_),
    .B2(_01430_),
    .ZN(_00652_));
 NAND3_X1 _11485_ (.A1(_04938_),
    .A2(\registers[17][13] ),
    .A3(_04945_),
    .ZN(_04951_));
 OAI21_X1 _11486_ (.A(_04951_),
    .B1(_04947_),
    .B2(_01432_),
    .ZN(_00653_));
 NAND3_X1 _11487_ (.A1(_04938_),
    .A2(\registers[17][14] ),
    .A3(_04945_),
    .ZN(_04952_));
 OAI21_X1 _11488_ (.A(_04952_),
    .B1(_04947_),
    .B2(_01434_),
    .ZN(_00654_));
 CLKBUF_X3 _11489_ (.A(_04595_),
    .Z(_04953_));
 NAND3_X1 _11490_ (.A1(_04953_),
    .A2(\registers[17][15] ),
    .A3(_04945_),
    .ZN(_04954_));
 OAI21_X1 _11491_ (.A(_04954_),
    .B1(_04947_),
    .B2(_01436_),
    .ZN(_00655_));
 NAND3_X1 _11492_ (.A1(_04953_),
    .A2(\registers[17][16] ),
    .A3(_04945_),
    .ZN(_04955_));
 OAI21_X1 _11493_ (.A(_04955_),
    .B1(_04947_),
    .B2(_01438_),
    .ZN(_00656_));
 CLKBUF_X3 _11494_ (.A(_04944_),
    .Z(_04956_));
 NAND3_X1 _11495_ (.A1(_04953_),
    .A2(\registers[17][17] ),
    .A3(_04956_),
    .ZN(_04957_));
 OAI21_X1 _11496_ (.A(_04957_),
    .B1(_04947_),
    .B2(_01441_),
    .ZN(_00657_));
 NAND3_X1 _11497_ (.A1(_04953_),
    .A2(\registers[17][18] ),
    .A3(_04956_),
    .ZN(_04958_));
 OAI21_X1 _11498_ (.A(_04958_),
    .B1(_04947_),
    .B2(_01443_),
    .ZN(_00658_));
 NAND3_X1 _11499_ (.A1(_04953_),
    .A2(\registers[17][19] ),
    .A3(_04956_),
    .ZN(_04959_));
 CLKBUF_X3 _11500_ (.A(_04944_),
    .Z(_04960_));
 OAI21_X1 _11501_ (.A(_04959_),
    .B1(_04960_),
    .B2(_01447_),
    .ZN(_00659_));
 NAND3_X1 _11502_ (.A1(_04953_),
    .A2(\registers[17][1] ),
    .A3(_04956_),
    .ZN(_04961_));
 OAI21_X1 _11503_ (.A(_04961_),
    .B1(_04960_),
    .B2(_01449_),
    .ZN(_00660_));
 NAND3_X1 _11504_ (.A1(_04953_),
    .A2(\registers[17][20] ),
    .A3(_04956_),
    .ZN(_04962_));
 OAI21_X1 _11505_ (.A(_04962_),
    .B1(_04960_),
    .B2(_01451_),
    .ZN(_00661_));
 NAND3_X1 _11506_ (.A1(_04953_),
    .A2(\registers[17][21] ),
    .A3(_04956_),
    .ZN(_04963_));
 OAI21_X1 _11507_ (.A(_04963_),
    .B1(_04960_),
    .B2(_01453_),
    .ZN(_00662_));
 NAND3_X1 _11508_ (.A1(_04953_),
    .A2(\registers[17][22] ),
    .A3(_04956_),
    .ZN(_04964_));
 OAI21_X1 _11509_ (.A(_04964_),
    .B1(_04960_),
    .B2(_01455_),
    .ZN(_00663_));
 NAND3_X1 _11510_ (.A1(_04953_),
    .A2(\registers[17][23] ),
    .A3(_04956_),
    .ZN(_04965_));
 OAI21_X1 _11511_ (.A(_04965_),
    .B1(_04960_),
    .B2(_01457_),
    .ZN(_00664_));
 CLKBUF_X3 _11512_ (.A(_04595_),
    .Z(_04966_));
 NAND3_X1 _11513_ (.A1(_04966_),
    .A2(\registers[17][24] ),
    .A3(_04956_),
    .ZN(_04967_));
 OAI21_X1 _11514_ (.A(_04967_),
    .B1(_04960_),
    .B2(_01459_),
    .ZN(_00665_));
 NAND3_X1 _11515_ (.A1(_04966_),
    .A2(\registers[17][25] ),
    .A3(_04956_),
    .ZN(_04968_));
 OAI21_X1 _11516_ (.A(_04968_),
    .B1(_04960_),
    .B2(_01461_),
    .ZN(_00666_));
 CLKBUF_X3 _11517_ (.A(_04944_),
    .Z(_04969_));
 NAND3_X1 _11518_ (.A1(_04966_),
    .A2(\registers[17][26] ),
    .A3(_04969_),
    .ZN(_04970_));
 OAI21_X1 _11519_ (.A(_04970_),
    .B1(_04960_),
    .B2(_01464_),
    .ZN(_00667_));
 NAND3_X1 _11520_ (.A1(_04966_),
    .A2(\registers[17][27] ),
    .A3(_04969_),
    .ZN(_04971_));
 OAI21_X1 _11521_ (.A(_04971_),
    .B1(_04960_),
    .B2(_01466_),
    .ZN(_00668_));
 NAND3_X1 _11522_ (.A1(_04966_),
    .A2(\registers[17][28] ),
    .A3(_04969_),
    .ZN(_04972_));
 CLKBUF_X3 _11523_ (.A(_04944_),
    .Z(_04973_));
 OAI21_X1 _11524_ (.A(_04972_),
    .B1(_04973_),
    .B2(_01470_),
    .ZN(_00669_));
 NAND3_X1 _11525_ (.A1(_04966_),
    .A2(\registers[17][29] ),
    .A3(_04969_),
    .ZN(_04974_));
 OAI21_X1 _11526_ (.A(_04974_),
    .B1(_04973_),
    .B2(_01472_),
    .ZN(_00670_));
 NAND3_X1 _11527_ (.A1(_04966_),
    .A2(\registers[17][2] ),
    .A3(_04969_),
    .ZN(_04975_));
 OAI21_X1 _11528_ (.A(_04975_),
    .B1(_04973_),
    .B2(_01474_),
    .ZN(_00671_));
 NAND3_X1 _11529_ (.A1(_04966_),
    .A2(\registers[17][30] ),
    .A3(_04969_),
    .ZN(_04976_));
 OAI21_X1 _11530_ (.A(_04976_),
    .B1(_04973_),
    .B2(_01476_),
    .ZN(_00672_));
 NAND3_X1 _11531_ (.A1(_04966_),
    .A2(\registers[17][31] ),
    .A3(_04969_),
    .ZN(_04977_));
 OAI21_X1 _11532_ (.A(_04977_),
    .B1(_04973_),
    .B2(_01478_),
    .ZN(_00673_));
 NAND3_X1 _11533_ (.A1(_04966_),
    .A2(\registers[17][3] ),
    .A3(_04969_),
    .ZN(_04978_));
 OAI21_X1 _11534_ (.A(_04978_),
    .B1(_04973_),
    .B2(_01480_),
    .ZN(_00674_));
 BUF_X4 _11535_ (.A(_04595_),
    .Z(_04979_));
 NAND3_X1 _11536_ (.A1(_04979_),
    .A2(\registers[17][4] ),
    .A3(_04969_),
    .ZN(_04980_));
 OAI21_X1 _11537_ (.A(_04980_),
    .B1(_04973_),
    .B2(_01482_),
    .ZN(_00675_));
 NAND3_X1 _11538_ (.A1(_04979_),
    .A2(\registers[17][5] ),
    .A3(_04969_),
    .ZN(_04981_));
 OAI21_X1 _11539_ (.A(_04981_),
    .B1(_04973_),
    .B2(_01484_),
    .ZN(_00676_));
 NAND3_X1 _11540_ (.A1(_04979_),
    .A2(\registers[17][6] ),
    .A3(_04944_),
    .ZN(_04982_));
 OAI21_X1 _11541_ (.A(_04982_),
    .B1(_04973_),
    .B2(_01486_),
    .ZN(_00677_));
 NAND3_X1 _11542_ (.A1(_04979_),
    .A2(\registers[17][7] ),
    .A3(_04944_),
    .ZN(_04983_));
 OAI21_X1 _11543_ (.A(_04983_),
    .B1(_04973_),
    .B2(_01488_),
    .ZN(_00678_));
 NAND3_X1 _11544_ (.A1(_04979_),
    .A2(\registers[17][8] ),
    .A3(_04944_),
    .ZN(_04984_));
 OAI21_X1 _11545_ (.A(_04984_),
    .B1(_04945_),
    .B2(_01491_),
    .ZN(_00679_));
 NAND3_X1 _11546_ (.A1(_04979_),
    .A2(\registers[17][9] ),
    .A3(_04944_),
    .ZN(_04985_));
 OAI21_X1 _11547_ (.A(_04985_),
    .B1(_04945_),
    .B2(_01493_),
    .ZN(_00680_));
 NOR4_X4 _11548_ (.A1(_01090_),
    .A2(_01738_),
    .A3(_01092_),
    .A4(_01141_),
    .ZN(_04986_));
 BUF_X4 _11549_ (.A(_04986_),
    .Z(_04987_));
 BUF_X4 _11550_ (.A(_04987_),
    .Z(_04988_));
 NAND2_X1 _11551_ (.A1(_04799_),
    .A2(_04988_),
    .ZN(_04989_));
 CLKBUF_X3 _11552_ (.A(_04844_),
    .Z(_04990_));
 NAND2_X1 _11553_ (.A1(_04990_),
    .A2(\registers[18][0] ),
    .ZN(_04991_));
 CLKBUF_X3 _11554_ (.A(_04987_),
    .Z(_04992_));
 OAI21_X1 _11555_ (.A(_04989_),
    .B1(_04991_),
    .B2(_04992_),
    .ZN(_00681_));
 NAND2_X1 _11556_ (.A1(_04806_),
    .A2(_04988_),
    .ZN(_04993_));
 NAND2_X1 _11557_ (.A1(_04990_),
    .A2(\registers[18][10] ),
    .ZN(_04994_));
 OAI21_X1 _11558_ (.A(_04993_),
    .B1(_04994_),
    .B2(_04992_),
    .ZN(_00682_));
 NAND2_X1 _11559_ (.A1(_04809_),
    .A2(_04988_),
    .ZN(_04995_));
 NAND2_X1 _11560_ (.A1(_04990_),
    .A2(\registers[18][11] ),
    .ZN(_04996_));
 OAI21_X1 _11561_ (.A(_04995_),
    .B1(_04996_),
    .B2(_04992_),
    .ZN(_00683_));
 NAND2_X1 _11562_ (.A1(_04813_),
    .A2(_04988_),
    .ZN(_04997_));
 NAND2_X1 _11563_ (.A1(_04990_),
    .A2(\registers[18][12] ),
    .ZN(_04998_));
 OAI21_X1 _11564_ (.A(_04997_),
    .B1(_04998_),
    .B2(_04992_),
    .ZN(_00684_));
 NAND2_X1 _11565_ (.A1(_04816_),
    .A2(_04988_),
    .ZN(_04999_));
 NAND2_X1 _11566_ (.A1(_04990_),
    .A2(\registers[18][13] ),
    .ZN(_05000_));
 OAI21_X1 _11567_ (.A(_04999_),
    .B1(_05000_),
    .B2(_04992_),
    .ZN(_00685_));
 NAND2_X1 _11568_ (.A1(_04819_),
    .A2(_04988_),
    .ZN(_05001_));
 NAND2_X1 _11569_ (.A1(_04990_),
    .A2(\registers[18][14] ),
    .ZN(_05002_));
 OAI21_X1 _11570_ (.A(_05001_),
    .B1(_05002_),
    .B2(_04992_),
    .ZN(_00686_));
 NAND2_X1 _11571_ (.A1(_04822_),
    .A2(_04988_),
    .ZN(_05003_));
 NAND2_X1 _11572_ (.A1(_04990_),
    .A2(\registers[18][15] ),
    .ZN(_05004_));
 OAI21_X1 _11573_ (.A(_05003_),
    .B1(_05004_),
    .B2(_04992_),
    .ZN(_00687_));
 NAND2_X1 _11574_ (.A1(_04825_),
    .A2(_04988_),
    .ZN(_05005_));
 NAND2_X1 _11575_ (.A1(_04990_),
    .A2(\registers[18][16] ),
    .ZN(_05006_));
 OAI21_X1 _11576_ (.A(_05005_),
    .B1(_05006_),
    .B2(_04992_),
    .ZN(_00688_));
 BUF_X4 _11577_ (.A(_04987_),
    .Z(_05007_));
 NAND2_X1 _11578_ (.A1(_04828_),
    .A2(_05007_),
    .ZN(_05008_));
 NAND2_X1 _11579_ (.A1(_04990_),
    .A2(\registers[18][17] ),
    .ZN(_05009_));
 OAI21_X1 _11580_ (.A(_05008_),
    .B1(_05009_),
    .B2(_04992_),
    .ZN(_00689_));
 NAND2_X1 _11581_ (.A1(_04832_),
    .A2(_05007_),
    .ZN(_05010_));
 NAND2_X1 _11582_ (.A1(_04990_),
    .A2(\registers[18][18] ),
    .ZN(_05011_));
 OAI21_X1 _11583_ (.A(_05010_),
    .B1(_05011_),
    .B2(_04992_),
    .ZN(_00690_));
 NAND2_X1 _11584_ (.A1(_04835_),
    .A2(_05007_),
    .ZN(_05012_));
 CLKBUF_X3 _11585_ (.A(_04844_),
    .Z(_05013_));
 NAND2_X1 _11586_ (.A1(_05013_),
    .A2(\registers[18][19] ),
    .ZN(_05014_));
 CLKBUF_X3 _11587_ (.A(_04987_),
    .Z(_05015_));
 OAI21_X1 _11588_ (.A(_05012_),
    .B1(_05014_),
    .B2(_05015_),
    .ZN(_00691_));
 NAND2_X1 _11589_ (.A1(_04839_),
    .A2(_05007_),
    .ZN(_05016_));
 NAND2_X1 _11590_ (.A1(_05013_),
    .A2(\registers[18][1] ),
    .ZN(_05017_));
 OAI21_X1 _11591_ (.A(_05016_),
    .B1(_05017_),
    .B2(_05015_),
    .ZN(_00692_));
 NAND2_X1 _11592_ (.A1(_04842_),
    .A2(_05007_),
    .ZN(_05018_));
 NAND2_X1 _11593_ (.A1(_05013_),
    .A2(\registers[18][20] ),
    .ZN(_05019_));
 OAI21_X1 _11594_ (.A(_05018_),
    .B1(_05019_),
    .B2(_05015_),
    .ZN(_00693_));
 NAND2_X1 _11595_ (.A1(_04847_),
    .A2(_05007_),
    .ZN(_05020_));
 NAND2_X1 _11596_ (.A1(_05013_),
    .A2(\registers[18][21] ),
    .ZN(_05021_));
 OAI21_X1 _11597_ (.A(_05020_),
    .B1(_05021_),
    .B2(_05015_),
    .ZN(_00694_));
 NAND2_X1 _11598_ (.A1(_04850_),
    .A2(_05007_),
    .ZN(_05022_));
 NAND2_X1 _11599_ (.A1(_05013_),
    .A2(\registers[18][22] ),
    .ZN(_05023_));
 OAI21_X1 _11600_ (.A(_05022_),
    .B1(_05023_),
    .B2(_05015_),
    .ZN(_00695_));
 NAND2_X1 _11601_ (.A1(_04853_),
    .A2(_05007_),
    .ZN(_05024_));
 NAND2_X1 _11602_ (.A1(_05013_),
    .A2(\registers[18][23] ),
    .ZN(_05025_));
 OAI21_X1 _11603_ (.A(_05024_),
    .B1(_05025_),
    .B2(_05015_),
    .ZN(_00696_));
 NAND2_X1 _11604_ (.A1(_04856_),
    .A2(_05007_),
    .ZN(_05026_));
 NAND2_X1 _11605_ (.A1(_05013_),
    .A2(\registers[18][24] ),
    .ZN(_05027_));
 OAI21_X1 _11606_ (.A(_05026_),
    .B1(_05027_),
    .B2(_05015_),
    .ZN(_00697_));
 NAND2_X1 _11607_ (.A1(_04859_),
    .A2(_05007_),
    .ZN(_05028_));
 NAND2_X1 _11608_ (.A1(_05013_),
    .A2(\registers[18][25] ),
    .ZN(_05029_));
 OAI21_X1 _11609_ (.A(_05028_),
    .B1(_05029_),
    .B2(_05015_),
    .ZN(_00698_));
 BUF_X4 _11610_ (.A(_04987_),
    .Z(_05030_));
 NAND2_X1 _11611_ (.A1(_04862_),
    .A2(_05030_),
    .ZN(_05031_));
 NAND2_X1 _11612_ (.A1(_05013_),
    .A2(\registers[18][26] ),
    .ZN(_05032_));
 OAI21_X1 _11613_ (.A(_05031_),
    .B1(_05032_),
    .B2(_05015_),
    .ZN(_00699_));
 NAND2_X1 _11614_ (.A1(_04866_),
    .A2(_05030_),
    .ZN(_05033_));
 NAND2_X1 _11615_ (.A1(_05013_),
    .A2(\registers[18][27] ),
    .ZN(_05034_));
 OAI21_X1 _11616_ (.A(_05033_),
    .B1(_05034_),
    .B2(_05015_),
    .ZN(_00700_));
 NAND2_X1 _11617_ (.A1(_04869_),
    .A2(_05030_),
    .ZN(_05035_));
 CLKBUF_X3 _11618_ (.A(_04844_),
    .Z(_05036_));
 NAND2_X1 _11619_ (.A1(_05036_),
    .A2(\registers[18][28] ),
    .ZN(_05037_));
 CLKBUF_X3 _11620_ (.A(_04987_),
    .Z(_05038_));
 OAI21_X1 _11621_ (.A(_05035_),
    .B1(_05037_),
    .B2(_05038_),
    .ZN(_00701_));
 NAND2_X1 _11622_ (.A1(_04873_),
    .A2(_05030_),
    .ZN(_05039_));
 NAND2_X1 _11623_ (.A1(_05036_),
    .A2(\registers[18][29] ),
    .ZN(_05040_));
 OAI21_X1 _11624_ (.A(_05039_),
    .B1(_05040_),
    .B2(_05038_),
    .ZN(_00702_));
 NAND2_X1 _11625_ (.A1(_04876_),
    .A2(_05030_),
    .ZN(_05041_));
 NAND2_X1 _11626_ (.A1(_05036_),
    .A2(\registers[18][2] ),
    .ZN(_05042_));
 OAI21_X1 _11627_ (.A(_05041_),
    .B1(_05042_),
    .B2(_05038_),
    .ZN(_00703_));
 NAND2_X1 _11628_ (.A1(_04880_),
    .A2(_05030_),
    .ZN(_05043_));
 NAND2_X1 _11629_ (.A1(_05036_),
    .A2(\registers[18][30] ),
    .ZN(_05044_));
 OAI21_X1 _11630_ (.A(_05043_),
    .B1(_05044_),
    .B2(_05038_),
    .ZN(_00704_));
 NAND2_X1 _11631_ (.A1(_04774_),
    .A2(_05030_),
    .ZN(_05045_));
 NAND2_X1 _11632_ (.A1(_05036_),
    .A2(\registers[18][31] ),
    .ZN(_05046_));
 OAI21_X1 _11633_ (.A(_05045_),
    .B1(_05046_),
    .B2(_05038_),
    .ZN(_00705_));
 NAND2_X1 _11634_ (.A1(_04778_),
    .A2(_05030_),
    .ZN(_05047_));
 NAND2_X1 _11635_ (.A1(_05036_),
    .A2(\registers[18][3] ),
    .ZN(_05048_));
 OAI21_X1 _11636_ (.A(_05047_),
    .B1(_05048_),
    .B2(_05038_),
    .ZN(_00706_));
 NAND2_X1 _11637_ (.A1(_04781_),
    .A2(_05030_),
    .ZN(_05049_));
 NAND2_X1 _11638_ (.A1(_05036_),
    .A2(\registers[18][4] ),
    .ZN(_05050_));
 OAI21_X1 _11639_ (.A(_05049_),
    .B1(_05050_),
    .B2(_05038_),
    .ZN(_00707_));
 NAND2_X1 _11640_ (.A1(_04784_),
    .A2(_05030_),
    .ZN(_05051_));
 NAND2_X1 _11641_ (.A1(_05036_),
    .A2(\registers[18][5] ),
    .ZN(_05052_));
 OAI21_X1 _11642_ (.A(_05051_),
    .B1(_05052_),
    .B2(_05038_),
    .ZN(_00708_));
 NAND2_X1 _11643_ (.A1(_04787_),
    .A2(_04987_),
    .ZN(_05053_));
 NAND2_X1 _11644_ (.A1(_05036_),
    .A2(\registers[18][6] ),
    .ZN(_05054_));
 OAI21_X1 _11645_ (.A(_05053_),
    .B1(_05054_),
    .B2(_05038_),
    .ZN(_00709_));
 NAND2_X1 _11646_ (.A1(_04790_),
    .A2(_04987_),
    .ZN(_05055_));
 NAND2_X1 _11647_ (.A1(_05036_),
    .A2(\registers[18][7] ),
    .ZN(_05056_));
 OAI21_X1 _11648_ (.A(_05055_),
    .B1(_05056_),
    .B2(_05038_),
    .ZN(_00710_));
 NAND2_X1 _11649_ (.A1(_04793_),
    .A2(_04987_),
    .ZN(_05057_));
 CLKBUF_X3 _11650_ (.A(_04844_),
    .Z(_05058_));
 NAND2_X1 _11651_ (.A1(_05058_),
    .A2(\registers[18][8] ),
    .ZN(_05059_));
 OAI21_X1 _11652_ (.A(_05057_),
    .B1(_05059_),
    .B2(_04988_),
    .ZN(_00711_));
 NAND2_X1 _11653_ (.A1(_04796_),
    .A2(_04987_),
    .ZN(_05060_));
 NAND2_X1 _11654_ (.A1(_05058_),
    .A2(\registers[18][9] ),
    .ZN(_05061_));
 OAI21_X1 _11655_ (.A(_05060_),
    .B1(_05061_),
    .B2(_04988_),
    .ZN(_00712_));
 NOR4_X4 _11656_ (.A1(_01090_),
    .A2(_01738_),
    .A3(_01092_),
    .A4(_01340_),
    .ZN(_05062_));
 BUF_X4 _11657_ (.A(_05062_),
    .Z(_05063_));
 BUF_X4 _11658_ (.A(_05063_),
    .Z(_05064_));
 NAND2_X1 _11659_ (.A1(_04799_),
    .A2(_05064_),
    .ZN(_05065_));
 NAND2_X1 _11660_ (.A1(_05058_),
    .A2(\registers[19][0] ),
    .ZN(_05066_));
 CLKBUF_X3 _11661_ (.A(_05063_),
    .Z(_05067_));
 OAI21_X1 _11662_ (.A(_05065_),
    .B1(_05066_),
    .B2(_05067_),
    .ZN(_00713_));
 NAND2_X1 _11663_ (.A1(_04806_),
    .A2(_05064_),
    .ZN(_05068_));
 NAND2_X1 _11664_ (.A1(_05058_),
    .A2(\registers[19][10] ),
    .ZN(_05069_));
 OAI21_X1 _11665_ (.A(_05068_),
    .B1(_05069_),
    .B2(_05067_),
    .ZN(_00714_));
 NAND2_X1 _11666_ (.A1(_04809_),
    .A2(_05064_),
    .ZN(_05070_));
 NAND2_X1 _11667_ (.A1(_05058_),
    .A2(\registers[19][11] ),
    .ZN(_05071_));
 OAI21_X1 _11668_ (.A(_05070_),
    .B1(_05071_),
    .B2(_05067_),
    .ZN(_00715_));
 NAND2_X1 _11669_ (.A1(_04813_),
    .A2(_05064_),
    .ZN(_05072_));
 NAND2_X1 _11670_ (.A1(_05058_),
    .A2(\registers[19][12] ),
    .ZN(_05073_));
 OAI21_X1 _11671_ (.A(_05072_),
    .B1(_05073_),
    .B2(_05067_),
    .ZN(_00716_));
 NAND2_X1 _11672_ (.A1(_04816_),
    .A2(_05064_),
    .ZN(_05074_));
 NAND2_X1 _11673_ (.A1(_05058_),
    .A2(\registers[19][13] ),
    .ZN(_05075_));
 OAI21_X1 _11674_ (.A(_05074_),
    .B1(_05075_),
    .B2(_05067_),
    .ZN(_00717_));
 NAND2_X1 _11675_ (.A1(_04819_),
    .A2(_05064_),
    .ZN(_05076_));
 NAND2_X1 _11676_ (.A1(_05058_),
    .A2(\registers[19][14] ),
    .ZN(_05077_));
 OAI21_X1 _11677_ (.A(_05076_),
    .B1(_05077_),
    .B2(_05067_),
    .ZN(_00718_));
 NAND2_X1 _11678_ (.A1(_04822_),
    .A2(_05064_),
    .ZN(_05078_));
 NAND2_X1 _11679_ (.A1(_05058_),
    .A2(\registers[19][15] ),
    .ZN(_05079_));
 OAI21_X1 _11680_ (.A(_05078_),
    .B1(_05079_),
    .B2(_05067_),
    .ZN(_00719_));
 NAND2_X1 _11681_ (.A1(_04825_),
    .A2(_05064_),
    .ZN(_05080_));
 NAND2_X1 _11682_ (.A1(_05058_),
    .A2(\registers[19][16] ),
    .ZN(_05081_));
 OAI21_X1 _11683_ (.A(_05080_),
    .B1(_05081_),
    .B2(_05067_),
    .ZN(_00720_));
 BUF_X4 _11684_ (.A(_05063_),
    .Z(_05082_));
 NAND2_X1 _11685_ (.A1(_04828_),
    .A2(_05082_),
    .ZN(_05083_));
 CLKBUF_X3 _11686_ (.A(_04844_),
    .Z(_05084_));
 NAND2_X1 _11687_ (.A1(_05084_),
    .A2(\registers[19][17] ),
    .ZN(_05085_));
 OAI21_X1 _11688_ (.A(_05083_),
    .B1(_05085_),
    .B2(_05067_),
    .ZN(_00721_));
 NAND2_X1 _11689_ (.A1(_04832_),
    .A2(_05082_),
    .ZN(_05086_));
 NAND2_X1 _11690_ (.A1(_05084_),
    .A2(\registers[19][18] ),
    .ZN(_05087_));
 OAI21_X1 _11691_ (.A(_05086_),
    .B1(_05087_),
    .B2(_05067_),
    .ZN(_00722_));
 NAND2_X1 _11692_ (.A1(_04835_),
    .A2(_05082_),
    .ZN(_05088_));
 NAND2_X1 _11693_ (.A1(_05084_),
    .A2(\registers[19][19] ),
    .ZN(_05089_));
 CLKBUF_X3 _11694_ (.A(_05063_),
    .Z(_05090_));
 OAI21_X1 _11695_ (.A(_05088_),
    .B1(_05089_),
    .B2(_05090_),
    .ZN(_00723_));
 NAND2_X1 _11696_ (.A1(_04839_),
    .A2(_05082_),
    .ZN(_05091_));
 NAND2_X1 _11697_ (.A1(_05084_),
    .A2(\registers[19][1] ),
    .ZN(_05092_));
 OAI21_X1 _11698_ (.A(_05091_),
    .B1(_05092_),
    .B2(_05090_),
    .ZN(_00724_));
 NAND2_X1 _11699_ (.A1(_04842_),
    .A2(_05082_),
    .ZN(_05093_));
 NAND2_X1 _11700_ (.A1(_05084_),
    .A2(\registers[19][20] ),
    .ZN(_05094_));
 OAI21_X1 _11701_ (.A(_05093_),
    .B1(_05094_),
    .B2(_05090_),
    .ZN(_00725_));
 NAND2_X1 _11702_ (.A1(_04847_),
    .A2(_05082_),
    .ZN(_05095_));
 NAND2_X1 _11703_ (.A1(_05084_),
    .A2(\registers[19][21] ),
    .ZN(_05096_));
 OAI21_X1 _11704_ (.A(_05095_),
    .B1(_05096_),
    .B2(_05090_),
    .ZN(_00726_));
 NAND2_X1 _11705_ (.A1(_04850_),
    .A2(_05082_),
    .ZN(_05097_));
 NAND2_X1 _11706_ (.A1(_05084_),
    .A2(\registers[19][22] ),
    .ZN(_05098_));
 OAI21_X1 _11707_ (.A(_05097_),
    .B1(_05098_),
    .B2(_05090_),
    .ZN(_00727_));
 NAND2_X1 _11708_ (.A1(_04853_),
    .A2(_05082_),
    .ZN(_05099_));
 NAND2_X1 _11709_ (.A1(_05084_),
    .A2(\registers[19][23] ),
    .ZN(_05100_));
 OAI21_X1 _11710_ (.A(_05099_),
    .B1(_05100_),
    .B2(_05090_),
    .ZN(_00728_));
 NAND2_X1 _11711_ (.A1(_04856_),
    .A2(_05082_),
    .ZN(_05101_));
 NAND2_X1 _11712_ (.A1(_05084_),
    .A2(\registers[19][24] ),
    .ZN(_05102_));
 OAI21_X1 _11713_ (.A(_05101_),
    .B1(_05102_),
    .B2(_05090_),
    .ZN(_00729_));
 NAND2_X1 _11714_ (.A1(_04859_),
    .A2(_05082_),
    .ZN(_05103_));
 NAND2_X1 _11715_ (.A1(_05084_),
    .A2(\registers[19][25] ),
    .ZN(_05104_));
 OAI21_X1 _11716_ (.A(_05103_),
    .B1(_05104_),
    .B2(_05090_),
    .ZN(_00730_));
 BUF_X4 _11717_ (.A(_05063_),
    .Z(_05105_));
 NAND2_X1 _11718_ (.A1(_04862_),
    .A2(_05105_),
    .ZN(_05106_));
 CLKBUF_X3 _11719_ (.A(_04844_),
    .Z(_05107_));
 NAND2_X1 _11720_ (.A1(_05107_),
    .A2(\registers[19][26] ),
    .ZN(_05108_));
 OAI21_X1 _11721_ (.A(_05106_),
    .B1(_05108_),
    .B2(_05090_),
    .ZN(_00731_));
 NAND2_X1 _11722_ (.A1(_04866_),
    .A2(_05105_),
    .ZN(_05109_));
 NAND2_X1 _11723_ (.A1(_05107_),
    .A2(\registers[19][27] ),
    .ZN(_05110_));
 OAI21_X1 _11724_ (.A(_05109_),
    .B1(_05110_),
    .B2(_05090_),
    .ZN(_00732_));
 NAND2_X1 _11725_ (.A1(_04869_),
    .A2(_05105_),
    .ZN(_05111_));
 NAND2_X1 _11726_ (.A1(_05107_),
    .A2(\registers[19][28] ),
    .ZN(_05112_));
 CLKBUF_X3 _11727_ (.A(_05063_),
    .Z(_05113_));
 OAI21_X1 _11728_ (.A(_05111_),
    .B1(_05112_),
    .B2(_05113_),
    .ZN(_00733_));
 NAND2_X1 _11729_ (.A1(_04873_),
    .A2(_05105_),
    .ZN(_05114_));
 NAND2_X1 _11730_ (.A1(_05107_),
    .A2(\registers[19][29] ),
    .ZN(_05115_));
 OAI21_X1 _11731_ (.A(_05114_),
    .B1(_05115_),
    .B2(_05113_),
    .ZN(_00734_));
 NAND2_X1 _11732_ (.A1(_04876_),
    .A2(_05105_),
    .ZN(_05116_));
 NAND2_X1 _11733_ (.A1(_05107_),
    .A2(\registers[19][2] ),
    .ZN(_05117_));
 OAI21_X1 _11734_ (.A(_05116_),
    .B1(_05117_),
    .B2(_05113_),
    .ZN(_00735_));
 NAND2_X1 _11735_ (.A1(_04880_),
    .A2(_05105_),
    .ZN(_05118_));
 NAND2_X1 _11736_ (.A1(_05107_),
    .A2(\registers[19][30] ),
    .ZN(_05119_));
 OAI21_X1 _11737_ (.A(_05118_),
    .B1(_05119_),
    .B2(_05113_),
    .ZN(_00736_));
 NAND2_X1 _11738_ (.A1(_04774_),
    .A2(_05105_),
    .ZN(_05120_));
 NAND2_X1 _11739_ (.A1(_05107_),
    .A2(\registers[19][31] ),
    .ZN(_05121_));
 OAI21_X1 _11740_ (.A(_05120_),
    .B1(_05121_),
    .B2(_05113_),
    .ZN(_00737_));
 NAND2_X1 _11741_ (.A1(_04778_),
    .A2(_05105_),
    .ZN(_05122_));
 NAND2_X1 _11742_ (.A1(_05107_),
    .A2(\registers[19][3] ),
    .ZN(_05123_));
 OAI21_X1 _11743_ (.A(_05122_),
    .B1(_05123_),
    .B2(_05113_),
    .ZN(_00738_));
 NAND2_X1 _11744_ (.A1(_04781_),
    .A2(_05105_),
    .ZN(_05124_));
 NAND2_X1 _11745_ (.A1(_05107_),
    .A2(\registers[19][4] ),
    .ZN(_05125_));
 OAI21_X1 _11746_ (.A(_05124_),
    .B1(_05125_),
    .B2(_05113_),
    .ZN(_00739_));
 NAND2_X1 _11747_ (.A1(_04784_),
    .A2(_05105_),
    .ZN(_05126_));
 NAND2_X1 _11748_ (.A1(_05107_),
    .A2(\registers[19][5] ),
    .ZN(_05127_));
 OAI21_X1 _11749_ (.A(_05126_),
    .B1(_05127_),
    .B2(_05113_),
    .ZN(_00740_));
 NAND2_X1 _11750_ (.A1(_04787_),
    .A2(_05063_),
    .ZN(_05128_));
 BUF_X4 _11751_ (.A(_04844_),
    .Z(_05129_));
 NAND2_X1 _11752_ (.A1(_05129_),
    .A2(\registers[19][6] ),
    .ZN(_05130_));
 OAI21_X1 _11753_ (.A(_05128_),
    .B1(_05130_),
    .B2(_05113_),
    .ZN(_00741_));
 NAND2_X1 _11754_ (.A1(_04790_),
    .A2(_05063_),
    .ZN(_05131_));
 NAND2_X1 _11755_ (.A1(_05129_),
    .A2(\registers[19][7] ),
    .ZN(_05132_));
 OAI21_X1 _11756_ (.A(_05131_),
    .B1(_05132_),
    .B2(_05113_),
    .ZN(_00742_));
 NAND2_X1 _11757_ (.A1(_04793_),
    .A2(_05063_),
    .ZN(_05133_));
 NAND2_X1 _11758_ (.A1(_05129_),
    .A2(\registers[19][8] ),
    .ZN(_05134_));
 OAI21_X1 _11759_ (.A(_05133_),
    .B1(_05134_),
    .B2(_05064_),
    .ZN(_00743_));
 NAND2_X1 _11760_ (.A1(_04796_),
    .A2(_05063_),
    .ZN(_05135_));
 NAND2_X1 _11761_ (.A1(_05129_),
    .A2(\registers[19][9] ),
    .ZN(_05136_));
 OAI21_X1 _11762_ (.A(_05135_),
    .B1(_05136_),
    .B2(_05064_),
    .ZN(_00744_));
 NOR2_X1 _11763_ (.A1(_01098_),
    .A2(_01138_),
    .ZN(_05137_));
 CLKBUF_X3 _11764_ (.A(_05137_),
    .Z(_05138_));
 CLKBUF_X3 _11765_ (.A(_05138_),
    .Z(_05139_));
 NAND2_X1 _11766_ (.A1(_04799_),
    .A2(_05139_),
    .ZN(_05140_));
 NAND2_X1 _11767_ (.A1(_05129_),
    .A2(\registers[1][0] ),
    .ZN(_05141_));
 CLKBUF_X3 _11768_ (.A(_05138_),
    .Z(_05142_));
 OAI21_X1 _11769_ (.A(_05140_),
    .B1(_05141_),
    .B2(_05142_),
    .ZN(_00745_));
 NAND2_X1 _11770_ (.A1(_04806_),
    .A2(_05139_),
    .ZN(_05143_));
 NAND2_X1 _11771_ (.A1(_05129_),
    .A2(\registers[1][10] ),
    .ZN(_05144_));
 OAI21_X1 _11772_ (.A(_05143_),
    .B1(_05144_),
    .B2(_05142_),
    .ZN(_00746_));
 NAND2_X1 _11773_ (.A1(_04809_),
    .A2(_05139_),
    .ZN(_05145_));
 NAND2_X1 _11774_ (.A1(_05129_),
    .A2(\registers[1][11] ),
    .ZN(_05146_));
 OAI21_X1 _11775_ (.A(_05145_),
    .B1(_05146_),
    .B2(_05142_),
    .ZN(_00747_));
 NAND2_X1 _11776_ (.A1(_04813_),
    .A2(_05139_),
    .ZN(_05147_));
 NAND2_X1 _11777_ (.A1(_05129_),
    .A2(\registers[1][12] ),
    .ZN(_05148_));
 OAI21_X1 _11778_ (.A(_05147_),
    .B1(_05148_),
    .B2(_05142_),
    .ZN(_00748_));
 NAND2_X1 _11779_ (.A1(_04816_),
    .A2(_05139_),
    .ZN(_05149_));
 NAND2_X1 _11780_ (.A1(_05129_),
    .A2(\registers[1][13] ),
    .ZN(_05150_));
 OAI21_X1 _11781_ (.A(_05149_),
    .B1(_05150_),
    .B2(_05142_),
    .ZN(_00749_));
 NAND2_X1 _11782_ (.A1(_04819_),
    .A2(_05139_),
    .ZN(_05151_));
 NAND2_X1 _11783_ (.A1(_05129_),
    .A2(\registers[1][14] ),
    .ZN(_05152_));
 OAI21_X1 _11784_ (.A(_05151_),
    .B1(_05152_),
    .B2(_05142_),
    .ZN(_00750_));
 NAND2_X1 _11785_ (.A1(_04822_),
    .A2(_05139_),
    .ZN(_05153_));
 CLKBUF_X3 _11786_ (.A(_04844_),
    .Z(_05154_));
 NAND2_X1 _11787_ (.A1(_05154_),
    .A2(\registers[1][15] ),
    .ZN(_05155_));
 OAI21_X1 _11788_ (.A(_05153_),
    .B1(_05155_),
    .B2(_05142_),
    .ZN(_00751_));
 NAND2_X1 _11789_ (.A1(_04825_),
    .A2(_05139_),
    .ZN(_05156_));
 NAND2_X1 _11790_ (.A1(_05154_),
    .A2(\registers[1][16] ),
    .ZN(_05157_));
 OAI21_X1 _11791_ (.A(_05156_),
    .B1(_05157_),
    .B2(_05142_),
    .ZN(_00752_));
 CLKBUF_X3 _11792_ (.A(_05138_),
    .Z(_05158_));
 NAND2_X1 _11793_ (.A1(_04828_),
    .A2(_05158_),
    .ZN(_05159_));
 NAND2_X1 _11794_ (.A1(_05154_),
    .A2(\registers[1][17] ),
    .ZN(_05160_));
 OAI21_X1 _11795_ (.A(_05159_),
    .B1(_05160_),
    .B2(_05142_),
    .ZN(_00753_));
 NAND2_X1 _11796_ (.A1(_04832_),
    .A2(_05158_),
    .ZN(_05161_));
 NAND2_X1 _11797_ (.A1(_05154_),
    .A2(\registers[1][18] ),
    .ZN(_05162_));
 OAI21_X1 _11798_ (.A(_05161_),
    .B1(_05162_),
    .B2(_05142_),
    .ZN(_00754_));
 NAND2_X1 _11799_ (.A1(_04835_),
    .A2(_05158_),
    .ZN(_05163_));
 NAND2_X1 _11800_ (.A1(_05154_),
    .A2(\registers[1][19] ),
    .ZN(_05164_));
 CLKBUF_X3 _11801_ (.A(_05138_),
    .Z(_05165_));
 OAI21_X1 _11802_ (.A(_05163_),
    .B1(_05164_),
    .B2(_05165_),
    .ZN(_00755_));
 NAND2_X1 _11803_ (.A1(_04839_),
    .A2(_05158_),
    .ZN(_05166_));
 NAND2_X1 _11804_ (.A1(_05154_),
    .A2(\registers[1][1] ),
    .ZN(_05167_));
 OAI21_X1 _11805_ (.A(_05166_),
    .B1(_05167_),
    .B2(_05165_),
    .ZN(_00756_));
 NAND2_X1 _11806_ (.A1(_04842_),
    .A2(_05158_),
    .ZN(_05168_));
 NAND2_X1 _11807_ (.A1(_05154_),
    .A2(\registers[1][20] ),
    .ZN(_05169_));
 OAI21_X1 _11808_ (.A(_05168_),
    .B1(_05169_),
    .B2(_05165_),
    .ZN(_00757_));
 NAND2_X1 _11809_ (.A1(_04847_),
    .A2(_05158_),
    .ZN(_05170_));
 NAND2_X1 _11810_ (.A1(_05154_),
    .A2(\registers[1][21] ),
    .ZN(_05171_));
 OAI21_X1 _11811_ (.A(_05170_),
    .B1(_05171_),
    .B2(_05165_),
    .ZN(_00758_));
 NAND2_X1 _11812_ (.A1(_04850_),
    .A2(_05158_),
    .ZN(_05172_));
 NAND2_X1 _11813_ (.A1(_05154_),
    .A2(\registers[1][22] ),
    .ZN(_05173_));
 OAI21_X1 _11814_ (.A(_05172_),
    .B1(_05173_),
    .B2(_05165_),
    .ZN(_00759_));
 NAND2_X1 _11815_ (.A1(_04853_),
    .A2(_05158_),
    .ZN(_05174_));
 NAND2_X1 _11816_ (.A1(_05154_),
    .A2(\registers[1][23] ),
    .ZN(_05175_));
 OAI21_X1 _11817_ (.A(_05174_),
    .B1(_05175_),
    .B2(_05165_),
    .ZN(_00760_));
 NAND2_X1 _11818_ (.A1(_04856_),
    .A2(_05158_),
    .ZN(_05176_));
 BUF_X4 _11819_ (.A(_01103_),
    .Z(_05177_));
 CLKBUF_X3 _11820_ (.A(_05177_),
    .Z(_05178_));
 NAND2_X1 _11821_ (.A1(_05178_),
    .A2(\registers[1][24] ),
    .ZN(_05179_));
 OAI21_X1 _11822_ (.A(_05176_),
    .B1(_05179_),
    .B2(_05165_),
    .ZN(_00761_));
 NAND2_X1 _11823_ (.A1(_04859_),
    .A2(_05158_),
    .ZN(_05180_));
 NAND2_X1 _11824_ (.A1(_05178_),
    .A2(\registers[1][25] ),
    .ZN(_05181_));
 OAI21_X1 _11825_ (.A(_05180_),
    .B1(_05181_),
    .B2(_05165_),
    .ZN(_00762_));
 CLKBUF_X3 _11826_ (.A(_05138_),
    .Z(_05182_));
 NAND2_X1 _11827_ (.A1(_04862_),
    .A2(_05182_),
    .ZN(_05183_));
 NAND2_X1 _11828_ (.A1(_05178_),
    .A2(\registers[1][26] ),
    .ZN(_05184_));
 OAI21_X1 _11829_ (.A(_05183_),
    .B1(_05184_),
    .B2(_05165_),
    .ZN(_00763_));
 NAND2_X1 _11830_ (.A1(_04866_),
    .A2(_05182_),
    .ZN(_05185_));
 NAND2_X1 _11831_ (.A1(_05178_),
    .A2(\registers[1][27] ),
    .ZN(_05186_));
 OAI21_X1 _11832_ (.A(_05185_),
    .B1(_05186_),
    .B2(_05165_),
    .ZN(_00764_));
 NAND2_X1 _11833_ (.A1(_04869_),
    .A2(_05182_),
    .ZN(_05187_));
 NAND2_X1 _11834_ (.A1(_05178_),
    .A2(\registers[1][28] ),
    .ZN(_05188_));
 CLKBUF_X3 _11835_ (.A(_05138_),
    .Z(_05189_));
 OAI21_X1 _11836_ (.A(_05187_),
    .B1(_05188_),
    .B2(_05189_),
    .ZN(_00765_));
 NAND2_X1 _11837_ (.A1(_04873_),
    .A2(_05182_),
    .ZN(_05190_));
 NAND2_X1 _11838_ (.A1(_05178_),
    .A2(\registers[1][29] ),
    .ZN(_05191_));
 OAI21_X1 _11839_ (.A(_05190_),
    .B1(_05191_),
    .B2(_05189_),
    .ZN(_00766_));
 NAND2_X1 _11840_ (.A1(_04876_),
    .A2(_05182_),
    .ZN(_05192_));
 NAND2_X1 _11841_ (.A1(_05178_),
    .A2(\registers[1][2] ),
    .ZN(_05193_));
 OAI21_X1 _11842_ (.A(_05192_),
    .B1(_05193_),
    .B2(_05189_),
    .ZN(_00767_));
 NAND2_X1 _11843_ (.A1(_04880_),
    .A2(_05182_),
    .ZN(_05194_));
 NAND2_X1 _11844_ (.A1(_05178_),
    .A2(\registers[1][30] ),
    .ZN(_05195_));
 OAI21_X1 _11845_ (.A(_05194_),
    .B1(_05195_),
    .B2(_05189_),
    .ZN(_00768_));
 NAND2_X1 _11846_ (.A1(_04774_),
    .A2(_05182_),
    .ZN(_05196_));
 NAND2_X1 _11847_ (.A1(_05178_),
    .A2(\registers[1][31] ),
    .ZN(_05197_));
 OAI21_X1 _11848_ (.A(_05196_),
    .B1(_05197_),
    .B2(_05189_),
    .ZN(_00769_));
 NAND2_X1 _11849_ (.A1(_04778_),
    .A2(_05182_),
    .ZN(_05198_));
 NAND2_X1 _11850_ (.A1(_05178_),
    .A2(\registers[1][3] ),
    .ZN(_05199_));
 OAI21_X1 _11851_ (.A(_05198_),
    .B1(_05199_),
    .B2(_05189_),
    .ZN(_00770_));
 NAND2_X1 _11852_ (.A1(_04781_),
    .A2(_05182_),
    .ZN(_05200_));
 BUF_X4 _11853_ (.A(_05177_),
    .Z(_05201_));
 NAND2_X1 _11854_ (.A1(_05201_),
    .A2(\registers[1][4] ),
    .ZN(_05202_));
 OAI21_X1 _11855_ (.A(_05200_),
    .B1(_05202_),
    .B2(_05189_),
    .ZN(_00771_));
 NAND2_X1 _11856_ (.A1(_04784_),
    .A2(_05182_),
    .ZN(_05203_));
 NAND2_X1 _11857_ (.A1(_05201_),
    .A2(\registers[1][5] ),
    .ZN(_05204_));
 OAI21_X1 _11858_ (.A(_05203_),
    .B1(_05204_),
    .B2(_05189_),
    .ZN(_00772_));
 NAND2_X1 _11859_ (.A1(_04787_),
    .A2(_05138_),
    .ZN(_05205_));
 NAND2_X1 _11860_ (.A1(_05201_),
    .A2(\registers[1][6] ),
    .ZN(_05206_));
 OAI21_X1 _11861_ (.A(_05205_),
    .B1(_05206_),
    .B2(_05189_),
    .ZN(_00773_));
 NAND2_X1 _11862_ (.A1(_04790_),
    .A2(_05138_),
    .ZN(_05207_));
 NAND2_X1 _11863_ (.A1(_05201_),
    .A2(\registers[1][7] ),
    .ZN(_05208_));
 OAI21_X1 _11864_ (.A(_05207_),
    .B1(_05208_),
    .B2(_05189_),
    .ZN(_00774_));
 NAND2_X1 _11865_ (.A1(_04793_),
    .A2(_05138_),
    .ZN(_05209_));
 NAND2_X1 _11866_ (.A1(_05201_),
    .A2(\registers[1][8] ),
    .ZN(_05210_));
 OAI21_X1 _11867_ (.A(_05209_),
    .B1(_05210_),
    .B2(_05139_),
    .ZN(_00775_));
 NAND2_X1 _11868_ (.A1(_04796_),
    .A2(_05138_),
    .ZN(_05211_));
 NAND2_X1 _11869_ (.A1(_05201_),
    .A2(\registers[1][9] ),
    .ZN(_05212_));
 OAI21_X1 _11870_ (.A(_05211_),
    .B1(_05212_),
    .B2(_05139_),
    .ZN(_00776_));
 OR3_X2 _11871_ (.A1(net3),
    .A2(_01738_),
    .A3(_01494_),
    .ZN(_05213_));
 OR2_X1 _11872_ (.A1(_01737_),
    .A2(_05213_),
    .ZN(_05214_));
 CLKBUF_X3 _11873_ (.A(_05214_),
    .Z(_05215_));
 CLKBUF_X3 _11874_ (.A(_05215_),
    .Z(_05216_));
 NAND3_X1 _11875_ (.A1(_04979_),
    .A2(\registers[20][0] ),
    .A3(_05216_),
    .ZN(_05217_));
 CLKBUF_X3 _11876_ (.A(_05215_),
    .Z(_05218_));
 OAI21_X1 _11877_ (.A(_05217_),
    .B1(_05218_),
    .B2(_01424_),
    .ZN(_00777_));
 NAND3_X1 _11878_ (.A1(_04979_),
    .A2(\registers[20][10] ),
    .A3(_05216_),
    .ZN(_05219_));
 OAI21_X1 _11879_ (.A(_05219_),
    .B1(_05218_),
    .B2(_01426_),
    .ZN(_00778_));
 NAND3_X1 _11880_ (.A1(_04979_),
    .A2(\registers[20][11] ),
    .A3(_05216_),
    .ZN(_05220_));
 OAI21_X1 _11881_ (.A(_05220_),
    .B1(_05218_),
    .B2(_01428_),
    .ZN(_00779_));
 NAND3_X1 _11882_ (.A1(_04979_),
    .A2(\registers[20][12] ),
    .A3(_05216_),
    .ZN(_05221_));
 OAI21_X1 _11883_ (.A(_05221_),
    .B1(_05218_),
    .B2(_01430_),
    .ZN(_00780_));
 CLKBUF_X3 _11884_ (.A(_01104_),
    .Z(_05222_));
 NAND3_X1 _11885_ (.A1(_05222_),
    .A2(\registers[20][13] ),
    .A3(_05216_),
    .ZN(_05223_));
 OAI21_X1 _11886_ (.A(_05223_),
    .B1(_05218_),
    .B2(_01432_),
    .ZN(_00781_));
 NAND3_X1 _11887_ (.A1(_05222_),
    .A2(\registers[20][14] ),
    .A3(_05216_),
    .ZN(_05224_));
 OAI21_X1 _11888_ (.A(_05224_),
    .B1(_05218_),
    .B2(_01434_),
    .ZN(_00782_));
 NAND3_X1 _11889_ (.A1(_05222_),
    .A2(\registers[20][15] ),
    .A3(_05216_),
    .ZN(_05225_));
 OAI21_X1 _11890_ (.A(_05225_),
    .B1(_05218_),
    .B2(_01436_),
    .ZN(_00783_));
 NAND3_X1 _11891_ (.A1(_05222_),
    .A2(\registers[20][16] ),
    .A3(_05216_),
    .ZN(_05226_));
 OAI21_X1 _11892_ (.A(_05226_),
    .B1(_05218_),
    .B2(_01438_),
    .ZN(_00784_));
 CLKBUF_X3 _11893_ (.A(_05215_),
    .Z(_05227_));
 NAND3_X1 _11894_ (.A1(_05222_),
    .A2(\registers[20][17] ),
    .A3(_05227_),
    .ZN(_05228_));
 OAI21_X1 _11895_ (.A(_05228_),
    .B1(_05218_),
    .B2(_01441_),
    .ZN(_00785_));
 NAND3_X1 _11896_ (.A1(_05222_),
    .A2(\registers[20][18] ),
    .A3(_05227_),
    .ZN(_05229_));
 OAI21_X1 _11897_ (.A(_05229_),
    .B1(_05218_),
    .B2(_01443_),
    .ZN(_00786_));
 NAND3_X1 _11898_ (.A1(_05222_),
    .A2(\registers[20][19] ),
    .A3(_05227_),
    .ZN(_05230_));
 CLKBUF_X3 _11899_ (.A(_05215_),
    .Z(_05231_));
 OAI21_X1 _11900_ (.A(_05230_),
    .B1(_05231_),
    .B2(_01447_),
    .ZN(_00787_));
 NAND3_X1 _11901_ (.A1(_05222_),
    .A2(\registers[20][1] ),
    .A3(_05227_),
    .ZN(_05232_));
 OAI21_X1 _11902_ (.A(_05232_),
    .B1(_05231_),
    .B2(_01449_),
    .ZN(_00788_));
 NAND3_X1 _11903_ (.A1(_05222_),
    .A2(\registers[20][20] ),
    .A3(_05227_),
    .ZN(_05233_));
 OAI21_X1 _11904_ (.A(_05233_),
    .B1(_05231_),
    .B2(_01451_),
    .ZN(_00789_));
 NAND3_X1 _11905_ (.A1(_05222_),
    .A2(\registers[20][21] ),
    .A3(_05227_),
    .ZN(_05234_));
 OAI21_X1 _11906_ (.A(_05234_),
    .B1(_05231_),
    .B2(_01453_),
    .ZN(_00790_));
 CLKBUF_X3 _11907_ (.A(_01104_),
    .Z(_05235_));
 NAND3_X1 _11908_ (.A1(_05235_),
    .A2(\registers[20][22] ),
    .A3(_05227_),
    .ZN(_05236_));
 OAI21_X1 _11909_ (.A(_05236_),
    .B1(_05231_),
    .B2(_01455_),
    .ZN(_00791_));
 NAND3_X1 _11910_ (.A1(_05235_),
    .A2(\registers[20][23] ),
    .A3(_05227_),
    .ZN(_05237_));
 OAI21_X1 _11911_ (.A(_05237_),
    .B1(_05231_),
    .B2(_01457_),
    .ZN(_00792_));
 NAND3_X1 _11912_ (.A1(_05235_),
    .A2(\registers[20][24] ),
    .A3(_05227_),
    .ZN(_05238_));
 OAI21_X1 _11913_ (.A(_05238_),
    .B1(_05231_),
    .B2(_01459_),
    .ZN(_00793_));
 NAND3_X1 _11914_ (.A1(_05235_),
    .A2(\registers[20][25] ),
    .A3(_05227_),
    .ZN(_05239_));
 OAI21_X1 _11915_ (.A(_05239_),
    .B1(_05231_),
    .B2(_01461_),
    .ZN(_00794_));
 CLKBUF_X3 _11916_ (.A(_05215_),
    .Z(_05240_));
 NAND3_X1 _11917_ (.A1(_05235_),
    .A2(\registers[20][26] ),
    .A3(_05240_),
    .ZN(_05241_));
 OAI21_X1 _11918_ (.A(_05241_),
    .B1(_05231_),
    .B2(_01464_),
    .ZN(_00795_));
 NAND3_X1 _11919_ (.A1(_05235_),
    .A2(\registers[20][27] ),
    .A3(_05240_),
    .ZN(_05242_));
 OAI21_X1 _11920_ (.A(_05242_),
    .B1(_05231_),
    .B2(_01466_),
    .ZN(_00796_));
 NAND3_X1 _11921_ (.A1(_05235_),
    .A2(\registers[20][28] ),
    .A3(_05240_),
    .ZN(_05243_));
 CLKBUF_X3 _11922_ (.A(_05215_),
    .Z(_05244_));
 OAI21_X1 _11923_ (.A(_05243_),
    .B1(_05244_),
    .B2(_01470_),
    .ZN(_00797_));
 NAND3_X1 _11924_ (.A1(_05235_),
    .A2(\registers[20][29] ),
    .A3(_05240_),
    .ZN(_05245_));
 OAI21_X1 _11925_ (.A(_05245_),
    .B1(_05244_),
    .B2(_01472_),
    .ZN(_00798_));
 NAND3_X1 _11926_ (.A1(_05235_),
    .A2(\registers[20][2] ),
    .A3(_05240_),
    .ZN(_05246_));
 OAI21_X1 _11927_ (.A(_05246_),
    .B1(_05244_),
    .B2(_01474_),
    .ZN(_00799_));
 NAND3_X1 _11928_ (.A1(_05235_),
    .A2(\registers[20][30] ),
    .A3(_05240_),
    .ZN(_05247_));
 OAI21_X1 _11929_ (.A(_05247_),
    .B1(_05244_),
    .B2(_01476_),
    .ZN(_00800_));
 BUF_X4 _11930_ (.A(_01104_),
    .Z(_05248_));
 NAND3_X1 _11931_ (.A1(_05248_),
    .A2(\registers[20][31] ),
    .A3(_05240_),
    .ZN(_05249_));
 OAI21_X1 _11932_ (.A(_05249_),
    .B1(_05244_),
    .B2(_01478_),
    .ZN(_00801_));
 NAND3_X1 _11933_ (.A1(_05248_),
    .A2(\registers[20][3] ),
    .A3(_05240_),
    .ZN(_05250_));
 OAI21_X1 _11934_ (.A(_05250_),
    .B1(_05244_),
    .B2(_01480_),
    .ZN(_00802_));
 NAND3_X1 _11935_ (.A1(_05248_),
    .A2(\registers[20][4] ),
    .A3(_05240_),
    .ZN(_05251_));
 OAI21_X1 _11936_ (.A(_05251_),
    .B1(_05244_),
    .B2(_01482_),
    .ZN(_00803_));
 NAND3_X1 _11937_ (.A1(_05248_),
    .A2(\registers[20][5] ),
    .A3(_05240_),
    .ZN(_05252_));
 OAI21_X1 _11938_ (.A(_05252_),
    .B1(_05244_),
    .B2(_01484_),
    .ZN(_00804_));
 NAND3_X1 _11939_ (.A1(_05248_),
    .A2(\registers[20][6] ),
    .A3(_05215_),
    .ZN(_05253_));
 OAI21_X1 _11940_ (.A(_05253_),
    .B1(_05244_),
    .B2(_01486_),
    .ZN(_00805_));
 NAND3_X1 _11941_ (.A1(_05248_),
    .A2(\registers[20][7] ),
    .A3(_05215_),
    .ZN(_05254_));
 OAI21_X1 _11942_ (.A(_05254_),
    .B1(_05244_),
    .B2(_01488_),
    .ZN(_00806_));
 NAND3_X1 _11943_ (.A1(_05248_),
    .A2(\registers[20][8] ),
    .A3(_05215_),
    .ZN(_05255_));
 OAI21_X1 _11944_ (.A(_05255_),
    .B1(_05216_),
    .B2(_01491_),
    .ZN(_00807_));
 NAND3_X1 _11945_ (.A1(_05248_),
    .A2(\registers[20][9] ),
    .A3(_05215_),
    .ZN(_05256_));
 OAI21_X1 _11946_ (.A(_05256_),
    .B1(_05216_),
    .B2(_01493_),
    .ZN(_00808_));
 NOR2_X1 _11947_ (.A1(_01098_),
    .A2(_05213_),
    .ZN(_05257_));
 CLKBUF_X3 _11948_ (.A(_05257_),
    .Z(_05258_));
 CLKBUF_X3 _11949_ (.A(_05258_),
    .Z(_05259_));
 NAND2_X1 _11950_ (.A1(_04799_),
    .A2(_05259_),
    .ZN(_05260_));
 NAND2_X1 _11951_ (.A1(_05201_),
    .A2(\registers[21][0] ),
    .ZN(_05261_));
 CLKBUF_X3 _11952_ (.A(_05258_),
    .Z(_05262_));
 OAI21_X1 _11953_ (.A(_05260_),
    .B1(_05261_),
    .B2(_05262_),
    .ZN(_00809_));
 NAND2_X1 _11954_ (.A1(_04806_),
    .A2(_05259_),
    .ZN(_05263_));
 NAND2_X1 _11955_ (.A1(_05201_),
    .A2(\registers[21][10] ),
    .ZN(_05264_));
 OAI21_X1 _11956_ (.A(_05263_),
    .B1(_05264_),
    .B2(_05262_),
    .ZN(_00810_));
 NAND2_X1 _11957_ (.A1(_04809_),
    .A2(_05259_),
    .ZN(_05265_));
 NAND2_X1 _11958_ (.A1(_05201_),
    .A2(\registers[21][11] ),
    .ZN(_05266_));
 OAI21_X1 _11959_ (.A(_05265_),
    .B1(_05266_),
    .B2(_05262_),
    .ZN(_00811_));
 NAND2_X1 _11960_ (.A1(_04813_),
    .A2(_05259_),
    .ZN(_05267_));
 NAND2_X1 _11961_ (.A1(_05201_),
    .A2(\registers[21][12] ),
    .ZN(_05268_));
 OAI21_X1 _11962_ (.A(_05267_),
    .B1(_05268_),
    .B2(_05262_),
    .ZN(_00812_));
 NAND2_X1 _11963_ (.A1(_04816_),
    .A2(_05259_),
    .ZN(_05269_));
 CLKBUF_X3 _11964_ (.A(_05177_),
    .Z(_05270_));
 NAND2_X1 _11965_ (.A1(_05270_),
    .A2(\registers[21][13] ),
    .ZN(_05271_));
 OAI21_X1 _11966_ (.A(_05269_),
    .B1(_05271_),
    .B2(_05262_),
    .ZN(_00813_));
 NAND2_X1 _11967_ (.A1(_04819_),
    .A2(_05259_),
    .ZN(_05272_));
 NAND2_X1 _11968_ (.A1(_05270_),
    .A2(\registers[21][14] ),
    .ZN(_05273_));
 OAI21_X1 _11969_ (.A(_05272_),
    .B1(_05273_),
    .B2(_05262_),
    .ZN(_00814_));
 NAND2_X1 _11970_ (.A1(_04822_),
    .A2(_05259_),
    .ZN(_05274_));
 NAND2_X1 _11971_ (.A1(_05270_),
    .A2(\registers[21][15] ),
    .ZN(_05275_));
 OAI21_X1 _11972_ (.A(_05274_),
    .B1(_05275_),
    .B2(_05262_),
    .ZN(_00815_));
 NAND2_X1 _11973_ (.A1(_04825_),
    .A2(_05259_),
    .ZN(_05276_));
 NAND2_X1 _11974_ (.A1(_05270_),
    .A2(\registers[21][16] ),
    .ZN(_05277_));
 OAI21_X1 _11975_ (.A(_05276_),
    .B1(_05277_),
    .B2(_05262_),
    .ZN(_00816_));
 CLKBUF_X3 _11976_ (.A(_05258_),
    .Z(_05278_));
 NAND2_X1 _11977_ (.A1(_04828_),
    .A2(_05278_),
    .ZN(_05279_));
 NAND2_X1 _11978_ (.A1(_05270_),
    .A2(\registers[21][17] ),
    .ZN(_05280_));
 OAI21_X1 _11979_ (.A(_05279_),
    .B1(_05280_),
    .B2(_05262_),
    .ZN(_00817_));
 NAND2_X1 _11980_ (.A1(_04832_),
    .A2(_05278_),
    .ZN(_05281_));
 NAND2_X1 _11981_ (.A1(_05270_),
    .A2(\registers[21][18] ),
    .ZN(_05282_));
 OAI21_X1 _11982_ (.A(_05281_),
    .B1(_05282_),
    .B2(_05262_),
    .ZN(_00818_));
 NAND2_X1 _11983_ (.A1(_04835_),
    .A2(_05278_),
    .ZN(_05283_));
 NAND2_X1 _11984_ (.A1(_05270_),
    .A2(\registers[21][19] ),
    .ZN(_05284_));
 CLKBUF_X3 _11985_ (.A(_05258_),
    .Z(_05285_));
 OAI21_X1 _11986_ (.A(_05283_),
    .B1(_05284_),
    .B2(_05285_),
    .ZN(_00819_));
 NAND2_X1 _11987_ (.A1(_04839_),
    .A2(_05278_),
    .ZN(_05286_));
 NAND2_X1 _11988_ (.A1(_05270_),
    .A2(\registers[21][1] ),
    .ZN(_05287_));
 OAI21_X1 _11989_ (.A(_05286_),
    .B1(_05287_),
    .B2(_05285_),
    .ZN(_00820_));
 NAND2_X1 _11990_ (.A1(_04842_),
    .A2(_05278_),
    .ZN(_05288_));
 NAND2_X1 _11991_ (.A1(_05270_),
    .A2(\registers[21][20] ),
    .ZN(_05289_));
 OAI21_X1 _11992_ (.A(_05288_),
    .B1(_05289_),
    .B2(_05285_),
    .ZN(_00821_));
 NAND2_X1 _11993_ (.A1(_04847_),
    .A2(_05278_),
    .ZN(_05290_));
 NAND2_X1 _11994_ (.A1(_05270_),
    .A2(\registers[21][21] ),
    .ZN(_05291_));
 OAI21_X1 _11995_ (.A(_05290_),
    .B1(_05291_),
    .B2(_05285_),
    .ZN(_00822_));
 NAND2_X1 _11996_ (.A1(_04850_),
    .A2(_05278_),
    .ZN(_05292_));
 CLKBUF_X3 _11997_ (.A(_05177_),
    .Z(_05293_));
 NAND2_X1 _11998_ (.A1(_05293_),
    .A2(\registers[21][22] ),
    .ZN(_05294_));
 OAI21_X1 _11999_ (.A(_05292_),
    .B1(_05294_),
    .B2(_05285_),
    .ZN(_00823_));
 NAND2_X1 _12000_ (.A1(_04853_),
    .A2(_05278_),
    .ZN(_05295_));
 NAND2_X1 _12001_ (.A1(_05293_),
    .A2(\registers[21][23] ),
    .ZN(_05296_));
 OAI21_X1 _12002_ (.A(_05295_),
    .B1(_05296_),
    .B2(_05285_),
    .ZN(_00824_));
 NAND2_X1 _12003_ (.A1(_04856_),
    .A2(_05278_),
    .ZN(_05297_));
 NAND2_X1 _12004_ (.A1(_05293_),
    .A2(\registers[21][24] ),
    .ZN(_05298_));
 OAI21_X1 _12005_ (.A(_05297_),
    .B1(_05298_),
    .B2(_05285_),
    .ZN(_00825_));
 NAND2_X1 _12006_ (.A1(_04859_),
    .A2(_05278_),
    .ZN(_05299_));
 NAND2_X1 _12007_ (.A1(_05293_),
    .A2(\registers[21][25] ),
    .ZN(_05300_));
 OAI21_X1 _12008_ (.A(_05299_),
    .B1(_05300_),
    .B2(_05285_),
    .ZN(_00826_));
 CLKBUF_X3 _12009_ (.A(_05258_),
    .Z(_05301_));
 NAND2_X1 _12010_ (.A1(_04862_),
    .A2(_05301_),
    .ZN(_05302_));
 NAND2_X1 _12011_ (.A1(_05293_),
    .A2(\registers[21][26] ),
    .ZN(_05303_));
 OAI21_X1 _12012_ (.A(_05302_),
    .B1(_05303_),
    .B2(_05285_),
    .ZN(_00827_));
 NAND2_X1 _12013_ (.A1(_04866_),
    .A2(_05301_),
    .ZN(_05304_));
 NAND2_X1 _12014_ (.A1(_05293_),
    .A2(\registers[21][27] ),
    .ZN(_05305_));
 OAI21_X1 _12015_ (.A(_05304_),
    .B1(_05305_),
    .B2(_05285_),
    .ZN(_00828_));
 NAND2_X1 _12016_ (.A1(_04869_),
    .A2(_05301_),
    .ZN(_05306_));
 NAND2_X1 _12017_ (.A1(_05293_),
    .A2(\registers[21][28] ),
    .ZN(_05307_));
 CLKBUF_X3 _12018_ (.A(_05258_),
    .Z(_05308_));
 OAI21_X1 _12019_ (.A(_05306_),
    .B1(_05307_),
    .B2(_05308_),
    .ZN(_00829_));
 NAND2_X1 _12020_ (.A1(_04873_),
    .A2(_05301_),
    .ZN(_05309_));
 NAND2_X1 _12021_ (.A1(_05293_),
    .A2(\registers[21][29] ),
    .ZN(_05310_));
 OAI21_X1 _12022_ (.A(_05309_),
    .B1(_05310_),
    .B2(_05308_),
    .ZN(_00830_));
 NAND2_X1 _12023_ (.A1(_04876_),
    .A2(_05301_),
    .ZN(_05311_));
 NAND2_X1 _12024_ (.A1(_05293_),
    .A2(\registers[21][2] ),
    .ZN(_05312_));
 OAI21_X1 _12025_ (.A(_05311_),
    .B1(_05312_),
    .B2(_05308_),
    .ZN(_00831_));
 NAND2_X1 _12026_ (.A1(_04880_),
    .A2(_05301_),
    .ZN(_05313_));
 NAND2_X1 _12027_ (.A1(_05293_),
    .A2(\registers[21][30] ),
    .ZN(_05314_));
 OAI21_X1 _12028_ (.A(_05313_),
    .B1(_05314_),
    .B2(_05308_),
    .ZN(_00832_));
 NAND2_X1 _12029_ (.A1(_04774_),
    .A2(_05301_),
    .ZN(_05315_));
 BUF_X4 _12030_ (.A(_05177_),
    .Z(_05316_));
 NAND2_X1 _12031_ (.A1(_05316_),
    .A2(\registers[21][31] ),
    .ZN(_05317_));
 OAI21_X1 _12032_ (.A(_05315_),
    .B1(_05317_),
    .B2(_05308_),
    .ZN(_00833_));
 NAND2_X1 _12033_ (.A1(_04778_),
    .A2(_05301_),
    .ZN(_05318_));
 NAND2_X1 _12034_ (.A1(_05316_),
    .A2(\registers[21][3] ),
    .ZN(_05319_));
 OAI21_X1 _12035_ (.A(_05318_),
    .B1(_05319_),
    .B2(_05308_),
    .ZN(_00834_));
 NAND2_X1 _12036_ (.A1(_04781_),
    .A2(_05301_),
    .ZN(_05320_));
 NAND2_X1 _12037_ (.A1(_05316_),
    .A2(\registers[21][4] ),
    .ZN(_05321_));
 OAI21_X1 _12038_ (.A(_05320_),
    .B1(_05321_),
    .B2(_05308_),
    .ZN(_00835_));
 NAND2_X1 _12039_ (.A1(_04784_),
    .A2(_05301_),
    .ZN(_05322_));
 NAND2_X1 _12040_ (.A1(_05316_),
    .A2(\registers[21][5] ),
    .ZN(_05323_));
 OAI21_X1 _12041_ (.A(_05322_),
    .B1(_05323_),
    .B2(_05308_),
    .ZN(_00836_));
 NAND2_X1 _12042_ (.A1(_04787_),
    .A2(_05258_),
    .ZN(_05324_));
 NAND2_X1 _12043_ (.A1(_05316_),
    .A2(\registers[21][6] ),
    .ZN(_05325_));
 OAI21_X1 _12044_ (.A(_05324_),
    .B1(_05325_),
    .B2(_05308_),
    .ZN(_00837_));
 NAND2_X1 _12045_ (.A1(_04790_),
    .A2(_05258_),
    .ZN(_05326_));
 NAND2_X1 _12046_ (.A1(_05316_),
    .A2(\registers[21][7] ),
    .ZN(_05327_));
 OAI21_X1 _12047_ (.A(_05326_),
    .B1(_05327_),
    .B2(_05308_),
    .ZN(_00838_));
 NAND2_X1 _12048_ (.A1(_04793_),
    .A2(_05258_),
    .ZN(_05328_));
 NAND2_X1 _12049_ (.A1(_05316_),
    .A2(\registers[21][8] ),
    .ZN(_05329_));
 OAI21_X1 _12050_ (.A(_05328_),
    .B1(_05329_),
    .B2(_05259_),
    .ZN(_00839_));
 NAND2_X1 _12051_ (.A1(_04796_),
    .A2(_05258_),
    .ZN(_05330_));
 NAND2_X1 _12052_ (.A1(_05316_),
    .A2(\registers[21][9] ),
    .ZN(_05331_));
 OAI21_X1 _12053_ (.A(_05330_),
    .B1(_05331_),
    .B2(_05259_),
    .ZN(_00840_));
 NOR2_X1 _12054_ (.A1(_01141_),
    .A2(_05213_),
    .ZN(_05332_));
 CLKBUF_X3 _12055_ (.A(_05332_),
    .Z(_05333_));
 CLKBUF_X3 _12056_ (.A(_05333_),
    .Z(_05334_));
 NAND2_X1 _12057_ (.A1(_04799_),
    .A2(_05334_),
    .ZN(_05335_));
 NAND2_X1 _12058_ (.A1(_05316_),
    .A2(\registers[22][0] ),
    .ZN(_05336_));
 CLKBUF_X3 _12059_ (.A(_05333_),
    .Z(_05337_));
 OAI21_X1 _12060_ (.A(_05335_),
    .B1(_05336_),
    .B2(_05337_),
    .ZN(_00841_));
 NAND2_X1 _12061_ (.A1(_04806_),
    .A2(_05334_),
    .ZN(_05338_));
 NAND2_X1 _12062_ (.A1(_05316_),
    .A2(\registers[22][10] ),
    .ZN(_05339_));
 OAI21_X1 _12063_ (.A(_05338_),
    .B1(_05339_),
    .B2(_05337_),
    .ZN(_00842_));
 NAND2_X1 _12064_ (.A1(_04809_),
    .A2(_05334_),
    .ZN(_05340_));
 CLKBUF_X3 _12065_ (.A(_05177_),
    .Z(_05341_));
 NAND2_X1 _12066_ (.A1(_05341_),
    .A2(\registers[22][11] ),
    .ZN(_05342_));
 OAI21_X1 _12067_ (.A(_05340_),
    .B1(_05342_),
    .B2(_05337_),
    .ZN(_00843_));
 NAND2_X1 _12068_ (.A1(_04813_),
    .A2(_05334_),
    .ZN(_05343_));
 NAND2_X1 _12069_ (.A1(_05341_),
    .A2(\registers[22][12] ),
    .ZN(_05344_));
 OAI21_X1 _12070_ (.A(_05343_),
    .B1(_05344_),
    .B2(_05337_),
    .ZN(_00844_));
 NAND2_X1 _12071_ (.A1(_04816_),
    .A2(_05334_),
    .ZN(_05345_));
 NAND2_X1 _12072_ (.A1(_05341_),
    .A2(\registers[22][13] ),
    .ZN(_05346_));
 OAI21_X1 _12073_ (.A(_05345_),
    .B1(_05346_),
    .B2(_05337_),
    .ZN(_00845_));
 NAND2_X1 _12074_ (.A1(_04819_),
    .A2(_05334_),
    .ZN(_05347_));
 NAND2_X1 _12075_ (.A1(_05341_),
    .A2(\registers[22][14] ),
    .ZN(_05348_));
 OAI21_X1 _12076_ (.A(_05347_),
    .B1(_05348_),
    .B2(_05337_),
    .ZN(_00846_));
 NAND2_X1 _12077_ (.A1(_04822_),
    .A2(_05334_),
    .ZN(_05349_));
 NAND2_X1 _12078_ (.A1(_05341_),
    .A2(\registers[22][15] ),
    .ZN(_05350_));
 OAI21_X1 _12079_ (.A(_05349_),
    .B1(_05350_),
    .B2(_05337_),
    .ZN(_00847_));
 NAND2_X1 _12080_ (.A1(_04825_),
    .A2(_05334_),
    .ZN(_05351_));
 NAND2_X1 _12081_ (.A1(_05341_),
    .A2(\registers[22][16] ),
    .ZN(_05352_));
 OAI21_X1 _12082_ (.A(_05351_),
    .B1(_05352_),
    .B2(_05337_),
    .ZN(_00848_));
 CLKBUF_X3 _12083_ (.A(_05333_),
    .Z(_05353_));
 NAND2_X1 _12084_ (.A1(_04828_),
    .A2(_05353_),
    .ZN(_05354_));
 NAND2_X1 _12085_ (.A1(_05341_),
    .A2(\registers[22][17] ),
    .ZN(_05355_));
 OAI21_X1 _12086_ (.A(_05354_),
    .B1(_05355_),
    .B2(_05337_),
    .ZN(_00849_));
 NAND2_X1 _12087_ (.A1(_04832_),
    .A2(_05353_),
    .ZN(_05356_));
 NAND2_X1 _12088_ (.A1(_05341_),
    .A2(\registers[22][18] ),
    .ZN(_05357_));
 OAI21_X1 _12089_ (.A(_05356_),
    .B1(_05357_),
    .B2(_05337_),
    .ZN(_00850_));
 NAND2_X1 _12090_ (.A1(_04835_),
    .A2(_05353_),
    .ZN(_05358_));
 NAND2_X1 _12091_ (.A1(_05341_),
    .A2(\registers[22][19] ),
    .ZN(_05359_));
 CLKBUF_X3 _12092_ (.A(_05333_),
    .Z(_05360_));
 OAI21_X1 _12093_ (.A(_05358_),
    .B1(_05359_),
    .B2(_05360_),
    .ZN(_00851_));
 NAND2_X1 _12094_ (.A1(_04839_),
    .A2(_05353_),
    .ZN(_05361_));
 NAND2_X1 _12095_ (.A1(_05341_),
    .A2(\registers[22][1] ),
    .ZN(_05362_));
 OAI21_X1 _12096_ (.A(_05361_),
    .B1(_05362_),
    .B2(_05360_),
    .ZN(_00852_));
 NAND2_X1 _12097_ (.A1(_04842_),
    .A2(_05353_),
    .ZN(_05363_));
 CLKBUF_X3 _12098_ (.A(_05177_),
    .Z(_05364_));
 NAND2_X1 _12099_ (.A1(_05364_),
    .A2(\registers[22][20] ),
    .ZN(_05365_));
 OAI21_X1 _12100_ (.A(_05363_),
    .B1(_05365_),
    .B2(_05360_),
    .ZN(_00853_));
 NAND2_X1 _12101_ (.A1(_04847_),
    .A2(_05353_),
    .ZN(_05366_));
 NAND2_X1 _12102_ (.A1(_05364_),
    .A2(\registers[22][21] ),
    .ZN(_05367_));
 OAI21_X1 _12103_ (.A(_05366_),
    .B1(_05367_),
    .B2(_05360_),
    .ZN(_00854_));
 NAND2_X1 _12104_ (.A1(_04850_),
    .A2(_05353_),
    .ZN(_05368_));
 NAND2_X1 _12105_ (.A1(_05364_),
    .A2(\registers[22][22] ),
    .ZN(_05369_));
 OAI21_X1 _12106_ (.A(_05368_),
    .B1(_05369_),
    .B2(_05360_),
    .ZN(_00855_));
 NAND2_X1 _12107_ (.A1(_04853_),
    .A2(_05353_),
    .ZN(_05370_));
 NAND2_X1 _12108_ (.A1(_05364_),
    .A2(\registers[22][23] ),
    .ZN(_05371_));
 OAI21_X1 _12109_ (.A(_05370_),
    .B1(_05371_),
    .B2(_05360_),
    .ZN(_00856_));
 NAND2_X1 _12110_ (.A1(_04856_),
    .A2(_05353_),
    .ZN(_05372_));
 NAND2_X1 _12111_ (.A1(_05364_),
    .A2(\registers[22][24] ),
    .ZN(_05373_));
 OAI21_X1 _12112_ (.A(_05372_),
    .B1(_05373_),
    .B2(_05360_),
    .ZN(_00857_));
 NAND2_X1 _12113_ (.A1(_04859_),
    .A2(_05353_),
    .ZN(_05374_));
 NAND2_X1 _12114_ (.A1(_05364_),
    .A2(\registers[22][25] ),
    .ZN(_05375_));
 OAI21_X1 _12115_ (.A(_05374_),
    .B1(_05375_),
    .B2(_05360_),
    .ZN(_00858_));
 CLKBUF_X3 _12116_ (.A(_05333_),
    .Z(_05376_));
 NAND2_X1 _12117_ (.A1(_04862_),
    .A2(_05376_),
    .ZN(_05377_));
 NAND2_X1 _12118_ (.A1(_05364_),
    .A2(\registers[22][26] ),
    .ZN(_05378_));
 OAI21_X1 _12119_ (.A(_05377_),
    .B1(_05378_),
    .B2(_05360_),
    .ZN(_00859_));
 NAND2_X1 _12120_ (.A1(_04866_),
    .A2(_05376_),
    .ZN(_05379_));
 NAND2_X1 _12121_ (.A1(_05364_),
    .A2(\registers[22][27] ),
    .ZN(_05380_));
 OAI21_X1 _12122_ (.A(_05379_),
    .B1(_05380_),
    .B2(_05360_),
    .ZN(_00860_));
 NAND2_X1 _12123_ (.A1(_04869_),
    .A2(_05376_),
    .ZN(_05381_));
 NAND2_X1 _12124_ (.A1(_05364_),
    .A2(\registers[22][28] ),
    .ZN(_05382_));
 CLKBUF_X3 _12125_ (.A(_05333_),
    .Z(_05383_));
 OAI21_X1 _12126_ (.A(_05381_),
    .B1(_05382_),
    .B2(_05383_),
    .ZN(_00861_));
 NAND2_X1 _12127_ (.A1(_04873_),
    .A2(_05376_),
    .ZN(_05384_));
 NAND2_X1 _12128_ (.A1(_05364_),
    .A2(\registers[22][29] ),
    .ZN(_05385_));
 OAI21_X1 _12129_ (.A(_05384_),
    .B1(_05385_),
    .B2(_05383_),
    .ZN(_00862_));
 NAND2_X1 _12130_ (.A1(_04876_),
    .A2(_05376_),
    .ZN(_05386_));
 BUF_X4 _12131_ (.A(_05177_),
    .Z(_05387_));
 NAND2_X1 _12132_ (.A1(_05387_),
    .A2(\registers[22][2] ),
    .ZN(_05388_));
 OAI21_X1 _12133_ (.A(_05386_),
    .B1(_05388_),
    .B2(_05383_),
    .ZN(_00863_));
 NAND2_X1 _12134_ (.A1(_04880_),
    .A2(_05376_),
    .ZN(_05389_));
 NAND2_X1 _12135_ (.A1(_05387_),
    .A2(\registers[22][30] ),
    .ZN(_05390_));
 OAI21_X1 _12136_ (.A(_05389_),
    .B1(_05390_),
    .B2(_05383_),
    .ZN(_00864_));
 NAND2_X1 _12137_ (.A1(_04774_),
    .A2(_05376_),
    .ZN(_05391_));
 NAND2_X1 _12138_ (.A1(_05387_),
    .A2(\registers[22][31] ),
    .ZN(_05392_));
 OAI21_X1 _12139_ (.A(_05391_),
    .B1(_05392_),
    .B2(_05383_),
    .ZN(_00865_));
 NAND2_X1 _12140_ (.A1(_04778_),
    .A2(_05376_),
    .ZN(_05393_));
 NAND2_X1 _12141_ (.A1(_05387_),
    .A2(\registers[22][3] ),
    .ZN(_05394_));
 OAI21_X1 _12142_ (.A(_05393_),
    .B1(_05394_),
    .B2(_05383_),
    .ZN(_00866_));
 NAND2_X1 _12143_ (.A1(_04781_),
    .A2(_05376_),
    .ZN(_05395_));
 NAND2_X1 _12144_ (.A1(_05387_),
    .A2(\registers[22][4] ),
    .ZN(_05396_));
 OAI21_X1 _12145_ (.A(_05395_),
    .B1(_05396_),
    .B2(_05383_),
    .ZN(_00867_));
 NAND2_X1 _12146_ (.A1(_04784_),
    .A2(_05376_),
    .ZN(_05397_));
 NAND2_X1 _12147_ (.A1(_05387_),
    .A2(\registers[22][5] ),
    .ZN(_05398_));
 OAI21_X1 _12148_ (.A(_05397_),
    .B1(_05398_),
    .B2(_05383_),
    .ZN(_00868_));
 NAND2_X1 _12149_ (.A1(_04787_),
    .A2(_05333_),
    .ZN(_05399_));
 NAND2_X1 _12150_ (.A1(_05387_),
    .A2(\registers[22][6] ),
    .ZN(_05400_));
 OAI21_X1 _12151_ (.A(_05399_),
    .B1(_05400_),
    .B2(_05383_),
    .ZN(_00869_));
 NAND2_X1 _12152_ (.A1(_04790_),
    .A2(_05333_),
    .ZN(_05401_));
 NAND2_X1 _12153_ (.A1(_05387_),
    .A2(\registers[22][7] ),
    .ZN(_05402_));
 OAI21_X1 _12154_ (.A(_05401_),
    .B1(_05402_),
    .B2(_05383_),
    .ZN(_00870_));
 NAND2_X1 _12155_ (.A1(_04793_),
    .A2(_05333_),
    .ZN(_05403_));
 NAND2_X1 _12156_ (.A1(_05387_),
    .A2(\registers[22][8] ),
    .ZN(_05404_));
 OAI21_X1 _12157_ (.A(_05403_),
    .B1(_05404_),
    .B2(_05334_),
    .ZN(_00871_));
 NAND2_X1 _12158_ (.A1(_04796_),
    .A2(_05333_),
    .ZN(_05405_));
 NAND2_X1 _12159_ (.A1(_05387_),
    .A2(\registers[22][9] ),
    .ZN(_05406_));
 OAI21_X1 _12160_ (.A(_05405_),
    .B1(_05406_),
    .B2(_05334_),
    .ZN(_00872_));
 NOR2_X2 _12161_ (.A1(_01340_),
    .A2(_05213_),
    .ZN(_05407_));
 BUF_X4 _12162_ (.A(_05407_),
    .Z(_05408_));
 CLKBUF_X3 _12163_ (.A(_05408_),
    .Z(_05409_));
 NAND2_X1 _12164_ (.A1(_04799_),
    .A2(_05409_),
    .ZN(_05410_));
 CLKBUF_X3 _12165_ (.A(_05177_),
    .Z(_05411_));
 NAND2_X1 _12166_ (.A1(_05411_),
    .A2(\registers[23][0] ),
    .ZN(_05412_));
 CLKBUF_X3 _12167_ (.A(_05408_),
    .Z(_05413_));
 OAI21_X1 _12168_ (.A(_05410_),
    .B1(_05412_),
    .B2(_05413_),
    .ZN(_00873_));
 NAND2_X1 _12169_ (.A1(_04806_),
    .A2(_05409_),
    .ZN(_05414_));
 NAND2_X1 _12170_ (.A1(_05411_),
    .A2(\registers[23][10] ),
    .ZN(_05415_));
 OAI21_X1 _12171_ (.A(_05414_),
    .B1(_05415_),
    .B2(_05413_),
    .ZN(_00874_));
 NAND2_X1 _12172_ (.A1(_04809_),
    .A2(_05409_),
    .ZN(_05416_));
 NAND2_X1 _12173_ (.A1(_05411_),
    .A2(\registers[23][11] ),
    .ZN(_05417_));
 OAI21_X1 _12174_ (.A(_05416_),
    .B1(_05417_),
    .B2(_05413_),
    .ZN(_00875_));
 NAND2_X1 _12175_ (.A1(_04813_),
    .A2(_05409_),
    .ZN(_05418_));
 NAND2_X1 _12176_ (.A1(_05411_),
    .A2(\registers[23][12] ),
    .ZN(_05419_));
 OAI21_X1 _12177_ (.A(_05418_),
    .B1(_05419_),
    .B2(_05413_),
    .ZN(_00876_));
 NAND2_X1 _12178_ (.A1(_04816_),
    .A2(_05409_),
    .ZN(_05420_));
 NAND2_X1 _12179_ (.A1(_05411_),
    .A2(\registers[23][13] ),
    .ZN(_05421_));
 OAI21_X1 _12180_ (.A(_05420_),
    .B1(_05421_),
    .B2(_05413_),
    .ZN(_00877_));
 NAND2_X1 _12181_ (.A1(_04819_),
    .A2(_05409_),
    .ZN(_05422_));
 NAND2_X1 _12182_ (.A1(_05411_),
    .A2(\registers[23][14] ),
    .ZN(_05423_));
 OAI21_X1 _12183_ (.A(_05422_),
    .B1(_05423_),
    .B2(_05413_),
    .ZN(_00878_));
 NAND2_X1 _12184_ (.A1(_04822_),
    .A2(_05409_),
    .ZN(_05424_));
 NAND2_X1 _12185_ (.A1(_05411_),
    .A2(\registers[23][15] ),
    .ZN(_05425_));
 OAI21_X1 _12186_ (.A(_05424_),
    .B1(_05425_),
    .B2(_05413_),
    .ZN(_00879_));
 NAND2_X1 _12187_ (.A1(_04825_),
    .A2(_05409_),
    .ZN(_05426_));
 NAND2_X1 _12188_ (.A1(_05411_),
    .A2(\registers[23][16] ),
    .ZN(_05427_));
 OAI21_X1 _12189_ (.A(_05426_),
    .B1(_05427_),
    .B2(_05413_),
    .ZN(_00880_));
 CLKBUF_X3 _12190_ (.A(_05408_),
    .Z(_05428_));
 NAND2_X1 _12191_ (.A1(_04828_),
    .A2(_05428_),
    .ZN(_05429_));
 NAND2_X1 _12192_ (.A1(_05411_),
    .A2(\registers[23][17] ),
    .ZN(_05430_));
 OAI21_X1 _12193_ (.A(_05429_),
    .B1(_05430_),
    .B2(_05413_),
    .ZN(_00881_));
 NAND2_X1 _12194_ (.A1(_04832_),
    .A2(_05428_),
    .ZN(_05431_));
 NAND2_X1 _12195_ (.A1(_05411_),
    .A2(\registers[23][18] ),
    .ZN(_05432_));
 OAI21_X1 _12196_ (.A(_05431_),
    .B1(_05432_),
    .B2(_05413_),
    .ZN(_00882_));
 NAND2_X1 _12197_ (.A1(_04835_),
    .A2(_05428_),
    .ZN(_05433_));
 CLKBUF_X3 _12198_ (.A(_05177_),
    .Z(_05434_));
 NAND2_X1 _12199_ (.A1(_05434_),
    .A2(\registers[23][19] ),
    .ZN(_05435_));
 CLKBUF_X3 _12200_ (.A(_05408_),
    .Z(_05436_));
 OAI21_X1 _12201_ (.A(_05433_),
    .B1(_05435_),
    .B2(_05436_),
    .ZN(_00883_));
 NAND2_X1 _12202_ (.A1(_04839_),
    .A2(_05428_),
    .ZN(_05437_));
 NAND2_X1 _12203_ (.A1(_05434_),
    .A2(\registers[23][1] ),
    .ZN(_05438_));
 OAI21_X1 _12204_ (.A(_05437_),
    .B1(_05438_),
    .B2(_05436_),
    .ZN(_00884_));
 NAND2_X1 _12205_ (.A1(_04842_),
    .A2(_05428_),
    .ZN(_05439_));
 NAND2_X1 _12206_ (.A1(_05434_),
    .A2(\registers[23][20] ),
    .ZN(_05440_));
 OAI21_X1 _12207_ (.A(_05439_),
    .B1(_05440_),
    .B2(_05436_),
    .ZN(_00885_));
 NAND2_X1 _12208_ (.A1(_04847_),
    .A2(_05428_),
    .ZN(_05441_));
 NAND2_X1 _12209_ (.A1(_05434_),
    .A2(\registers[23][21] ),
    .ZN(_05442_));
 OAI21_X1 _12210_ (.A(_05441_),
    .B1(_05442_),
    .B2(_05436_),
    .ZN(_00886_));
 NAND2_X1 _12211_ (.A1(_04850_),
    .A2(_05428_),
    .ZN(_05443_));
 NAND2_X1 _12212_ (.A1(_05434_),
    .A2(\registers[23][22] ),
    .ZN(_05444_));
 OAI21_X1 _12213_ (.A(_05443_),
    .B1(_05444_),
    .B2(_05436_),
    .ZN(_00887_));
 NAND2_X1 _12214_ (.A1(_04853_),
    .A2(_05428_),
    .ZN(_05445_));
 NAND2_X1 _12215_ (.A1(_05434_),
    .A2(\registers[23][23] ),
    .ZN(_05446_));
 OAI21_X1 _12216_ (.A(_05445_),
    .B1(_05446_),
    .B2(_05436_),
    .ZN(_00888_));
 NAND2_X1 _12217_ (.A1(_04856_),
    .A2(_05428_),
    .ZN(_05447_));
 NAND2_X1 _12218_ (.A1(_05434_),
    .A2(\registers[23][24] ),
    .ZN(_05448_));
 OAI21_X1 _12219_ (.A(_05447_),
    .B1(_05448_),
    .B2(_05436_),
    .ZN(_00889_));
 NAND2_X1 _12220_ (.A1(_04859_),
    .A2(_05428_),
    .ZN(_05449_));
 NAND2_X1 _12221_ (.A1(_05434_),
    .A2(\registers[23][25] ),
    .ZN(_05450_));
 OAI21_X1 _12222_ (.A(_05449_),
    .B1(_05450_),
    .B2(_05436_),
    .ZN(_00890_));
 CLKBUF_X3 _12223_ (.A(_05408_),
    .Z(_05451_));
 NAND2_X1 _12224_ (.A1(_04862_),
    .A2(_05451_),
    .ZN(_05452_));
 NAND2_X1 _12225_ (.A1(_05434_),
    .A2(\registers[23][26] ),
    .ZN(_05453_));
 OAI21_X1 _12226_ (.A(_05452_),
    .B1(_05453_),
    .B2(_05436_),
    .ZN(_00891_));
 NAND2_X1 _12227_ (.A1(_04866_),
    .A2(_05451_),
    .ZN(_05454_));
 NAND2_X1 _12228_ (.A1(_05434_),
    .A2(\registers[23][27] ),
    .ZN(_05455_));
 OAI21_X1 _12229_ (.A(_05454_),
    .B1(_05455_),
    .B2(_05436_),
    .ZN(_00892_));
 NAND2_X1 _12230_ (.A1(_04869_),
    .A2(_05451_),
    .ZN(_05456_));
 BUF_X4 _12231_ (.A(_01103_),
    .Z(_05457_));
 BUF_X2 _12232_ (.A(_05457_),
    .Z(_05458_));
 NAND2_X1 _12233_ (.A1(_05458_),
    .A2(\registers[23][28] ),
    .ZN(_05459_));
 BUF_X2 _12234_ (.A(_05408_),
    .Z(_05460_));
 OAI21_X1 _12235_ (.A(_05456_),
    .B1(_05459_),
    .B2(_05460_),
    .ZN(_00893_));
 NAND2_X1 _12236_ (.A1(_04873_),
    .A2(_05451_),
    .ZN(_05461_));
 NAND2_X1 _12237_ (.A1(_05458_),
    .A2(\registers[23][29] ),
    .ZN(_05462_));
 OAI21_X1 _12238_ (.A(_05461_),
    .B1(_05462_),
    .B2(_05460_),
    .ZN(_00894_));
 NAND2_X1 _12239_ (.A1(_04876_),
    .A2(_05451_),
    .ZN(_05463_));
 NAND2_X1 _12240_ (.A1(_05458_),
    .A2(\registers[23][2] ),
    .ZN(_05464_));
 OAI21_X1 _12241_ (.A(_05463_),
    .B1(_05464_),
    .B2(_05460_),
    .ZN(_00895_));
 NAND2_X1 _12242_ (.A1(_04880_),
    .A2(_05451_),
    .ZN(_05465_));
 NAND2_X1 _12243_ (.A1(_05458_),
    .A2(\registers[23][30] ),
    .ZN(_05466_));
 OAI21_X1 _12244_ (.A(_05465_),
    .B1(_05466_),
    .B2(_05460_),
    .ZN(_00896_));
 NAND2_X1 _12245_ (.A1(_04774_),
    .A2(_05451_),
    .ZN(_05467_));
 NAND2_X1 _12246_ (.A1(_05458_),
    .A2(\registers[23][31] ),
    .ZN(_05468_));
 OAI21_X1 _12247_ (.A(_05467_),
    .B1(_05468_),
    .B2(_05460_),
    .ZN(_00897_));
 NAND2_X1 _12248_ (.A1(_04778_),
    .A2(_05451_),
    .ZN(_05469_));
 NAND2_X1 _12249_ (.A1(_05458_),
    .A2(\registers[23][3] ),
    .ZN(_05470_));
 OAI21_X1 _12250_ (.A(_05469_),
    .B1(_05470_),
    .B2(_05460_),
    .ZN(_00898_));
 NAND2_X1 _12251_ (.A1(_04781_),
    .A2(_05451_),
    .ZN(_05471_));
 NAND2_X1 _12252_ (.A1(_05458_),
    .A2(\registers[23][4] ),
    .ZN(_05472_));
 OAI21_X1 _12253_ (.A(_05471_),
    .B1(_05472_),
    .B2(_05460_),
    .ZN(_00899_));
 NAND2_X1 _12254_ (.A1(_04784_),
    .A2(_05451_),
    .ZN(_05473_));
 NAND2_X1 _12255_ (.A1(_05458_),
    .A2(\registers[23][5] ),
    .ZN(_05474_));
 OAI21_X1 _12256_ (.A(_05473_),
    .B1(_05474_),
    .B2(_05460_),
    .ZN(_00900_));
 NAND2_X1 _12257_ (.A1(_04787_),
    .A2(_05408_),
    .ZN(_05475_));
 NAND2_X1 _12258_ (.A1(_05458_),
    .A2(\registers[23][6] ),
    .ZN(_05476_));
 OAI21_X1 _12259_ (.A(_05475_),
    .B1(_05476_),
    .B2(_05460_),
    .ZN(_00901_));
 NAND2_X1 _12260_ (.A1(_04790_),
    .A2(_05408_),
    .ZN(_05477_));
 NAND2_X1 _12261_ (.A1(_05458_),
    .A2(\registers[23][7] ),
    .ZN(_05478_));
 OAI21_X1 _12262_ (.A(_05477_),
    .B1(_05478_),
    .B2(_05460_),
    .ZN(_00902_));
 NAND2_X1 _12263_ (.A1(_04793_),
    .A2(_05408_),
    .ZN(_05479_));
 BUF_X4 _12264_ (.A(_05457_),
    .Z(_05480_));
 NAND2_X1 _12265_ (.A1(_05480_),
    .A2(\registers[23][8] ),
    .ZN(_05481_));
 OAI21_X1 _12266_ (.A(_05479_),
    .B1(_05481_),
    .B2(_05409_),
    .ZN(_00903_));
 NAND2_X1 _12267_ (.A1(_04796_),
    .A2(_05408_),
    .ZN(_05482_));
 NAND2_X1 _12268_ (.A1(_05480_),
    .A2(\registers[23][9] ),
    .ZN(_05483_));
 OAI21_X1 _12269_ (.A(_05482_),
    .B1(_05483_),
    .B2(_05409_),
    .ZN(_00904_));
 NAND3_X1 _12270_ (.A1(_01090_),
    .A2(_01091_),
    .A3(_01494_),
    .ZN(_05484_));
 OR2_X1 _12271_ (.A1(_01737_),
    .A2(_05484_),
    .ZN(_05485_));
 CLKBUF_X3 _12272_ (.A(_05485_),
    .Z(_05486_));
 CLKBUF_X3 _12273_ (.A(_05486_),
    .Z(_05487_));
 NAND3_X1 _12274_ (.A1(_05248_),
    .A2(\registers[24][0] ),
    .A3(_05487_),
    .ZN(_05488_));
 CLKBUF_X3 _12275_ (.A(_05486_),
    .Z(_05489_));
 OAI21_X1 _12276_ (.A(_05488_),
    .B1(_05489_),
    .B2(_01424_),
    .ZN(_00905_));
 NAND3_X1 _12277_ (.A1(_05248_),
    .A2(\registers[24][10] ),
    .A3(_05487_),
    .ZN(_05490_));
 OAI21_X1 _12278_ (.A(_05490_),
    .B1(_05489_),
    .B2(_01426_),
    .ZN(_00906_));
 CLKBUF_X3 _12279_ (.A(_01104_),
    .Z(_05491_));
 NAND3_X1 _12280_ (.A1(_05491_),
    .A2(\registers[24][11] ),
    .A3(_05487_),
    .ZN(_05492_));
 OAI21_X1 _12281_ (.A(_05492_),
    .B1(_05489_),
    .B2(_01428_),
    .ZN(_00907_));
 NAND3_X1 _12282_ (.A1(_05491_),
    .A2(\registers[24][12] ),
    .A3(_05487_),
    .ZN(_05493_));
 OAI21_X1 _12283_ (.A(_05493_),
    .B1(_05489_),
    .B2(_01430_),
    .ZN(_00908_));
 NAND3_X1 _12284_ (.A1(_05491_),
    .A2(\registers[24][13] ),
    .A3(_05487_),
    .ZN(_05494_));
 OAI21_X1 _12285_ (.A(_05494_),
    .B1(_05489_),
    .B2(_01432_),
    .ZN(_00909_));
 NAND3_X1 _12286_ (.A1(_05491_),
    .A2(\registers[24][14] ),
    .A3(_05487_),
    .ZN(_05495_));
 OAI21_X1 _12287_ (.A(_05495_),
    .B1(_05489_),
    .B2(_01434_),
    .ZN(_00910_));
 NAND3_X1 _12288_ (.A1(_05491_),
    .A2(\registers[24][15] ),
    .A3(_05487_),
    .ZN(_05496_));
 OAI21_X1 _12289_ (.A(_05496_),
    .B1(_05489_),
    .B2(_01436_),
    .ZN(_00911_));
 NAND3_X1 _12290_ (.A1(_05491_),
    .A2(\registers[24][16] ),
    .A3(_05487_),
    .ZN(_05497_));
 OAI21_X1 _12291_ (.A(_05497_),
    .B1(_05489_),
    .B2(_01438_),
    .ZN(_00912_));
 CLKBUF_X3 _12292_ (.A(_05486_),
    .Z(_05498_));
 NAND3_X1 _12293_ (.A1(_05491_),
    .A2(\registers[24][17] ),
    .A3(_05498_),
    .ZN(_05499_));
 OAI21_X1 _12294_ (.A(_05499_),
    .B1(_05489_),
    .B2(_01441_),
    .ZN(_00913_));
 NAND3_X1 _12295_ (.A1(_05491_),
    .A2(\registers[24][18] ),
    .A3(_05498_),
    .ZN(_05500_));
 OAI21_X1 _12296_ (.A(_05500_),
    .B1(_05489_),
    .B2(_01443_),
    .ZN(_00914_));
 NAND3_X1 _12297_ (.A1(_05491_),
    .A2(\registers[24][19] ),
    .A3(_05498_),
    .ZN(_05501_));
 CLKBUF_X3 _12298_ (.A(_05486_),
    .Z(_05502_));
 OAI21_X1 _12299_ (.A(_05501_),
    .B1(_05502_),
    .B2(_01447_),
    .ZN(_00915_));
 NAND3_X1 _12300_ (.A1(_05491_),
    .A2(\registers[24][1] ),
    .A3(_05498_),
    .ZN(_05503_));
 OAI21_X1 _12301_ (.A(_05503_),
    .B1(_05502_),
    .B2(_01449_),
    .ZN(_00916_));
 BUF_X4 _12302_ (.A(_01104_),
    .Z(_05504_));
 NAND3_X1 _12303_ (.A1(_05504_),
    .A2(\registers[24][20] ),
    .A3(_05498_),
    .ZN(_05505_));
 OAI21_X1 _12304_ (.A(_05505_),
    .B1(_05502_),
    .B2(_01451_),
    .ZN(_00917_));
 NAND3_X1 _12305_ (.A1(_05504_),
    .A2(\registers[24][21] ),
    .A3(_05498_),
    .ZN(_05506_));
 OAI21_X1 _12306_ (.A(_05506_),
    .B1(_05502_),
    .B2(_01453_),
    .ZN(_00918_));
 NAND3_X1 _12307_ (.A1(_05504_),
    .A2(\registers[24][22] ),
    .A3(_05498_),
    .ZN(_05507_));
 OAI21_X1 _12308_ (.A(_05507_),
    .B1(_05502_),
    .B2(_01455_),
    .ZN(_00919_));
 NAND3_X1 _12309_ (.A1(_05504_),
    .A2(\registers[24][23] ),
    .A3(_05498_),
    .ZN(_05508_));
 OAI21_X1 _12310_ (.A(_05508_),
    .B1(_05502_),
    .B2(_01457_),
    .ZN(_00920_));
 NAND3_X1 _12311_ (.A1(_05504_),
    .A2(\registers[24][24] ),
    .A3(_05498_),
    .ZN(_05509_));
 OAI21_X1 _12312_ (.A(_05509_),
    .B1(_05502_),
    .B2(_01459_),
    .ZN(_00921_));
 NAND3_X1 _12313_ (.A1(_05504_),
    .A2(\registers[24][25] ),
    .A3(_05498_),
    .ZN(_05510_));
 OAI21_X1 _12314_ (.A(_05510_),
    .B1(_05502_),
    .B2(_01461_),
    .ZN(_00922_));
 CLKBUF_X3 _12315_ (.A(_05486_),
    .Z(_05511_));
 NAND3_X1 _12316_ (.A1(_05504_),
    .A2(\registers[24][26] ),
    .A3(_05511_),
    .ZN(_05512_));
 OAI21_X1 _12317_ (.A(_05512_),
    .B1(_05502_),
    .B2(_01464_),
    .ZN(_00923_));
 NAND3_X1 _12318_ (.A1(_05504_),
    .A2(\registers[24][27] ),
    .A3(_05511_),
    .ZN(_05513_));
 OAI21_X1 _12319_ (.A(_05513_),
    .B1(_05502_),
    .B2(_01466_),
    .ZN(_00924_));
 NAND3_X1 _12320_ (.A1(_05504_),
    .A2(\registers[24][28] ),
    .A3(_05511_),
    .ZN(_05514_));
 CLKBUF_X3 _12321_ (.A(_05486_),
    .Z(_05515_));
 OAI21_X1 _12322_ (.A(_05514_),
    .B1(_05515_),
    .B2(_01470_),
    .ZN(_00925_));
 NAND3_X1 _12323_ (.A1(_05504_),
    .A2(\registers[24][29] ),
    .A3(_05511_),
    .ZN(_05516_));
 OAI21_X1 _12324_ (.A(_05516_),
    .B1(_05515_),
    .B2(_01472_),
    .ZN(_00926_));
 BUF_X4 _12325_ (.A(_01104_),
    .Z(_05517_));
 NAND3_X1 _12326_ (.A1(_05517_),
    .A2(\registers[24][2] ),
    .A3(_05511_),
    .ZN(_05518_));
 OAI21_X1 _12327_ (.A(_05518_),
    .B1(_05515_),
    .B2(_01474_),
    .ZN(_00927_));
 NAND3_X1 _12328_ (.A1(_05517_),
    .A2(\registers[24][30] ),
    .A3(_05511_),
    .ZN(_05519_));
 OAI21_X1 _12329_ (.A(_05519_),
    .B1(_05515_),
    .B2(_01476_),
    .ZN(_00928_));
 NAND3_X1 _12330_ (.A1(_05517_),
    .A2(\registers[24][31] ),
    .A3(_05511_),
    .ZN(_05520_));
 OAI21_X1 _12331_ (.A(_05520_),
    .B1(_05515_),
    .B2(_01478_),
    .ZN(_00929_));
 NAND3_X1 _12332_ (.A1(_05517_),
    .A2(\registers[24][3] ),
    .A3(_05511_),
    .ZN(_05521_));
 OAI21_X1 _12333_ (.A(_05521_),
    .B1(_05515_),
    .B2(_01480_),
    .ZN(_00930_));
 NAND3_X1 _12334_ (.A1(_05517_),
    .A2(\registers[24][4] ),
    .A3(_05511_),
    .ZN(_05522_));
 OAI21_X1 _12335_ (.A(_05522_),
    .B1(_05515_),
    .B2(_01482_),
    .ZN(_00931_));
 NAND3_X1 _12336_ (.A1(_05517_),
    .A2(\registers[24][5] ),
    .A3(_05511_),
    .ZN(_05523_));
 OAI21_X1 _12337_ (.A(_05523_),
    .B1(_05515_),
    .B2(_01484_),
    .ZN(_00932_));
 NAND3_X1 _12338_ (.A1(_05517_),
    .A2(\registers[24][6] ),
    .A3(_05486_),
    .ZN(_05524_));
 OAI21_X1 _12339_ (.A(_05524_),
    .B1(_05515_),
    .B2(_01486_),
    .ZN(_00933_));
 NAND3_X1 _12340_ (.A1(_05517_),
    .A2(\registers[24][7] ),
    .A3(_05486_),
    .ZN(_05525_));
 OAI21_X1 _12341_ (.A(_05525_),
    .B1(_05515_),
    .B2(_01488_),
    .ZN(_00934_));
 NAND3_X1 _12342_ (.A1(_05517_),
    .A2(\registers[24][8] ),
    .A3(_05486_),
    .ZN(_05526_));
 OAI21_X1 _12343_ (.A(_05526_),
    .B1(_05487_),
    .B2(_01491_),
    .ZN(_00935_));
 NAND3_X1 _12344_ (.A1(_05517_),
    .A2(\registers[24][9] ),
    .A3(_05486_),
    .ZN(_05527_));
 OAI21_X1 _12345_ (.A(_05527_),
    .B1(_05487_),
    .B2(_01493_),
    .ZN(_00936_));
 NOR2_X1 _12346_ (.A1(_01098_),
    .A2(_05484_),
    .ZN(_05528_));
 BUF_X4 _12347_ (.A(_05528_),
    .Z(_05529_));
 CLKBUF_X3 _12348_ (.A(_05529_),
    .Z(_05530_));
 NAND2_X1 _12349_ (.A1(_04799_),
    .A2(_05530_),
    .ZN(_05531_));
 NAND2_X1 _12350_ (.A1(_05480_),
    .A2(\registers[25][0] ),
    .ZN(_05532_));
 CLKBUF_X3 _12351_ (.A(_05529_),
    .Z(_05533_));
 OAI21_X1 _12352_ (.A(_05531_),
    .B1(_05532_),
    .B2(_05533_),
    .ZN(_00937_));
 NAND2_X1 _12353_ (.A1(_04806_),
    .A2(_05530_),
    .ZN(_05534_));
 NAND2_X1 _12354_ (.A1(_05480_),
    .A2(\registers[25][10] ),
    .ZN(_05535_));
 OAI21_X1 _12355_ (.A(_05534_),
    .B1(_05535_),
    .B2(_05533_),
    .ZN(_00938_));
 NAND2_X1 _12356_ (.A1(_04809_),
    .A2(_05530_),
    .ZN(_05536_));
 NAND2_X1 _12357_ (.A1(_05480_),
    .A2(\registers[25][11] ),
    .ZN(_05537_));
 OAI21_X1 _12358_ (.A(_05536_),
    .B1(_05537_),
    .B2(_05533_),
    .ZN(_00939_));
 NAND2_X1 _12359_ (.A1(_04813_),
    .A2(_05530_),
    .ZN(_05538_));
 NAND2_X1 _12360_ (.A1(_05480_),
    .A2(\registers[25][12] ),
    .ZN(_05539_));
 OAI21_X1 _12361_ (.A(_05538_),
    .B1(_05539_),
    .B2(_05533_),
    .ZN(_00940_));
 NAND2_X1 _12362_ (.A1(_04816_),
    .A2(_05530_),
    .ZN(_05540_));
 NAND2_X1 _12363_ (.A1(_05480_),
    .A2(\registers[25][13] ),
    .ZN(_05541_));
 OAI21_X1 _12364_ (.A(_05540_),
    .B1(_05541_),
    .B2(_05533_),
    .ZN(_00941_));
 NAND2_X1 _12365_ (.A1(_04819_),
    .A2(_05530_),
    .ZN(_05542_));
 NAND2_X1 _12366_ (.A1(_05480_),
    .A2(\registers[25][14] ),
    .ZN(_05543_));
 OAI21_X1 _12367_ (.A(_05542_),
    .B1(_05543_),
    .B2(_05533_),
    .ZN(_00942_));
 NAND2_X1 _12368_ (.A1(_04822_),
    .A2(_05530_),
    .ZN(_05544_));
 NAND2_X1 _12369_ (.A1(_05480_),
    .A2(\registers[25][15] ),
    .ZN(_05545_));
 OAI21_X1 _12370_ (.A(_05544_),
    .B1(_05545_),
    .B2(_05533_),
    .ZN(_00943_));
 NAND2_X1 _12371_ (.A1(_04825_),
    .A2(_05530_),
    .ZN(_05546_));
 NAND2_X1 _12372_ (.A1(_05480_),
    .A2(\registers[25][16] ),
    .ZN(_05547_));
 OAI21_X1 _12373_ (.A(_05546_),
    .B1(_05547_),
    .B2(_05533_),
    .ZN(_00944_));
 CLKBUF_X3 _12374_ (.A(_05529_),
    .Z(_05548_));
 NAND2_X1 _12375_ (.A1(_04828_),
    .A2(_05548_),
    .ZN(_05549_));
 CLKBUF_X3 _12376_ (.A(_05457_),
    .Z(_05550_));
 NAND2_X1 _12377_ (.A1(_05550_),
    .A2(\registers[25][17] ),
    .ZN(_05551_));
 OAI21_X1 _12378_ (.A(_05549_),
    .B1(_05551_),
    .B2(_05533_),
    .ZN(_00945_));
 NAND2_X1 _12379_ (.A1(_04832_),
    .A2(_05548_),
    .ZN(_05552_));
 NAND2_X1 _12380_ (.A1(_05550_),
    .A2(\registers[25][18] ),
    .ZN(_05553_));
 OAI21_X1 _12381_ (.A(_05552_),
    .B1(_05553_),
    .B2(_05533_),
    .ZN(_00946_));
 NAND2_X1 _12382_ (.A1(_04835_),
    .A2(_05548_),
    .ZN(_05554_));
 NAND2_X1 _12383_ (.A1(_05550_),
    .A2(\registers[25][19] ),
    .ZN(_05555_));
 CLKBUF_X3 _12384_ (.A(_05529_),
    .Z(_05556_));
 OAI21_X1 _12385_ (.A(_05554_),
    .B1(_05555_),
    .B2(_05556_),
    .ZN(_00947_));
 NAND2_X1 _12386_ (.A1(_04839_),
    .A2(_05548_),
    .ZN(_05557_));
 NAND2_X1 _12387_ (.A1(_05550_),
    .A2(\registers[25][1] ),
    .ZN(_05558_));
 OAI21_X1 _12388_ (.A(_05557_),
    .B1(_05558_),
    .B2(_05556_),
    .ZN(_00948_));
 NAND2_X1 _12389_ (.A1(_04842_),
    .A2(_05548_),
    .ZN(_05559_));
 NAND2_X1 _12390_ (.A1(_05550_),
    .A2(\registers[25][20] ),
    .ZN(_05560_));
 OAI21_X1 _12391_ (.A(_05559_),
    .B1(_05560_),
    .B2(_05556_),
    .ZN(_00949_));
 NAND2_X1 _12392_ (.A1(_04847_),
    .A2(_05548_),
    .ZN(_05561_));
 NAND2_X1 _12393_ (.A1(_05550_),
    .A2(\registers[25][21] ),
    .ZN(_05562_));
 OAI21_X1 _12394_ (.A(_05561_),
    .B1(_05562_),
    .B2(_05556_),
    .ZN(_00950_));
 NAND2_X1 _12395_ (.A1(_04850_),
    .A2(_05548_),
    .ZN(_05563_));
 NAND2_X1 _12396_ (.A1(_05550_),
    .A2(\registers[25][22] ),
    .ZN(_05564_));
 OAI21_X1 _12397_ (.A(_05563_),
    .B1(_05564_),
    .B2(_05556_),
    .ZN(_00951_));
 NAND2_X1 _12398_ (.A1(_04853_),
    .A2(_05548_),
    .ZN(_05565_));
 NAND2_X1 _12399_ (.A1(_05550_),
    .A2(\registers[25][23] ),
    .ZN(_05566_));
 OAI21_X1 _12400_ (.A(_05565_),
    .B1(_05566_),
    .B2(_05556_),
    .ZN(_00952_));
 NAND2_X1 _12401_ (.A1(_04856_),
    .A2(_05548_),
    .ZN(_05567_));
 NAND2_X1 _12402_ (.A1(_05550_),
    .A2(\registers[25][24] ),
    .ZN(_05568_));
 OAI21_X1 _12403_ (.A(_05567_),
    .B1(_05568_),
    .B2(_05556_),
    .ZN(_00953_));
 NAND2_X1 _12404_ (.A1(_04859_),
    .A2(_05548_),
    .ZN(_05569_));
 NAND2_X1 _12405_ (.A1(_05550_),
    .A2(\registers[25][25] ),
    .ZN(_05570_));
 OAI21_X1 _12406_ (.A(_05569_),
    .B1(_05570_),
    .B2(_05556_),
    .ZN(_00954_));
 CLKBUF_X3 _12407_ (.A(_05529_),
    .Z(_05571_));
 NAND2_X1 _12408_ (.A1(_04862_),
    .A2(_05571_),
    .ZN(_05572_));
 CLKBUF_X3 _12409_ (.A(_05457_),
    .Z(_05573_));
 NAND2_X1 _12410_ (.A1(_05573_),
    .A2(\registers[25][26] ),
    .ZN(_05574_));
 OAI21_X1 _12411_ (.A(_05572_),
    .B1(_05574_),
    .B2(_05556_),
    .ZN(_00955_));
 NAND2_X1 _12412_ (.A1(_04866_),
    .A2(_05571_),
    .ZN(_05575_));
 NAND2_X1 _12413_ (.A1(_05573_),
    .A2(\registers[25][27] ),
    .ZN(_05576_));
 OAI21_X1 _12414_ (.A(_05575_),
    .B1(_05576_),
    .B2(_05556_),
    .ZN(_00956_));
 NAND2_X1 _12415_ (.A1(_04869_),
    .A2(_05571_),
    .ZN(_05577_));
 NAND2_X1 _12416_ (.A1(_05573_),
    .A2(\registers[25][28] ),
    .ZN(_05578_));
 CLKBUF_X3 _12417_ (.A(_05529_),
    .Z(_05579_));
 OAI21_X1 _12418_ (.A(_05577_),
    .B1(_05578_),
    .B2(_05579_),
    .ZN(_00957_));
 NAND2_X1 _12419_ (.A1(_04873_),
    .A2(_05571_),
    .ZN(_05580_));
 NAND2_X1 _12420_ (.A1(_05573_),
    .A2(\registers[25][29] ),
    .ZN(_05581_));
 OAI21_X1 _12421_ (.A(_05580_),
    .B1(_05581_),
    .B2(_05579_),
    .ZN(_00958_));
 NAND2_X1 _12422_ (.A1(_04876_),
    .A2(_05571_),
    .ZN(_05582_));
 NAND2_X1 _12423_ (.A1(_05573_),
    .A2(\registers[25][2] ),
    .ZN(_05583_));
 OAI21_X1 _12424_ (.A(_05582_),
    .B1(_05583_),
    .B2(_05579_),
    .ZN(_00959_));
 NAND2_X1 _12425_ (.A1(_04880_),
    .A2(_05571_),
    .ZN(_05584_));
 NAND2_X1 _12426_ (.A1(_05573_),
    .A2(\registers[25][30] ),
    .ZN(_05585_));
 OAI21_X1 _12427_ (.A(_05584_),
    .B1(_05585_),
    .B2(_05579_),
    .ZN(_00960_));
 NAND2_X1 _12428_ (.A1(_04774_),
    .A2(_05571_),
    .ZN(_05586_));
 NAND2_X1 _12429_ (.A1(_05573_),
    .A2(\registers[25][31] ),
    .ZN(_05587_));
 OAI21_X1 _12430_ (.A(_05586_),
    .B1(_05587_),
    .B2(_05579_),
    .ZN(_00961_));
 NAND2_X1 _12431_ (.A1(_04778_),
    .A2(_05571_),
    .ZN(_05588_));
 NAND2_X1 _12432_ (.A1(_05573_),
    .A2(\registers[25][3] ),
    .ZN(_05589_));
 OAI21_X1 _12433_ (.A(_05588_),
    .B1(_05589_),
    .B2(_05579_),
    .ZN(_00962_));
 NAND2_X1 _12434_ (.A1(_04781_),
    .A2(_05571_),
    .ZN(_05590_));
 NAND2_X1 _12435_ (.A1(_05573_),
    .A2(\registers[25][4] ),
    .ZN(_05591_));
 OAI21_X1 _12436_ (.A(_05590_),
    .B1(_05591_),
    .B2(_05579_),
    .ZN(_00963_));
 NAND2_X1 _12437_ (.A1(_04784_),
    .A2(_05571_),
    .ZN(_05592_));
 NAND2_X1 _12438_ (.A1(_05573_),
    .A2(\registers[25][5] ),
    .ZN(_05593_));
 OAI21_X1 _12439_ (.A(_05592_),
    .B1(_05593_),
    .B2(_05579_),
    .ZN(_00964_));
 NAND2_X1 _12440_ (.A1(_04787_),
    .A2(_05529_),
    .ZN(_05594_));
 BUF_X4 _12441_ (.A(_05457_),
    .Z(_05595_));
 NAND2_X1 _12442_ (.A1(_05595_),
    .A2(\registers[25][6] ),
    .ZN(_05596_));
 OAI21_X1 _12443_ (.A(_05594_),
    .B1(_05596_),
    .B2(_05579_),
    .ZN(_00965_));
 NAND2_X1 _12444_ (.A1(_04790_),
    .A2(_05529_),
    .ZN(_05597_));
 NAND2_X1 _12445_ (.A1(_05595_),
    .A2(\registers[25][7] ),
    .ZN(_05598_));
 OAI21_X1 _12446_ (.A(_05597_),
    .B1(_05598_),
    .B2(_05579_),
    .ZN(_00966_));
 NAND2_X1 _12447_ (.A1(_04793_),
    .A2(_05529_),
    .ZN(_05599_));
 NAND2_X1 _12448_ (.A1(_05595_),
    .A2(\registers[25][8] ),
    .ZN(_05600_));
 OAI21_X1 _12449_ (.A(_05599_),
    .B1(_05600_),
    .B2(_05530_),
    .ZN(_00967_));
 NAND2_X1 _12450_ (.A1(_04796_),
    .A2(_05529_),
    .ZN(_05601_));
 NAND2_X1 _12451_ (.A1(_05595_),
    .A2(\registers[25][9] ),
    .ZN(_05602_));
 OAI21_X1 _12452_ (.A(_05601_),
    .B1(_05602_),
    .B2(_05530_),
    .ZN(_00968_));
 NOR2_X1 _12453_ (.A1(_01141_),
    .A2(_05484_),
    .ZN(_05603_));
 CLKBUF_X3 _12454_ (.A(_05603_),
    .Z(_05604_));
 CLKBUF_X3 _12455_ (.A(_05604_),
    .Z(_05605_));
 NAND2_X1 _12456_ (.A1(_04799_),
    .A2(_05605_),
    .ZN(_05606_));
 NAND2_X1 _12457_ (.A1(_05595_),
    .A2(\registers[26][0] ),
    .ZN(_05607_));
 CLKBUF_X3 _12458_ (.A(_05604_),
    .Z(_05608_));
 OAI21_X1 _12459_ (.A(_05606_),
    .B1(_05607_),
    .B2(_05608_),
    .ZN(_00969_));
 NAND2_X1 _12460_ (.A1(_04806_),
    .A2(_05605_),
    .ZN(_05609_));
 NAND2_X1 _12461_ (.A1(_05595_),
    .A2(\registers[26][10] ),
    .ZN(_05610_));
 OAI21_X1 _12462_ (.A(_05609_),
    .B1(_05610_),
    .B2(_05608_),
    .ZN(_00970_));
 NAND2_X1 _12463_ (.A1(_04809_),
    .A2(_05605_),
    .ZN(_05611_));
 NAND2_X1 _12464_ (.A1(_05595_),
    .A2(\registers[26][11] ),
    .ZN(_05612_));
 OAI21_X1 _12465_ (.A(_05611_),
    .B1(_05612_),
    .B2(_05608_),
    .ZN(_00971_));
 NAND2_X1 _12466_ (.A1(_04813_),
    .A2(_05605_),
    .ZN(_05613_));
 NAND2_X1 _12467_ (.A1(_05595_),
    .A2(\registers[26][12] ),
    .ZN(_05614_));
 OAI21_X1 _12468_ (.A(_05613_),
    .B1(_05614_),
    .B2(_05608_),
    .ZN(_00972_));
 NAND2_X1 _12469_ (.A1(_04816_),
    .A2(_05605_),
    .ZN(_05615_));
 NAND2_X1 _12470_ (.A1(_05595_),
    .A2(\registers[26][13] ),
    .ZN(_05616_));
 OAI21_X1 _12471_ (.A(_05615_),
    .B1(_05616_),
    .B2(_05608_),
    .ZN(_00973_));
 NAND2_X1 _12472_ (.A1(_04819_),
    .A2(_05605_),
    .ZN(_05617_));
 NAND2_X1 _12473_ (.A1(_05595_),
    .A2(\registers[26][14] ),
    .ZN(_05618_));
 OAI21_X1 _12474_ (.A(_05617_),
    .B1(_05618_),
    .B2(_05608_),
    .ZN(_00974_));
 NAND2_X1 _12475_ (.A1(_04822_),
    .A2(_05605_),
    .ZN(_05619_));
 CLKBUF_X3 _12476_ (.A(_05457_),
    .Z(_05620_));
 NAND2_X1 _12477_ (.A1(_05620_),
    .A2(\registers[26][15] ),
    .ZN(_05621_));
 OAI21_X1 _12478_ (.A(_05619_),
    .B1(_05621_),
    .B2(_05608_),
    .ZN(_00975_));
 NAND2_X1 _12479_ (.A1(_04825_),
    .A2(_05605_),
    .ZN(_05622_));
 NAND2_X1 _12480_ (.A1(_05620_),
    .A2(\registers[26][16] ),
    .ZN(_05623_));
 OAI21_X1 _12481_ (.A(_05622_),
    .B1(_05623_),
    .B2(_05608_),
    .ZN(_00976_));
 CLKBUF_X3 _12482_ (.A(_05604_),
    .Z(_05624_));
 NAND2_X1 _12483_ (.A1(_04828_),
    .A2(_05624_),
    .ZN(_05625_));
 NAND2_X1 _12484_ (.A1(_05620_),
    .A2(\registers[26][17] ),
    .ZN(_05626_));
 OAI21_X1 _12485_ (.A(_05625_),
    .B1(_05626_),
    .B2(_05608_),
    .ZN(_00977_));
 NAND2_X1 _12486_ (.A1(_04832_),
    .A2(_05624_),
    .ZN(_05627_));
 NAND2_X1 _12487_ (.A1(_05620_),
    .A2(\registers[26][18] ),
    .ZN(_05628_));
 OAI21_X1 _12488_ (.A(_05627_),
    .B1(_05628_),
    .B2(_05608_),
    .ZN(_00978_));
 NAND2_X1 _12489_ (.A1(_04835_),
    .A2(_05624_),
    .ZN(_05629_));
 NAND2_X1 _12490_ (.A1(_05620_),
    .A2(\registers[26][19] ),
    .ZN(_05630_));
 CLKBUF_X3 _12491_ (.A(_05604_),
    .Z(_05631_));
 OAI21_X1 _12492_ (.A(_05629_),
    .B1(_05630_),
    .B2(_05631_),
    .ZN(_00979_));
 NAND2_X1 _12493_ (.A1(_04839_),
    .A2(_05624_),
    .ZN(_05632_));
 NAND2_X1 _12494_ (.A1(_05620_),
    .A2(\registers[26][1] ),
    .ZN(_05633_));
 OAI21_X1 _12495_ (.A(_05632_),
    .B1(_05633_),
    .B2(_05631_),
    .ZN(_00980_));
 NAND2_X1 _12496_ (.A1(_04842_),
    .A2(_05624_),
    .ZN(_05634_));
 NAND2_X1 _12497_ (.A1(_05620_),
    .A2(\registers[26][20] ),
    .ZN(_05635_));
 OAI21_X1 _12498_ (.A(_05634_),
    .B1(_05635_),
    .B2(_05631_),
    .ZN(_00981_));
 NAND2_X1 _12499_ (.A1(_04847_),
    .A2(_05624_),
    .ZN(_05636_));
 NAND2_X1 _12500_ (.A1(_05620_),
    .A2(\registers[26][21] ),
    .ZN(_05637_));
 OAI21_X1 _12501_ (.A(_05636_),
    .B1(_05637_),
    .B2(_05631_),
    .ZN(_00982_));
 NAND2_X1 _12502_ (.A1(_04850_),
    .A2(_05624_),
    .ZN(_05638_));
 NAND2_X1 _12503_ (.A1(_05620_),
    .A2(\registers[26][22] ),
    .ZN(_05639_));
 OAI21_X1 _12504_ (.A(_05638_),
    .B1(_05639_),
    .B2(_05631_),
    .ZN(_00983_));
 NAND2_X1 _12505_ (.A1(_04853_),
    .A2(_05624_),
    .ZN(_05640_));
 NAND2_X1 _12506_ (.A1(_05620_),
    .A2(\registers[26][23] ),
    .ZN(_05641_));
 OAI21_X1 _12507_ (.A(_05640_),
    .B1(_05641_),
    .B2(_05631_),
    .ZN(_00984_));
 NAND2_X1 _12508_ (.A1(_04856_),
    .A2(_05624_),
    .ZN(_05642_));
 CLKBUF_X3 _12509_ (.A(_05457_),
    .Z(_05643_));
 NAND2_X1 _12510_ (.A1(_05643_),
    .A2(\registers[26][24] ),
    .ZN(_05644_));
 OAI21_X1 _12511_ (.A(_05642_),
    .B1(_05644_),
    .B2(_05631_),
    .ZN(_00985_));
 NAND2_X1 _12512_ (.A1(_04859_),
    .A2(_05624_),
    .ZN(_05645_));
 NAND2_X1 _12513_ (.A1(_05643_),
    .A2(\registers[26][25] ),
    .ZN(_05646_));
 OAI21_X1 _12514_ (.A(_05645_),
    .B1(_05646_),
    .B2(_05631_),
    .ZN(_00986_));
 CLKBUF_X3 _12515_ (.A(_05604_),
    .Z(_05647_));
 NAND2_X1 _12516_ (.A1(_04862_),
    .A2(_05647_),
    .ZN(_05648_));
 NAND2_X1 _12517_ (.A1(_05643_),
    .A2(\registers[26][26] ),
    .ZN(_05649_));
 OAI21_X1 _12518_ (.A(_05648_),
    .B1(_05649_),
    .B2(_05631_),
    .ZN(_00987_));
 NAND2_X1 _12519_ (.A1(_04866_),
    .A2(_05647_),
    .ZN(_05650_));
 NAND2_X1 _12520_ (.A1(_05643_),
    .A2(\registers[26][27] ),
    .ZN(_05651_));
 OAI21_X1 _12521_ (.A(_05650_),
    .B1(_05651_),
    .B2(_05631_),
    .ZN(_00988_));
 NAND2_X1 _12522_ (.A1(_04869_),
    .A2(_05647_),
    .ZN(_05652_));
 NAND2_X1 _12523_ (.A1(_05643_),
    .A2(\registers[26][28] ),
    .ZN(_05653_));
 CLKBUF_X3 _12524_ (.A(_05604_),
    .Z(_05654_));
 OAI21_X1 _12525_ (.A(_05652_),
    .B1(_05653_),
    .B2(_05654_),
    .ZN(_00989_));
 NAND2_X1 _12526_ (.A1(_04873_),
    .A2(_05647_),
    .ZN(_05655_));
 NAND2_X1 _12527_ (.A1(_05643_),
    .A2(\registers[26][29] ),
    .ZN(_05656_));
 OAI21_X1 _12528_ (.A(_05655_),
    .B1(_05656_),
    .B2(_05654_),
    .ZN(_00990_));
 NAND2_X1 _12529_ (.A1(_04876_),
    .A2(_05647_),
    .ZN(_05657_));
 NAND2_X1 _12530_ (.A1(_05643_),
    .A2(\registers[26][2] ),
    .ZN(_05658_));
 OAI21_X1 _12531_ (.A(_05657_),
    .B1(_05658_),
    .B2(_05654_),
    .ZN(_00991_));
 NAND2_X1 _12532_ (.A1(_04880_),
    .A2(_05647_),
    .ZN(_05659_));
 NAND2_X1 _12533_ (.A1(_05643_),
    .A2(\registers[26][30] ),
    .ZN(_05660_));
 OAI21_X1 _12534_ (.A(_05659_),
    .B1(_05660_),
    .B2(_05654_),
    .ZN(_00992_));
 NAND2_X1 _12535_ (.A1(_04774_),
    .A2(_05647_),
    .ZN(_05661_));
 NAND2_X1 _12536_ (.A1(_05643_),
    .A2(\registers[26][31] ),
    .ZN(_05662_));
 OAI21_X1 _12537_ (.A(_05661_),
    .B1(_05662_),
    .B2(_05654_),
    .ZN(_00993_));
 NAND2_X1 _12538_ (.A1(_04778_),
    .A2(_05647_),
    .ZN(_05663_));
 NAND2_X1 _12539_ (.A1(_05643_),
    .A2(\registers[26][3] ),
    .ZN(_05664_));
 OAI21_X1 _12540_ (.A(_05663_),
    .B1(_05664_),
    .B2(_05654_),
    .ZN(_00994_));
 NAND2_X1 _12541_ (.A1(_04781_),
    .A2(_05647_),
    .ZN(_05665_));
 BUF_X4 _12542_ (.A(_05457_),
    .Z(_05666_));
 NAND2_X1 _12543_ (.A1(_05666_),
    .A2(\registers[26][4] ),
    .ZN(_05667_));
 OAI21_X1 _12544_ (.A(_05665_),
    .B1(_05667_),
    .B2(_05654_),
    .ZN(_00995_));
 NAND2_X1 _12545_ (.A1(_04784_),
    .A2(_05647_),
    .ZN(_05668_));
 NAND2_X1 _12546_ (.A1(_05666_),
    .A2(\registers[26][5] ),
    .ZN(_05669_));
 OAI21_X1 _12547_ (.A(_05668_),
    .B1(_05669_),
    .B2(_05654_),
    .ZN(_00996_));
 NAND2_X1 _12548_ (.A1(_04787_),
    .A2(_05604_),
    .ZN(_05670_));
 NAND2_X1 _12549_ (.A1(_05666_),
    .A2(\registers[26][6] ),
    .ZN(_05671_));
 OAI21_X1 _12550_ (.A(_05670_),
    .B1(_05671_),
    .B2(_05654_),
    .ZN(_00997_));
 NAND2_X1 _12551_ (.A1(_04790_),
    .A2(_05604_),
    .ZN(_05672_));
 NAND2_X1 _12552_ (.A1(_05666_),
    .A2(\registers[26][7] ),
    .ZN(_05673_));
 OAI21_X1 _12553_ (.A(_05672_),
    .B1(_05673_),
    .B2(_05654_),
    .ZN(_00998_));
 NAND2_X1 _12554_ (.A1(_04793_),
    .A2(_05604_),
    .ZN(_05674_));
 NAND2_X1 _12555_ (.A1(_05666_),
    .A2(\registers[26][8] ),
    .ZN(_05675_));
 OAI21_X1 _12556_ (.A(_05674_),
    .B1(_05675_),
    .B2(_05605_),
    .ZN(_00999_));
 NAND2_X1 _12557_ (.A1(_04796_),
    .A2(_05604_),
    .ZN(_05676_));
 NAND2_X1 _12558_ (.A1(_05666_),
    .A2(\registers[26][9] ),
    .ZN(_05677_));
 OAI21_X1 _12559_ (.A(_05676_),
    .B1(_05677_),
    .B2(_05605_),
    .ZN(_01000_));
 NOR2_X1 _12560_ (.A1(_01340_),
    .A2(_05484_),
    .ZN(_05678_));
 BUF_X4 _12561_ (.A(_05678_),
    .Z(_05679_));
 CLKBUF_X3 _12562_ (.A(_05679_),
    .Z(_05680_));
 NAND2_X1 _12563_ (.A1(_04799_),
    .A2(_05680_),
    .ZN(_05681_));
 NAND2_X1 _12564_ (.A1(_05666_),
    .A2(\registers[27][0] ),
    .ZN(_05682_));
 CLKBUF_X3 _12565_ (.A(_05679_),
    .Z(_05683_));
 OAI21_X1 _12566_ (.A(_05681_),
    .B1(_05682_),
    .B2(_05683_),
    .ZN(_01001_));
 NAND2_X1 _12567_ (.A1(_04806_),
    .A2(_05680_),
    .ZN(_05684_));
 NAND2_X1 _12568_ (.A1(_05666_),
    .A2(\registers[27][10] ),
    .ZN(_05685_));
 OAI21_X1 _12569_ (.A(_05684_),
    .B1(_05685_),
    .B2(_05683_),
    .ZN(_01002_));
 NAND2_X1 _12570_ (.A1(_04809_),
    .A2(_05680_),
    .ZN(_05686_));
 NAND2_X1 _12571_ (.A1(_05666_),
    .A2(\registers[27][11] ),
    .ZN(_05687_));
 OAI21_X1 _12572_ (.A(_05686_),
    .B1(_05687_),
    .B2(_05683_),
    .ZN(_01003_));
 NAND2_X1 _12573_ (.A1(_04813_),
    .A2(_05680_),
    .ZN(_05688_));
 NAND2_X1 _12574_ (.A1(_05666_),
    .A2(\registers[27][12] ),
    .ZN(_05689_));
 OAI21_X1 _12575_ (.A(_05688_),
    .B1(_05689_),
    .B2(_05683_),
    .ZN(_01004_));
 NAND2_X1 _12576_ (.A1(_04816_),
    .A2(_05680_),
    .ZN(_05690_));
 CLKBUF_X3 _12577_ (.A(_05457_),
    .Z(_05691_));
 NAND2_X1 _12578_ (.A1(_05691_),
    .A2(\registers[27][13] ),
    .ZN(_05692_));
 OAI21_X1 _12579_ (.A(_05690_),
    .B1(_05692_),
    .B2(_05683_),
    .ZN(_01005_));
 NAND2_X1 _12580_ (.A1(_04819_),
    .A2(_05680_),
    .ZN(_05693_));
 NAND2_X1 _12581_ (.A1(_05691_),
    .A2(\registers[27][14] ),
    .ZN(_05694_));
 OAI21_X1 _12582_ (.A(_05693_),
    .B1(_05694_),
    .B2(_05683_),
    .ZN(_01006_));
 NAND2_X1 _12583_ (.A1(_04822_),
    .A2(_05680_),
    .ZN(_05695_));
 NAND2_X1 _12584_ (.A1(_05691_),
    .A2(\registers[27][15] ),
    .ZN(_05696_));
 OAI21_X1 _12585_ (.A(_05695_),
    .B1(_05696_),
    .B2(_05683_),
    .ZN(_01007_));
 NAND2_X1 _12586_ (.A1(_04825_),
    .A2(_05680_),
    .ZN(_05697_));
 NAND2_X1 _12587_ (.A1(_05691_),
    .A2(\registers[27][16] ),
    .ZN(_05698_));
 OAI21_X1 _12588_ (.A(_05697_),
    .B1(_05698_),
    .B2(_05683_),
    .ZN(_01008_));
 CLKBUF_X3 _12589_ (.A(_05679_),
    .Z(_05699_));
 NAND2_X1 _12590_ (.A1(_04828_),
    .A2(_05699_),
    .ZN(_05700_));
 NAND2_X1 _12591_ (.A1(_05691_),
    .A2(\registers[27][17] ),
    .ZN(_05701_));
 OAI21_X1 _12592_ (.A(_05700_),
    .B1(_05701_),
    .B2(_05683_),
    .ZN(_01009_));
 NAND2_X1 _12593_ (.A1(_04832_),
    .A2(_05699_),
    .ZN(_05702_));
 NAND2_X1 _12594_ (.A1(_05691_),
    .A2(\registers[27][18] ),
    .ZN(_05703_));
 OAI21_X1 _12595_ (.A(_05702_),
    .B1(_05703_),
    .B2(_05683_),
    .ZN(_01010_));
 NAND2_X1 _12596_ (.A1(_04835_),
    .A2(_05699_),
    .ZN(_05704_));
 NAND2_X1 _12597_ (.A1(_05691_),
    .A2(\registers[27][19] ),
    .ZN(_05705_));
 CLKBUF_X3 _12598_ (.A(_05679_),
    .Z(_05706_));
 OAI21_X1 _12599_ (.A(_05704_),
    .B1(_05705_),
    .B2(_05706_),
    .ZN(_01011_));
 NAND2_X1 _12600_ (.A1(_04839_),
    .A2(_05699_),
    .ZN(_05707_));
 NAND2_X1 _12601_ (.A1(_05691_),
    .A2(\registers[27][1] ),
    .ZN(_05708_));
 OAI21_X1 _12602_ (.A(_05707_),
    .B1(_05708_),
    .B2(_05706_),
    .ZN(_01012_));
 NAND2_X1 _12603_ (.A1(_04842_),
    .A2(_05699_),
    .ZN(_05709_));
 NAND2_X1 _12604_ (.A1(_05691_),
    .A2(\registers[27][20] ),
    .ZN(_05710_));
 OAI21_X1 _12605_ (.A(_05709_),
    .B1(_05710_),
    .B2(_05706_),
    .ZN(_01013_));
 NAND2_X1 _12606_ (.A1(_04847_),
    .A2(_05699_),
    .ZN(_05711_));
 NAND2_X1 _12607_ (.A1(_05691_),
    .A2(\registers[27][21] ),
    .ZN(_05712_));
 OAI21_X1 _12608_ (.A(_05711_),
    .B1(_05712_),
    .B2(_05706_),
    .ZN(_01014_));
 NAND2_X1 _12609_ (.A1(_04850_),
    .A2(_05699_),
    .ZN(_05713_));
 CLKBUF_X3 _12610_ (.A(_05457_),
    .Z(_05714_));
 NAND2_X1 _12611_ (.A1(_05714_),
    .A2(\registers[27][22] ),
    .ZN(_05715_));
 OAI21_X1 _12612_ (.A(_05713_),
    .B1(_05715_),
    .B2(_05706_),
    .ZN(_01015_));
 NAND2_X1 _12613_ (.A1(_04853_),
    .A2(_05699_),
    .ZN(_05716_));
 NAND2_X1 _12614_ (.A1(_05714_),
    .A2(\registers[27][23] ),
    .ZN(_05717_));
 OAI21_X1 _12615_ (.A(_05716_),
    .B1(_05717_),
    .B2(_05706_),
    .ZN(_01016_));
 NAND2_X1 _12616_ (.A1(_04856_),
    .A2(_05699_),
    .ZN(_05718_));
 NAND2_X1 _12617_ (.A1(_05714_),
    .A2(\registers[27][24] ),
    .ZN(_05719_));
 OAI21_X1 _12618_ (.A(_05718_),
    .B1(_05719_),
    .B2(_05706_),
    .ZN(_01017_));
 NAND2_X1 _12619_ (.A1(_04859_),
    .A2(_05699_),
    .ZN(_05720_));
 NAND2_X1 _12620_ (.A1(_05714_),
    .A2(\registers[27][25] ),
    .ZN(_05721_));
 OAI21_X1 _12621_ (.A(_05720_),
    .B1(_05721_),
    .B2(_05706_),
    .ZN(_01018_));
 CLKBUF_X3 _12622_ (.A(_05679_),
    .Z(_05722_));
 NAND2_X1 _12623_ (.A1(_04862_),
    .A2(_05722_),
    .ZN(_05723_));
 NAND2_X1 _12624_ (.A1(_05714_),
    .A2(\registers[27][26] ),
    .ZN(_05724_));
 OAI21_X1 _12625_ (.A(_05723_),
    .B1(_05724_),
    .B2(_05706_),
    .ZN(_01019_));
 NAND2_X1 _12626_ (.A1(_04866_),
    .A2(_05722_),
    .ZN(_05725_));
 NAND2_X1 _12627_ (.A1(_05714_),
    .A2(\registers[27][27] ),
    .ZN(_05726_));
 OAI21_X1 _12628_ (.A(_05725_),
    .B1(_05726_),
    .B2(_05706_),
    .ZN(_01020_));
 NAND2_X1 _12629_ (.A1(_04869_),
    .A2(_05722_),
    .ZN(_05727_));
 NAND2_X1 _12630_ (.A1(_05714_),
    .A2(\registers[27][28] ),
    .ZN(_05728_));
 CLKBUF_X3 _12631_ (.A(_05679_),
    .Z(_05729_));
 OAI21_X1 _12632_ (.A(_05727_),
    .B1(_05728_),
    .B2(_05729_),
    .ZN(_01021_));
 NAND2_X1 _12633_ (.A1(_04873_),
    .A2(_05722_),
    .ZN(_05730_));
 NAND2_X1 _12634_ (.A1(_05714_),
    .A2(\registers[27][29] ),
    .ZN(_05731_));
 OAI21_X1 _12635_ (.A(_05730_),
    .B1(_05731_),
    .B2(_05729_),
    .ZN(_01022_));
 NAND2_X1 _12636_ (.A1(_04876_),
    .A2(_05722_),
    .ZN(_05732_));
 NAND2_X1 _12637_ (.A1(_05714_),
    .A2(\registers[27][2] ),
    .ZN(_05733_));
 OAI21_X1 _12638_ (.A(_05732_),
    .B1(_05733_),
    .B2(_05729_),
    .ZN(_01023_));
 NAND2_X1 _12639_ (.A1(_04880_),
    .A2(_05722_),
    .ZN(_05734_));
 NAND2_X1 _12640_ (.A1(_05714_),
    .A2(\registers[27][30] ),
    .ZN(_05735_));
 OAI21_X1 _12641_ (.A(_05734_),
    .B1(_05735_),
    .B2(_05729_),
    .ZN(_01024_));
 NAND2_X1 _12642_ (.A1(_01088_),
    .A2(_05722_),
    .ZN(_05736_));
 BUF_X4 _12643_ (.A(_01416_),
    .Z(_05737_));
 NAND2_X1 _12644_ (.A1(_05737_),
    .A2(\registers[27][31] ),
    .ZN(_05738_));
 OAI21_X1 _12645_ (.A(_05736_),
    .B1(_05738_),
    .B2(_05729_),
    .ZN(_01025_));
 NAND2_X1 _12646_ (.A1(_01108_),
    .A2(_05722_),
    .ZN(_05739_));
 NAND2_X1 _12647_ (.A1(_05737_),
    .A2(\registers[27][3] ),
    .ZN(_05740_));
 OAI21_X1 _12648_ (.A(_05739_),
    .B1(_05740_),
    .B2(_05729_),
    .ZN(_01026_));
 NAND2_X1 _12649_ (.A1(_01112_),
    .A2(_05722_),
    .ZN(_05741_));
 NAND2_X1 _12650_ (.A1(_05737_),
    .A2(\registers[27][4] ),
    .ZN(_05742_));
 OAI21_X1 _12651_ (.A(_05741_),
    .B1(_05742_),
    .B2(_05729_),
    .ZN(_01027_));
 NAND2_X1 _12652_ (.A1(_01116_),
    .A2(_05722_),
    .ZN(_05743_));
 NAND2_X1 _12653_ (.A1(_05737_),
    .A2(\registers[27][5] ),
    .ZN(_05744_));
 OAI21_X1 _12654_ (.A(_05743_),
    .B1(_05744_),
    .B2(_05729_),
    .ZN(_01028_));
 NAND2_X1 _12655_ (.A1(_01120_),
    .A2(_05679_),
    .ZN(_05745_));
 NAND2_X1 _12656_ (.A1(_05737_),
    .A2(\registers[27][6] ),
    .ZN(_05746_));
 OAI21_X1 _12657_ (.A(_05745_),
    .B1(_05746_),
    .B2(_05729_),
    .ZN(_01029_));
 NAND2_X1 _12658_ (.A1(_01124_),
    .A2(_05679_),
    .ZN(_05747_));
 NAND2_X1 _12659_ (.A1(_05737_),
    .A2(\registers[27][7] ),
    .ZN(_05748_));
 OAI21_X1 _12660_ (.A(_05747_),
    .B1(_05748_),
    .B2(_05729_),
    .ZN(_01030_));
 NAND2_X1 _12661_ (.A1(_01128_),
    .A2(_05679_),
    .ZN(_05749_));
 NAND2_X1 _12662_ (.A1(_05737_),
    .A2(\registers[27][8] ),
    .ZN(_05750_));
 OAI21_X1 _12663_ (.A(_05749_),
    .B1(_05750_),
    .B2(_05680_),
    .ZN(_01031_));
 NAND2_X1 _12664_ (.A1(_01132_),
    .A2(_05679_),
    .ZN(_05751_));
 NAND2_X1 _12665_ (.A1(_05737_),
    .A2(\registers[27][9] ),
    .ZN(_05752_));
 OAI21_X1 _12666_ (.A(_05751_),
    .B1(_05752_),
    .B2(_05680_),
    .ZN(_01032_));
 NOR2_X1 _12667_ (.A1(_01093_),
    .A2(_01737_),
    .ZN(_05753_));
 CLKBUF_X3 _12668_ (.A(_05753_),
    .Z(_05754_));
 CLKBUF_X3 _12669_ (.A(_05754_),
    .Z(_05755_));
 NAND2_X1 _12670_ (.A1(_01136_),
    .A2(_05755_),
    .ZN(_05756_));
 NAND2_X1 _12671_ (.A1(_05737_),
    .A2(\registers[28][0] ),
    .ZN(_05757_));
 CLKBUF_X3 _12672_ (.A(_05754_),
    .Z(_05758_));
 OAI21_X1 _12673_ (.A(_05756_),
    .B1(_05757_),
    .B2(_05758_),
    .ZN(_01033_));
 NAND2_X1 _12674_ (.A1(_01148_),
    .A2(_05755_),
    .ZN(_05759_));
 NAND2_X1 _12675_ (.A1(_05737_),
    .A2(\registers[28][10] ),
    .ZN(_05760_));
 OAI21_X1 _12676_ (.A(_05759_),
    .B1(_05760_),
    .B2(_05758_),
    .ZN(_01034_));
 NAND2_X1 _12677_ (.A1(_01152_),
    .A2(_05755_),
    .ZN(_05761_));
 CLKBUF_X3 _12678_ (.A(_01416_),
    .Z(_05762_));
 NAND2_X1 _12679_ (.A1(_05762_),
    .A2(\registers[28][11] ),
    .ZN(_05763_));
 OAI21_X1 _12680_ (.A(_05761_),
    .B1(_05763_),
    .B2(_05758_),
    .ZN(_01035_));
 NAND2_X1 _12681_ (.A1(_01157_),
    .A2(_05755_),
    .ZN(_05764_));
 NAND2_X1 _12682_ (.A1(_05762_),
    .A2(\registers[28][12] ),
    .ZN(_05765_));
 OAI21_X1 _12683_ (.A(_05764_),
    .B1(_05765_),
    .B2(_05758_),
    .ZN(_01036_));
 NAND2_X1 _12684_ (.A1(_01161_),
    .A2(_05755_),
    .ZN(_05766_));
 NAND2_X1 _12685_ (.A1(_05762_),
    .A2(\registers[28][13] ),
    .ZN(_05767_));
 OAI21_X1 _12686_ (.A(_05766_),
    .B1(_05767_),
    .B2(_05758_),
    .ZN(_01037_));
 NAND2_X1 _12687_ (.A1(_01165_),
    .A2(_05755_),
    .ZN(_05768_));
 NAND2_X1 _12688_ (.A1(_05762_),
    .A2(\registers[28][14] ),
    .ZN(_05769_));
 OAI21_X1 _12689_ (.A(_05768_),
    .B1(_05769_),
    .B2(_05758_),
    .ZN(_01038_));
 NAND2_X1 _12690_ (.A1(_01169_),
    .A2(_05755_),
    .ZN(_05770_));
 NAND2_X1 _12691_ (.A1(_05762_),
    .A2(\registers[28][15] ),
    .ZN(_05771_));
 OAI21_X1 _12692_ (.A(_05770_),
    .B1(_05771_),
    .B2(_05758_),
    .ZN(_01039_));
 NAND2_X1 _12693_ (.A1(_01173_),
    .A2(_05755_),
    .ZN(_05772_));
 NAND2_X1 _12694_ (.A1(_05762_),
    .A2(\registers[28][16] ),
    .ZN(_05773_));
 OAI21_X1 _12695_ (.A(_05772_),
    .B1(_05773_),
    .B2(_05758_),
    .ZN(_01040_));
 CLKBUF_X3 _12696_ (.A(_05754_),
    .Z(_05774_));
 NAND2_X1 _12697_ (.A1(_01177_),
    .A2(_05774_),
    .ZN(_05775_));
 NAND2_X1 _12698_ (.A1(_05762_),
    .A2(\registers[28][17] ),
    .ZN(_05776_));
 OAI21_X1 _12699_ (.A(_05775_),
    .B1(_05776_),
    .B2(_05758_),
    .ZN(_01041_));
 NAND2_X1 _12700_ (.A1(_01182_),
    .A2(_05774_),
    .ZN(_05777_));
 NAND2_X1 _12701_ (.A1(_05762_),
    .A2(\registers[28][18] ),
    .ZN(_05778_));
 OAI21_X1 _12702_ (.A(_05777_),
    .B1(_05778_),
    .B2(_05758_),
    .ZN(_01042_));
 NAND2_X1 _12703_ (.A1(_01186_),
    .A2(_05774_),
    .ZN(_05779_));
 NAND2_X1 _12704_ (.A1(_05762_),
    .A2(\registers[28][19] ),
    .ZN(_05780_));
 CLKBUF_X3 _12705_ (.A(_05754_),
    .Z(_05781_));
 OAI21_X1 _12706_ (.A(_05779_),
    .B1(_05780_),
    .B2(_05781_),
    .ZN(_01043_));
 NAND2_X1 _12707_ (.A1(_01191_),
    .A2(_05774_),
    .ZN(_05782_));
 NAND2_X1 _12708_ (.A1(_05762_),
    .A2(\registers[28][1] ),
    .ZN(_05783_));
 OAI21_X1 _12709_ (.A(_05782_),
    .B1(_05783_),
    .B2(_05781_),
    .ZN(_01044_));
 NAND2_X1 _12710_ (.A1(_01195_),
    .A2(_05774_),
    .ZN(_05784_));
 CLKBUF_X3 _12711_ (.A(_01416_),
    .Z(_05785_));
 NAND2_X1 _12712_ (.A1(_05785_),
    .A2(\registers[28][20] ),
    .ZN(_05786_));
 OAI21_X1 _12713_ (.A(_05784_),
    .B1(_05786_),
    .B2(_05781_),
    .ZN(_01045_));
 NAND2_X1 _12714_ (.A1(_01200_),
    .A2(_05774_),
    .ZN(_05787_));
 NAND2_X1 _12715_ (.A1(_05785_),
    .A2(\registers[28][21] ),
    .ZN(_05788_));
 OAI21_X1 _12716_ (.A(_05787_),
    .B1(_05788_),
    .B2(_05781_),
    .ZN(_01046_));
 NAND2_X1 _12717_ (.A1(_01204_),
    .A2(_05774_),
    .ZN(_05789_));
 NAND2_X1 _12718_ (.A1(_05785_),
    .A2(\registers[28][22] ),
    .ZN(_05790_));
 OAI21_X1 _12719_ (.A(_05789_),
    .B1(_05790_),
    .B2(_05781_),
    .ZN(_01047_));
 NAND2_X1 _12720_ (.A1(_01208_),
    .A2(_05774_),
    .ZN(_05791_));
 NAND2_X1 _12721_ (.A1(_05785_),
    .A2(\registers[28][23] ),
    .ZN(_05792_));
 OAI21_X1 _12722_ (.A(_05791_),
    .B1(_05792_),
    .B2(_05781_),
    .ZN(_01048_));
 NAND2_X1 _12723_ (.A1(_01212_),
    .A2(_05774_),
    .ZN(_05793_));
 NAND2_X1 _12724_ (.A1(_05785_),
    .A2(\registers[28][24] ),
    .ZN(_05794_));
 OAI21_X1 _12725_ (.A(_05793_),
    .B1(_05794_),
    .B2(_05781_),
    .ZN(_01049_));
 NAND2_X1 _12726_ (.A1(_01216_),
    .A2(_05774_),
    .ZN(_05795_));
 NAND2_X1 _12727_ (.A1(_05785_),
    .A2(\registers[28][25] ),
    .ZN(_05796_));
 OAI21_X1 _12728_ (.A(_05795_),
    .B1(_05796_),
    .B2(_05781_),
    .ZN(_01050_));
 CLKBUF_X3 _12729_ (.A(_05754_),
    .Z(_05797_));
 NAND2_X1 _12730_ (.A1(_01220_),
    .A2(_05797_),
    .ZN(_05798_));
 NAND2_X1 _12731_ (.A1(_05785_),
    .A2(\registers[28][26] ),
    .ZN(_05799_));
 OAI21_X1 _12732_ (.A(_05798_),
    .B1(_05799_),
    .B2(_05781_),
    .ZN(_01051_));
 NAND2_X1 _12733_ (.A1(_01225_),
    .A2(_05797_),
    .ZN(_05800_));
 NAND2_X1 _12734_ (.A1(_05785_),
    .A2(\registers[28][27] ),
    .ZN(_05801_));
 OAI21_X1 _12735_ (.A(_05800_),
    .B1(_05801_),
    .B2(_05781_),
    .ZN(_01052_));
 NAND2_X1 _12736_ (.A1(_01229_),
    .A2(_05797_),
    .ZN(_05802_));
 NAND2_X1 _12737_ (.A1(_05785_),
    .A2(\registers[28][28] ),
    .ZN(_05803_));
 CLKBUF_X3 _12738_ (.A(_05754_),
    .Z(_05804_));
 OAI21_X1 _12739_ (.A(_05802_),
    .B1(_05803_),
    .B2(_05804_),
    .ZN(_01053_));
 NAND2_X1 _12740_ (.A1(_01234_),
    .A2(_05797_),
    .ZN(_05805_));
 NAND2_X1 _12741_ (.A1(_05785_),
    .A2(\registers[28][29] ),
    .ZN(_05806_));
 OAI21_X1 _12742_ (.A(_05805_),
    .B1(_05806_),
    .B2(_05804_),
    .ZN(_01054_));
 NAND2_X1 _12743_ (.A1(_01238_),
    .A2(_05797_),
    .ZN(_05807_));
 BUF_X4 _12744_ (.A(_01416_),
    .Z(_05808_));
 NAND2_X1 _12745_ (.A1(_05808_),
    .A2(\registers[28][2] ),
    .ZN(_05809_));
 OAI21_X1 _12746_ (.A(_05807_),
    .B1(_05809_),
    .B2(_05804_),
    .ZN(_01055_));
 NAND2_X1 _12747_ (.A1(_01243_),
    .A2(_05797_),
    .ZN(_05810_));
 NAND2_X1 _12748_ (.A1(_05808_),
    .A2(\registers[28][30] ),
    .ZN(_05811_));
 OAI21_X1 _12749_ (.A(_05810_),
    .B1(_05811_),
    .B2(_05804_),
    .ZN(_01056_));
 NAND2_X1 _12750_ (.A1(_01088_),
    .A2(_05797_),
    .ZN(_05812_));
 NAND2_X1 _12751_ (.A1(_05808_),
    .A2(\registers[28][31] ),
    .ZN(_05813_));
 OAI21_X1 _12752_ (.A(_05812_),
    .B1(_05813_),
    .B2(_05804_),
    .ZN(_01057_));
 NAND2_X1 _12753_ (.A1(_01108_),
    .A2(_05797_),
    .ZN(_05814_));
 NAND2_X1 _12754_ (.A1(_05808_),
    .A2(\registers[28][3] ),
    .ZN(_05815_));
 OAI21_X1 _12755_ (.A(_05814_),
    .B1(_05815_),
    .B2(_05804_),
    .ZN(_01058_));
 NAND2_X1 _12756_ (.A1(_01112_),
    .A2(_05797_),
    .ZN(_05816_));
 NAND2_X1 _12757_ (.A1(_05808_),
    .A2(\registers[28][4] ),
    .ZN(_05817_));
 OAI21_X1 _12758_ (.A(_05816_),
    .B1(_05817_),
    .B2(_05804_),
    .ZN(_01059_));
 NAND2_X1 _12759_ (.A1(_01116_),
    .A2(_05797_),
    .ZN(_05818_));
 NAND2_X1 _12760_ (.A1(_05808_),
    .A2(\registers[28][5] ),
    .ZN(_05819_));
 OAI21_X1 _12761_ (.A(_05818_),
    .B1(_05819_),
    .B2(_05804_),
    .ZN(_01060_));
 NAND2_X1 _12762_ (.A1(_01120_),
    .A2(_05754_),
    .ZN(_05820_));
 NAND2_X1 _12763_ (.A1(_05808_),
    .A2(\registers[28][6] ),
    .ZN(_05821_));
 OAI21_X1 _12764_ (.A(_05820_),
    .B1(_05821_),
    .B2(_05804_),
    .ZN(_01061_));
 NAND2_X1 _12765_ (.A1(_01124_),
    .A2(_05754_),
    .ZN(_05822_));
 NAND2_X1 _12766_ (.A1(_05808_),
    .A2(\registers[28][7] ),
    .ZN(_05823_));
 OAI21_X1 _12767_ (.A(_05822_),
    .B1(_05823_),
    .B2(_05804_),
    .ZN(_01062_));
 NAND2_X1 _12768_ (.A1(_01128_),
    .A2(_05754_),
    .ZN(_05824_));
 NAND2_X1 _12769_ (.A1(_05808_),
    .A2(\registers[28][8] ),
    .ZN(_05825_));
 OAI21_X1 _12770_ (.A(_05824_),
    .B1(_05825_),
    .B2(_05755_),
    .ZN(_01063_));
 NAND2_X1 _12771_ (.A1(_01132_),
    .A2(_05754_),
    .ZN(_05826_));
 NAND2_X1 _12772_ (.A1(_05808_),
    .A2(\registers[28][9] ),
    .ZN(_05827_));
 OAI21_X1 _12773_ (.A(_05826_),
    .B1(_05827_),
    .B2(_05755_),
    .ZN(_01064_));
 CLKBUF_X3 _12774_ (.A(_01100_),
    .Z(_05828_));
 NAND2_X1 _12775_ (.A1(_01136_),
    .A2(_05828_),
    .ZN(_05829_));
 CLKBUF_X3 _12776_ (.A(_01416_),
    .Z(_05830_));
 NAND2_X1 _12777_ (.A1(_05830_),
    .A2(\registers[29][0] ),
    .ZN(_05831_));
 OAI21_X1 _12778_ (.A(_05829_),
    .B1(_05831_),
    .B2(_01107_),
    .ZN(_01065_));
 NAND2_X1 _12779_ (.A1(_01148_),
    .A2(_05828_),
    .ZN(_05832_));
 NAND2_X1 _12780_ (.A1(_05830_),
    .A2(\registers[29][10] ),
    .ZN(_05833_));
 OAI21_X1 _12781_ (.A(_05832_),
    .B1(_05833_),
    .B2(_01107_),
    .ZN(_01066_));
 NAND2_X1 _12782_ (.A1(_01152_),
    .A2(_05828_),
    .ZN(_05834_));
 NAND2_X1 _12783_ (.A1(_05830_),
    .A2(\registers[29][11] ),
    .ZN(_05835_));
 CLKBUF_X3 _12784_ (.A(_01100_),
    .Z(_05836_));
 OAI21_X1 _12785_ (.A(_05834_),
    .B1(_05835_),
    .B2(_05836_),
    .ZN(_01067_));
 NAND2_X1 _12786_ (.A1(_01157_),
    .A2(_05828_),
    .ZN(_05837_));
 NAND2_X1 _12787_ (.A1(_05830_),
    .A2(\registers[29][12] ),
    .ZN(_05838_));
 OAI21_X1 _12788_ (.A(_05837_),
    .B1(_05838_),
    .B2(_05836_),
    .ZN(_01068_));
 NAND2_X1 _12789_ (.A1(_01161_),
    .A2(_05828_),
    .ZN(_05839_));
 NAND2_X1 _12790_ (.A1(_05830_),
    .A2(\registers[29][13] ),
    .ZN(_05840_));
 OAI21_X1 _12791_ (.A(_05839_),
    .B1(_05840_),
    .B2(_05836_),
    .ZN(_01069_));
 NAND2_X1 _12792_ (.A1(_01165_),
    .A2(_05828_),
    .ZN(_05841_));
 NAND2_X1 _12793_ (.A1(_05830_),
    .A2(\registers[29][14] ),
    .ZN(_05842_));
 OAI21_X1 _12794_ (.A(_05841_),
    .B1(_05842_),
    .B2(_05836_),
    .ZN(_01070_));
 NAND2_X1 _12795_ (.A1(_01169_),
    .A2(_05828_),
    .ZN(_05843_));
 NAND2_X1 _12796_ (.A1(_05830_),
    .A2(\registers[29][15] ),
    .ZN(_05844_));
 OAI21_X1 _12797_ (.A(_05843_),
    .B1(_05844_),
    .B2(_05836_),
    .ZN(_01071_));
 NAND2_X1 _12798_ (.A1(_01173_),
    .A2(_05828_),
    .ZN(_05845_));
 NAND2_X1 _12799_ (.A1(_05830_),
    .A2(\registers[29][16] ),
    .ZN(_05846_));
 OAI21_X1 _12800_ (.A(_05845_),
    .B1(_05846_),
    .B2(_05836_),
    .ZN(_01072_));
 NAND2_X1 _12801_ (.A1(_01177_),
    .A2(_05828_),
    .ZN(_05847_));
 NAND2_X1 _12802_ (.A1(_05830_),
    .A2(\registers[29][17] ),
    .ZN(_05848_));
 OAI21_X1 _12803_ (.A(_05847_),
    .B1(_05848_),
    .B2(_05836_),
    .ZN(_01073_));
 NAND2_X1 _12804_ (.A1(_01182_),
    .A2(_05828_),
    .ZN(_05849_));
 NAND2_X1 _12805_ (.A1(_05830_),
    .A2(\registers[29][18] ),
    .ZN(_05850_));
 OAI21_X1 _12806_ (.A(_05849_),
    .B1(_05850_),
    .B2(_05836_),
    .ZN(_01074_));
 CLKBUF_X3 _12807_ (.A(_01100_),
    .Z(_05851_));
 NAND2_X1 _12808_ (.A1(_01186_),
    .A2(_05851_),
    .ZN(_05852_));
 CLKBUF_X3 _12809_ (.A(_01416_),
    .Z(_05853_));
 NAND2_X1 _12810_ (.A1(_05853_),
    .A2(\registers[29][19] ),
    .ZN(_05854_));
 OAI21_X1 _12811_ (.A(_05852_),
    .B1(_05854_),
    .B2(_05836_),
    .ZN(_01075_));
 NAND2_X1 _12812_ (.A1(_01191_),
    .A2(_05851_),
    .ZN(_05855_));
 NAND2_X1 _12813_ (.A1(_05853_),
    .A2(\registers[29][1] ),
    .ZN(_05856_));
 OAI21_X1 _12814_ (.A(_05855_),
    .B1(_05856_),
    .B2(_05836_),
    .ZN(_01076_));
 NAND2_X1 _12815_ (.A1(_01195_),
    .A2(_05851_),
    .ZN(_05857_));
 NAND2_X1 _12816_ (.A1(_05853_),
    .A2(\registers[29][20] ),
    .ZN(_05858_));
 CLKBUF_X3 _12817_ (.A(_01100_),
    .Z(_05859_));
 OAI21_X1 _12818_ (.A(_05857_),
    .B1(_05858_),
    .B2(_05859_),
    .ZN(_01077_));
 NAND2_X1 _12819_ (.A1(_01200_),
    .A2(_05851_),
    .ZN(_05860_));
 NAND2_X1 _12820_ (.A1(_05853_),
    .A2(\registers[29][21] ),
    .ZN(_05861_));
 OAI21_X1 _12821_ (.A(_05860_),
    .B1(_05861_),
    .B2(_05859_),
    .ZN(_01078_));
 NAND2_X1 _12822_ (.A1(_01204_),
    .A2(_05851_),
    .ZN(_05862_));
 NAND2_X1 _12823_ (.A1(_05853_),
    .A2(\registers[29][22] ),
    .ZN(_05863_));
 OAI21_X1 _12824_ (.A(_05862_),
    .B1(_05863_),
    .B2(_05859_),
    .ZN(_01079_));
 NAND2_X1 _12825_ (.A1(_01208_),
    .A2(_05851_),
    .ZN(_05864_));
 NAND2_X1 _12826_ (.A1(_05853_),
    .A2(\registers[29][23] ),
    .ZN(_05865_));
 OAI21_X1 _12827_ (.A(_05864_),
    .B1(_05865_),
    .B2(_05859_),
    .ZN(_01080_));
 NAND2_X1 _12828_ (.A1(_01212_),
    .A2(_05851_),
    .ZN(_05866_));
 NAND2_X1 _12829_ (.A1(_05853_),
    .A2(\registers[29][24] ),
    .ZN(_05867_));
 OAI21_X1 _12830_ (.A(_05866_),
    .B1(_05867_),
    .B2(_05859_),
    .ZN(_01081_));
 NAND2_X1 _12831_ (.A1(_01216_),
    .A2(_05851_),
    .ZN(_05868_));
 NAND2_X1 _12832_ (.A1(_05853_),
    .A2(\registers[29][25] ),
    .ZN(_05869_));
 OAI21_X1 _12833_ (.A(_05868_),
    .B1(_05869_),
    .B2(_05859_),
    .ZN(_01082_));
 NAND2_X1 _12834_ (.A1(_01220_),
    .A2(_05851_),
    .ZN(_05870_));
 NAND2_X1 _12835_ (.A1(_05853_),
    .A2(\registers[29][26] ),
    .ZN(_05871_));
 OAI21_X1 _12836_ (.A(_05870_),
    .B1(_05871_),
    .B2(_05859_),
    .ZN(_01083_));
 NAND2_X1 _12837_ (.A1(_01225_),
    .A2(_05851_),
    .ZN(_05872_));
 NAND2_X1 _12838_ (.A1(_05853_),
    .A2(\registers[29][27] ),
    .ZN(_05873_));
 OAI21_X1 _12839_ (.A(_05872_),
    .B1(_05873_),
    .B2(_05859_),
    .ZN(_01084_));
 NAND2_X1 _12840_ (.A1(_01229_),
    .A2(_01100_),
    .ZN(_05874_));
 NAND2_X1 _12841_ (.A1(_01417_),
    .A2(\registers[29][28] ),
    .ZN(_05875_));
 OAI21_X1 _12842_ (.A(_05874_),
    .B1(_05875_),
    .B2(_05859_),
    .ZN(_01085_));
 NAND2_X1 _12843_ (.A1(_01234_),
    .A2(_01100_),
    .ZN(_05876_));
 NAND2_X1 _12844_ (.A1(_01417_),
    .A2(\registers[29][29] ),
    .ZN(_05877_));
 OAI21_X1 _12845_ (.A(_05876_),
    .B1(_05877_),
    .B2(_05859_),
    .ZN(_01086_));
 NAND2_X1 _12846_ (.A1(_01238_),
    .A2(_01100_),
    .ZN(_05878_));
 NAND2_X1 _12847_ (.A1(_01417_),
    .A2(\registers[29][2] ),
    .ZN(_05879_));
 OAI21_X1 _12848_ (.A(_05878_),
    .B1(_05879_),
    .B2(_01101_),
    .ZN(_01087_));
 NAND2_X1 _12849_ (.A1(_01243_),
    .A2(_01100_),
    .ZN(_05880_));
 NAND2_X1 _12850_ (.A1(_01417_),
    .A2(\registers[29][30] ),
    .ZN(_05881_));
 OAI21_X1 _12851_ (.A(_05880_),
    .B1(_05881_),
    .B2(_01101_),
    .ZN(_00000_));
 DFF_X2 \read_data1[0]$_SDFFCE_PN0P_  (.D(_00329_),
    .CK(clknet_leaf_134_clk),
    .Q(net5),
    .QN(_06969_));
 DFF_X2 \read_data1[10]$_SDFFCE_PN0P_  (.D(_00330_),
    .CK(clknet_leaf_133_clk),
    .Q(net6),
    .QN(_06968_));
 DFF_X2 \read_data1[11]$_SDFFCE_PN0P_  (.D(_00331_),
    .CK(clknet_leaf_123_clk),
    .Q(net7),
    .QN(_06967_));
 DFF_X2 \read_data1[12]$_SDFFCE_PN0P_  (.D(_00332_),
    .CK(clknet_leaf_123_clk),
    .Q(net8),
    .QN(_06966_));
 DFF_X2 \read_data1[13]$_SDFFCE_PN0P_  (.D(_00333_),
    .CK(clknet_leaf_133_clk),
    .Q(net9),
    .QN(_06965_));
 DFF_X2 \read_data1[14]$_SDFFCE_PN0P_  (.D(_00334_),
    .CK(clknet_leaf_123_clk),
    .Q(net10),
    .QN(_06964_));
 DFF_X2 \read_data1[15]$_SDFFCE_PN0P_  (.D(_00335_),
    .CK(clknet_leaf_123_clk),
    .Q(net11),
    .QN(_06963_));
 DFF_X2 \read_data1[16]$_SDFFCE_PN0P_  (.D(_00336_),
    .CK(clknet_leaf_122_clk),
    .Q(net12),
    .QN(_06962_));
 DFF_X2 \read_data1[17]$_SDFFCE_PN0P_  (.D(_00337_),
    .CK(clknet_leaf_134_clk),
    .Q(net13),
    .QN(_06961_));
 DFF_X2 \read_data1[18]$_SDFFCE_PN0P_  (.D(_00338_),
    .CK(clknet_leaf_100_clk),
    .Q(net14),
    .QN(_06960_));
 DFF_X2 \read_data1[19]$_SDFFCE_PN0P_  (.D(_00339_),
    .CK(clknet_leaf_100_clk),
    .Q(net15),
    .QN(_06959_));
 DFF_X1 \read_data1[1]$_SDFFCE_PN0P_  (.D(_00340_),
    .CK(clknet_leaf_99_clk),
    .Q(net16),
    .QN(_06958_));
 DFF_X1 \read_data1[20]$_SDFFCE_PN0P_  (.D(_00341_),
    .CK(clknet_leaf_99_clk),
    .Q(net17),
    .QN(_06957_));
 DFF_X1 \read_data1[21]$_SDFFCE_PN0P_  (.D(_00342_),
    .CK(clknet_leaf_99_clk),
    .Q(net18),
    .QN(_06956_));
 DFF_X1 \read_data1[22]$_SDFFCE_PN0P_  (.D(_00343_),
    .CK(clknet_leaf_95_clk),
    .Q(net19),
    .QN(_06955_));
 DFF_X1 \read_data1[23]$_SDFFCE_PN0P_  (.D(_00344_),
    .CK(clknet_leaf_95_clk),
    .Q(net20),
    .QN(_06954_));
 DFF_X1 \read_data1[24]$_SDFFCE_PN0P_  (.D(_00345_),
    .CK(clknet_leaf_93_clk),
    .Q(net21),
    .QN(_06953_));
 DFF_X1 \read_data1[25]$_SDFFCE_PN0P_  (.D(_00346_),
    .CK(clknet_leaf_93_clk),
    .Q(net22),
    .QN(_06952_));
 DFF_X1 \read_data1[26]$_SDFFCE_PN0P_  (.D(_00347_),
    .CK(clknet_leaf_93_clk),
    .Q(net23),
    .QN(_06951_));
 DFF_X1 \read_data1[27]$_SDFFCE_PN0P_  (.D(_00348_),
    .CK(clknet_leaf_93_clk),
    .Q(net24),
    .QN(_06950_));
 DFF_X2 \read_data1[28]$_SDFFCE_PN0P_  (.D(_00349_),
    .CK(clknet_leaf_60_clk),
    .Q(net25),
    .QN(_06949_));
 DFF_X1 \read_data1[29]$_SDFFCE_PN0P_  (.D(_00350_),
    .CK(clknet_leaf_60_clk),
    .Q(net26),
    .QN(_06948_));
 DFF_X1 \read_data1[2]$_SDFFCE_PN0P_  (.D(_00351_),
    .CK(clknet_leaf_67_clk),
    .Q(net27),
    .QN(_06947_));
 DFF_X2 \read_data1[30]$_SDFFCE_PN0P_  (.D(_00352_),
    .CK(clknet_leaf_60_clk),
    .Q(net28),
    .QN(_06946_));
 DFF_X1 \read_data1[31]$_SDFFCE_PN0P_  (.D(_00353_),
    .CK(clknet_leaf_67_clk),
    .Q(net29),
    .QN(_06945_));
 DFF_X2 \read_data1[3]$_SDFFCE_PN0P_  (.D(_00354_),
    .CK(clknet_leaf_70_clk),
    .Q(net30),
    .QN(_06944_));
 DFF_X1 \read_data1[4]$_SDFFCE_PN0P_  (.D(_00355_),
    .CK(clknet_leaf_70_clk),
    .Q(net31),
    .QN(_06943_));
 DFF_X1 \read_data1[5]$_SDFFCE_PN0P_  (.D(_00356_),
    .CK(clknet_leaf_61_clk),
    .Q(net32),
    .QN(_06942_));
 DFF_X2 \read_data1[6]$_SDFFCE_PN0P_  (.D(_00357_),
    .CK(clknet_leaf_60_clk),
    .Q(net33),
    .QN(_06941_));
 DFF_X2 \read_data1[7]$_SDFFCE_PN0P_  (.D(_00358_),
    .CK(clknet_leaf_59_clk),
    .Q(net34),
    .QN(_06940_));
 DFF_X1 \read_data1[8]$_SDFFCE_PN0P_  (.D(_00359_),
    .CK(clknet_leaf_95_clk),
    .Q(net35),
    .QN(_06939_));
 DFF_X2 \read_data1[9]$_SDFFCE_PN0P_  (.D(_00360_),
    .CK(clknet_leaf_100_clk),
    .Q(net36),
    .QN(_06938_));
 DFF_X1 \read_data2[0]$_SDFFCE_PN0P_  (.D(_00361_),
    .CK(clknet_leaf_101_clk),
    .Q(net37),
    .QN(_06937_));
 DFF_X2 \read_data2[10]$_SDFFCE_PN0P_  (.D(_00362_),
    .CK(clknet_leaf_123_clk),
    .Q(net38),
    .QN(_06936_));
 DFF_X2 \read_data2[11]$_SDFFCE_PN0P_  (.D(_00363_),
    .CK(clknet_leaf_120_clk),
    .Q(net39),
    .QN(_06935_));
 DFF_X2 \read_data2[12]$_SDFFCE_PN0P_  (.D(_00364_),
    .CK(clknet_leaf_120_clk),
    .Q(net40),
    .QN(_06934_));
 DFF_X2 \read_data2[13]$_SDFFCE_PN0P_  (.D(_00365_),
    .CK(clknet_leaf_112_clk),
    .Q(net41),
    .QN(_06933_));
 DFF_X2 \read_data2[14]$_SDFFCE_PN0P_  (.D(_00366_),
    .CK(clknet_leaf_123_clk),
    .Q(net42),
    .QN(_06932_));
 DFF_X2 \read_data2[15]$_SDFFCE_PN0P_  (.D(_00367_),
    .CK(clknet_leaf_121_clk),
    .Q(net43),
    .QN(_06931_));
 DFF_X2 \read_data2[16]$_SDFFCE_PN0P_  (.D(_00368_),
    .CK(clknet_leaf_122_clk),
    .Q(net44),
    .QN(_06930_));
 DFF_X1 \read_data2[17]$_SDFFCE_PN0P_  (.D(_00369_),
    .CK(clknet_leaf_102_clk),
    .Q(net45),
    .QN(_06929_));
 DFF_X1 \read_data2[18]$_SDFFCE_PN0P_  (.D(_00370_),
    .CK(clknet_leaf_102_clk),
    .Q(net46),
    .QN(_06928_));
 DFF_X1 \read_data2[19]$_SDFFCE_PN0P_  (.D(_00371_),
    .CK(clknet_leaf_104_clk),
    .Q(net47),
    .QN(_06927_));
 DFF_X1 \read_data2[1]$_SDFFCE_PN0P_  (.D(_00372_),
    .CK(clknet_leaf_104_clk),
    .Q(net48),
    .QN(_06926_));
 DFF_X1 \read_data2[20]$_SDFFCE_PN0P_  (.D(_00373_),
    .CK(clknet_leaf_104_clk),
    .Q(net49),
    .QN(_06925_));
 DFF_X1 \read_data2[21]$_SDFFCE_PN0P_  (.D(_00374_),
    .CK(clknet_leaf_104_clk),
    .Q(net50),
    .QN(_06924_));
 DFF_X1 \read_data2[22]$_SDFFCE_PN0P_  (.D(_00375_),
    .CK(clknet_leaf_89_clk),
    .Q(net51),
    .QN(_06923_));
 DFF_X1 \read_data2[23]$_SDFFCE_PN0P_  (.D(_00376_),
    .CK(clknet_leaf_90_clk),
    .Q(net52),
    .QN(_06922_));
 DFF_X1 \read_data2[24]$_SDFFCE_PN0P_  (.D(_00377_),
    .CK(clknet_leaf_90_clk),
    .Q(net53),
    .QN(_06921_));
 DFF_X1 \read_data2[25]$_SDFFCE_PN0P_  (.D(_00378_),
    .CK(clknet_leaf_90_clk),
    .Q(net54),
    .QN(_06920_));
 DFF_X2 \read_data2[26]$_SDFFCE_PN0P_  (.D(_00379_),
    .CK(clknet_leaf_91_clk),
    .Q(net55),
    .QN(_06919_));
 DFF_X1 \read_data2[27]$_SDFFCE_PN0P_  (.D(_00380_),
    .CK(clknet_leaf_91_clk),
    .Q(net56),
    .QN(_06918_));
 DFF_X2 \read_data2[28]$_SDFFCE_PN0P_  (.D(_00381_),
    .CK(clknet_leaf_81_clk),
    .Q(net57),
    .QN(_06917_));
 DFF_X2 \read_data2[29]$_SDFFCE_PN0P_  (.D(_00382_),
    .CK(clknet_leaf_70_clk),
    .Q(net58),
    .QN(_06916_));
 DFF_X2 \read_data2[2]$_SDFFCE_PN0P_  (.D(_00383_),
    .CK(clknet_leaf_71_clk),
    .Q(net59),
    .QN(_06915_));
 DFF_X2 \read_data2[30]$_SDFFCE_PN0P_  (.D(_00384_),
    .CK(clknet_leaf_71_clk),
    .Q(net60),
    .QN(_06914_));
 DFF_X2 \read_data2[31]$_SDFFCE_PN0P_  (.D(_00385_),
    .CK(clknet_leaf_70_clk),
    .Q(net61),
    .QN(_06913_));
 DFF_X2 \read_data2[3]$_SDFFCE_PN0P_  (.D(_00386_),
    .CK(clknet_leaf_71_clk),
    .Q(net62),
    .QN(_06912_));
 DFF_X2 \read_data2[4]$_SDFFCE_PN0P_  (.D(_00387_),
    .CK(clknet_leaf_71_clk),
    .Q(net63),
    .QN(_06911_));
 DFF_X2 \read_data2[5]$_SDFFCE_PN0P_  (.D(_00388_),
    .CK(clknet_leaf_71_clk),
    .Q(net64),
    .QN(_06910_));
 DFF_X2 \read_data2[6]$_SDFFCE_PN0P_  (.D(_00389_),
    .CK(clknet_leaf_92_clk),
    .Q(net65),
    .QN(_06909_));
 DFF_X2 \read_data2[7]$_SDFFCE_PN0P_  (.D(_00390_),
    .CK(clknet_leaf_92_clk),
    .Q(net66),
    .QN(_06908_));
 DFF_X2 \read_data2[8]$_SDFFCE_PN0P_  (.D(_00391_),
    .CK(clknet_leaf_103_clk),
    .Q(net67),
    .QN(_06907_));
 DFF_X1 \read_data2[9]$_SDFFCE_PN0P_  (.D(_00392_),
    .CK(clknet_leaf_102_clk),
    .Q(net68),
    .QN(_06906_));
 DFF_X1 \registers[0][0]$_SDFFCE_PN0P_  (.D(_00393_),
    .CK(clknet_leaf_131_clk),
    .Q(\registers[0][0] ),
    .QN(_06905_));
 DFF_X1 \registers[0][10]$_SDFFCE_PN0P_  (.D(_00394_),
    .CK(clknet_leaf_127_clk),
    .Q(\registers[0][10] ),
    .QN(_06904_));
 DFF_X1 \registers[0][11]$_SDFFCE_PN0P_  (.D(_00395_),
    .CK(clknet_leaf_127_clk),
    .Q(\registers[0][11] ),
    .QN(_06903_));
 DFF_X1 \registers[0][12]$_SDFFCE_PN0P_  (.D(_00396_),
    .CK(clknet_leaf_126_clk),
    .Q(\registers[0][12] ),
    .QN(_06902_));
 DFF_X1 \registers[0][13]$_SDFFCE_PN0P_  (.D(_00397_),
    .CK(clknet_leaf_132_clk),
    .Q(\registers[0][13] ),
    .QN(_06901_));
 DFF_X1 \registers[0][14]$_SDFFCE_PN0P_  (.D(_00398_),
    .CK(clknet_leaf_126_clk),
    .Q(\registers[0][14] ),
    .QN(_06900_));
 DFF_X1 \registers[0][15]$_SDFFCE_PN0P_  (.D(_00399_),
    .CK(clknet_leaf_129_clk),
    .Q(\registers[0][15] ),
    .QN(_06899_));
 DFF_X1 \registers[0][16]$_SDFFCE_PN0P_  (.D(_00400_),
    .CK(clknet_leaf_132_clk),
    .Q(\registers[0][16] ),
    .QN(_06898_));
 DFF_X1 \registers[0][17]$_SDFFCE_PN0P_  (.D(_00401_),
    .CK(clknet_leaf_135_clk),
    .Q(\registers[0][17] ),
    .QN(_06897_));
 DFF_X1 \registers[0][18]$_SDFFCE_PN0P_  (.D(_00402_),
    .CK(clknet_leaf_135_clk),
    .Q(\registers[0][18] ),
    .QN(_06896_));
 DFF_X1 \registers[0][19]$_SDFFCE_PN0P_  (.D(_00403_),
    .CK(clknet_leaf_97_clk),
    .Q(\registers[0][19] ),
    .QN(_06895_));
 DFF_X1 \registers[0][1]$_SDFFCE_PN0P_  (.D(_00404_),
    .CK(clknet_leaf_139_clk),
    .Q(\registers[0][1] ),
    .QN(_06894_));
 DFF_X1 \registers[0][20]$_SDFFCE_PN0P_  (.D(_00405_),
    .CK(clknet_leaf_97_clk),
    .Q(\registers[0][20] ),
    .QN(_06893_));
 DFF_X1 \registers[0][21]$_SDFFCE_PN0P_  (.D(_00406_),
    .CK(clknet_leaf_97_clk),
    .Q(\registers[0][21] ),
    .QN(_06892_));
 DFF_X1 \registers[0][22]$_SDFFCE_PN0P_  (.D(_00407_),
    .CK(clknet_leaf_96_clk),
    .Q(\registers[0][22] ),
    .QN(_06891_));
 DFF_X1 \registers[0][23]$_SDFFCE_PN0P_  (.D(_00408_),
    .CK(clknet_leaf_55_clk),
    .Q(\registers[0][23] ),
    .QN(_06890_));
 DFF_X1 \registers[0][24]$_SDFFCE_PN0P_  (.D(_00409_),
    .CK(clknet_leaf_55_clk),
    .Q(\registers[0][24] ),
    .QN(_06889_));
 DFF_X1 \registers[0][25]$_SDFFCE_PN0P_  (.D(_00410_),
    .CK(clknet_leaf_56_clk),
    .Q(\registers[0][25] ),
    .QN(_06888_));
 DFF_X1 \registers[0][26]$_SDFFCE_PN0P_  (.D(_00411_),
    .CK(clknet_leaf_57_clk),
    .Q(\registers[0][26] ),
    .QN(_06887_));
 DFF_X1 \registers[0][27]$_SDFFCE_PN0P_  (.D(_00412_),
    .CK(clknet_leaf_57_clk),
    .Q(\registers[0][27] ),
    .QN(_06886_));
 DFF_X1 \registers[0][28]$_SDFFCE_PN0P_  (.D(_00413_),
    .CK(clknet_leaf_65_clk),
    .Q(\registers[0][28] ),
    .QN(_06885_));
 DFF_X1 \registers[0][29]$_SDFFCE_PN0P_  (.D(_00414_),
    .CK(clknet_leaf_63_clk),
    .Q(\registers[0][29] ),
    .QN(_06884_));
 DFF_X1 \registers[0][2]$_SDFFCE_PN0P_  (.D(_00415_),
    .CK(clknet_leaf_65_clk),
    .Q(\registers[0][2] ),
    .QN(_06883_));
 DFF_X1 \registers[0][30]$_SDFFCE_PN0P_  (.D(_00416_),
    .CK(clknet_leaf_65_clk),
    .Q(\registers[0][30] ),
    .QN(_06882_));
 DFF_X1 \registers[0][31]$_SDFFCE_PN0P_  (.D(_00417_),
    .CK(clknet_leaf_65_clk),
    .Q(\registers[0][31] ),
    .QN(_06881_));
 DFF_X1 \registers[0][3]$_SDFFCE_PN0P_  (.D(_00418_),
    .CK(clknet_leaf_66_clk),
    .Q(\registers[0][3] ),
    .QN(_06880_));
 DFF_X1 \registers[0][4]$_SDFFCE_PN0P_  (.D(_00419_),
    .CK(clknet_leaf_62_clk),
    .Q(\registers[0][4] ),
    .QN(_06879_));
 DFF_X1 \registers[0][5]$_SDFFCE_PN0P_  (.D(_00420_),
    .CK(clknet_leaf_62_clk),
    .Q(\registers[0][5] ),
    .QN(_06878_));
 DFF_X1 \registers[0][6]$_SDFFCE_PN0P_  (.D(_00421_),
    .CK(clknet_leaf_58_clk),
    .Q(\registers[0][6] ),
    .QN(_06877_));
 DFF_X1 \registers[0][7]$_SDFFCE_PN0P_  (.D(_00422_),
    .CK(clknet_leaf_58_clk),
    .Q(\registers[0][7] ),
    .QN(_06876_));
 DFF_X1 \registers[0][8]$_SDFFCE_PN0P_  (.D(_00423_),
    .CK(clknet_leaf_136_clk),
    .Q(\registers[0][8] ),
    .QN(_06875_));
 DFF_X1 \registers[0][9]$_SDFFCE_PN0P_  (.D(_00424_),
    .CK(clknet_leaf_136_clk),
    .Q(\registers[0][9] ),
    .QN(_06874_));
 DFF_X1 \registers[10][0]$_SDFFCE_PN0P_  (.D(_00425_),
    .CK(clknet_leaf_12_clk),
    .Q(\registers[10][0] ),
    .QN(_06873_));
 DFF_X1 \registers[10][10]$_SDFFCE_PN0P_  (.D(_00426_),
    .CK(clknet_leaf_154_clk),
    .Q(\registers[10][10] ),
    .QN(_06872_));
 DFF_X1 \registers[10][11]$_SDFFCE_PN0P_  (.D(_00427_),
    .CK(clknet_leaf_156_clk),
    .Q(\registers[10][11] ),
    .QN(_06871_));
 DFF_X1 \registers[10][12]$_SDFFCE_PN0P_  (.D(_00428_),
    .CK(clknet_leaf_154_clk),
    .Q(\registers[10][12] ),
    .QN(_06870_));
 DFF_X1 \registers[10][13]$_SDFFCE_PN0P_  (.D(_00429_),
    .CK(clknet_leaf_0_clk),
    .Q(\registers[10][13] ),
    .QN(_06869_));
 DFF_X1 \registers[10][14]$_SDFFCE_PN0P_  (.D(_00430_),
    .CK(clknet_leaf_1_clk),
    .Q(\registers[10][14] ),
    .QN(_06868_));
 DFF_X1 \registers[10][15]$_SDFFCE_PN0P_  (.D(_00431_),
    .CK(clknet_leaf_158_clk),
    .Q(\registers[10][15] ),
    .QN(_06867_));
 DFF_X1 \registers[10][16]$_SDFFCE_PN0P_  (.D(_00432_),
    .CK(clknet_leaf_0_clk),
    .Q(\registers[10][16] ),
    .QN(_06866_));
 DFF_X1 \registers[10][17]$_SDFFCE_PN0P_  (.D(_00433_),
    .CK(clknet_leaf_4_clk),
    .Q(\registers[10][17] ),
    .QN(_06865_));
 DFF_X1 \registers[10][18]$_SDFFCE_PN0P_  (.D(_00434_),
    .CK(clknet_leaf_5_clk),
    .Q(\registers[10][18] ),
    .QN(_06864_));
 DFF_X1 \registers[10][19]$_SDFFCE_PN0P_  (.D(_00435_),
    .CK(clknet_leaf_6_clk),
    .Q(\registers[10][19] ),
    .QN(_06863_));
 DFF_X1 \registers[10][1]$_SDFFCE_PN0P_  (.D(_00436_),
    .CK(clknet_leaf_6_clk),
    .Q(\registers[10][1] ),
    .QN(_06862_));
 DFF_X1 \registers[10][20]$_SDFFCE_PN0P_  (.D(_00437_),
    .CK(clknet_leaf_6_clk),
    .Q(\registers[10][20] ),
    .QN(_06861_));
 DFF_X1 \registers[10][21]$_SDFFCE_PN0P_  (.D(_00438_),
    .CK(clknet_leaf_7_clk),
    .Q(\registers[10][21] ),
    .QN(_06860_));
 DFF_X1 \registers[10][22]$_SDFFCE_PN0P_  (.D(_00439_),
    .CK(clknet_leaf_26_clk),
    .Q(\registers[10][22] ),
    .QN(_06859_));
 DFF_X1 \registers[10][23]$_SDFFCE_PN0P_  (.D(_00440_),
    .CK(clknet_leaf_26_clk),
    .Q(\registers[10][23] ),
    .QN(_06858_));
 DFF_X1 \registers[10][24]$_SDFFCE_PN0P_  (.D(_00441_),
    .CK(clknet_leaf_27_clk),
    .Q(\registers[10][24] ),
    .QN(_06857_));
 DFF_X1 \registers[10][25]$_SDFFCE_PN0P_  (.D(_00442_),
    .CK(clknet_leaf_27_clk),
    .Q(\registers[10][25] ),
    .QN(_06856_));
 DFF_X1 \registers[10][26]$_SDFFCE_PN0P_  (.D(_00443_),
    .CK(clknet_leaf_28_clk),
    .Q(\registers[10][26] ),
    .QN(_06855_));
 DFF_X1 \registers[10][27]$_SDFFCE_PN0P_  (.D(_00444_),
    .CK(clknet_leaf_28_clk),
    .Q(\registers[10][27] ),
    .QN(_06854_));
 DFF_X1 \registers[10][28]$_SDFFCE_PN0P_  (.D(_00445_),
    .CK(clknet_leaf_35_clk),
    .Q(\registers[10][28] ),
    .QN(_06853_));
 DFF_X1 \registers[10][29]$_SDFFCE_PN0P_  (.D(_00446_),
    .CK(clknet_leaf_35_clk),
    .Q(\registers[10][29] ),
    .QN(_06852_));
 DFF_X1 \registers[10][2]$_SDFFCE_PN0P_  (.D(_00447_),
    .CK(clknet_leaf_35_clk),
    .Q(\registers[10][2] ),
    .QN(_06851_));
 DFF_X1 \registers[10][30]$_SDFFCE_PN0P_  (.D(_00448_),
    .CK(clknet_leaf_37_clk),
    .Q(\registers[10][30] ),
    .QN(_06850_));
 DFF_X1 \registers[10][31]$_SDFFCE_PN0P_  (.D(_00449_),
    .CK(clknet_leaf_36_clk),
    .Q(\registers[10][31] ),
    .QN(_06849_));
 DFF_X1 \registers[10][3]$_SDFFCE_PN0P_  (.D(_00450_),
    .CK(clknet_leaf_37_clk),
    .Q(\registers[10][3] ),
    .QN(_06848_));
 DFF_X1 \registers[10][4]$_SDFFCE_PN0P_  (.D(_00451_),
    .CK(clknet_leaf_35_clk),
    .Q(\registers[10][4] ),
    .QN(_06847_));
 DFF_X1 \registers[10][5]$_SDFFCE_PN0P_  (.D(_00452_),
    .CK(clknet_leaf_35_clk),
    .Q(\registers[10][5] ),
    .QN(_06846_));
 DFF_X1 \registers[10][6]$_SDFFCE_PN0P_  (.D(_00453_),
    .CK(clknet_leaf_29_clk),
    .Q(\registers[10][6] ),
    .QN(_06845_));
 DFF_X1 \registers[10][7]$_SDFFCE_PN0P_  (.D(_00454_),
    .CK(clknet_leaf_29_clk),
    .Q(\registers[10][7] ),
    .QN(_06844_));
 DFF_X1 \registers[10][8]$_SDFFCE_PN0P_  (.D(_00455_),
    .CK(clknet_leaf_11_clk),
    .Q(\registers[10][8] ),
    .QN(_06843_));
 DFF_X1 \registers[10][9]$_SDFFCE_PN0P_  (.D(_00456_),
    .CK(clknet_leaf_3_clk),
    .Q(\registers[10][9] ),
    .QN(_06842_));
 DFF_X1 \registers[11][0]$_SDFFCE_PN0P_  (.D(_00457_),
    .CK(clknet_leaf_2_clk),
    .Q(\registers[11][0] ),
    .QN(_06841_));
 DFF_X1 \registers[11][10]$_SDFFCE_PN0P_  (.D(_00458_),
    .CK(clknet_leaf_155_clk),
    .Q(\registers[11][10] ),
    .QN(_06840_));
 DFF_X1 \registers[11][11]$_SDFFCE_PN0P_  (.D(_00459_),
    .CK(clknet_leaf_156_clk),
    .Q(\registers[11][11] ),
    .QN(_06839_));
 DFF_X1 \registers[11][12]$_SDFFCE_PN0P_  (.D(_00460_),
    .CK(clknet_leaf_156_clk),
    .Q(\registers[11][12] ),
    .QN(_06838_));
 DFF_X1 \registers[11][13]$_SDFFCE_PN0P_  (.D(_00461_),
    .CK(clknet_leaf_4_clk),
    .Q(\registers[11][13] ),
    .QN(_06837_));
 DFF_X1 \registers[11][14]$_SDFFCE_PN0P_  (.D(_00462_),
    .CK(clknet_leaf_1_clk),
    .Q(\registers[11][14] ),
    .QN(_06836_));
 DFF_X1 \registers[11][15]$_SDFFCE_PN0P_  (.D(_00463_),
    .CK(clknet_leaf_159_clk),
    .Q(\registers[11][15] ),
    .QN(_06835_));
 DFF_X1 \registers[11][16]$_SDFFCE_PN0P_  (.D(_00464_),
    .CK(clknet_leaf_0_clk),
    .Q(\registers[11][16] ),
    .QN(_06834_));
 DFF_X1 \registers[11][17]$_SDFFCE_PN0P_  (.D(_00465_),
    .CK(clknet_leaf_4_clk),
    .Q(\registers[11][17] ),
    .QN(_06833_));
 DFF_X1 \registers[11][18]$_SDFFCE_PN0P_  (.D(_00466_),
    .CK(clknet_leaf_4_clk),
    .Q(\registers[11][18] ),
    .QN(_06832_));
 DFF_X1 \registers[11][19]$_SDFFCE_PN0P_  (.D(_00467_),
    .CK(clknet_leaf_6_clk),
    .Q(\registers[11][19] ),
    .QN(_06831_));
 DFF_X1 \registers[11][1]$_SDFFCE_PN0P_  (.D(_00468_),
    .CK(clknet_leaf_6_clk),
    .Q(\registers[11][1] ),
    .QN(_06830_));
 DFF_X1 \registers[11][20]$_SDFFCE_PN0P_  (.D(_00469_),
    .CK(clknet_leaf_7_clk),
    .Q(\registers[11][20] ),
    .QN(_06829_));
 DFF_X1 \registers[11][21]$_SDFFCE_PN0P_  (.D(_00470_),
    .CK(clknet_leaf_7_clk),
    .Q(\registers[11][21] ),
    .QN(_06828_));
 DFF_X1 \registers[11][22]$_SDFFCE_PN0P_  (.D(_00471_),
    .CK(clknet_leaf_26_clk),
    .Q(\registers[11][22] ),
    .QN(_06827_));
 DFF_X1 \registers[11][23]$_SDFFCE_PN0P_  (.D(_00472_),
    .CK(clknet_leaf_26_clk),
    .Q(\registers[11][23] ),
    .QN(_06826_));
 DFF_X1 \registers[11][24]$_SDFFCE_PN0P_  (.D(_00473_),
    .CK(clknet_leaf_27_clk),
    .Q(\registers[11][24] ),
    .QN(_06825_));
 DFF_X1 \registers[11][25]$_SDFFCE_PN0P_  (.D(_00474_),
    .CK(clknet_leaf_27_clk),
    .Q(\registers[11][25] ),
    .QN(_06824_));
 DFF_X1 \registers[11][26]$_SDFFCE_PN0P_  (.D(_00475_),
    .CK(clknet_leaf_29_clk),
    .Q(\registers[11][26] ),
    .QN(_06823_));
 DFF_X1 \registers[11][27]$_SDFFCE_PN0P_  (.D(_00476_),
    .CK(clknet_leaf_29_clk),
    .Q(\registers[11][27] ),
    .QN(_06822_));
 DFF_X1 \registers[11][28]$_SDFFCE_PN0P_  (.D(_00477_),
    .CK(clknet_leaf_30_clk),
    .Q(\registers[11][28] ),
    .QN(_06821_));
 DFF_X1 \registers[11][29]$_SDFFCE_PN0P_  (.D(_00478_),
    .CK(clknet_leaf_34_clk),
    .Q(\registers[11][29] ),
    .QN(_06820_));
 DFF_X1 \registers[11][2]$_SDFFCE_PN0P_  (.D(_00479_),
    .CK(clknet_leaf_37_clk),
    .Q(\registers[11][2] ),
    .QN(_06819_));
 DFF_X1 \registers[11][30]$_SDFFCE_PN0P_  (.D(_00480_),
    .CK(clknet_leaf_38_clk),
    .Q(\registers[11][30] ),
    .QN(_06818_));
 DFF_X1 \registers[11][31]$_SDFFCE_PN0P_  (.D(_00481_),
    .CK(clknet_leaf_38_clk),
    .Q(\registers[11][31] ),
    .QN(_06817_));
 DFF_X1 \registers[11][3]$_SDFFCE_PN0P_  (.D(_00482_),
    .CK(clknet_leaf_38_clk),
    .Q(\registers[11][3] ),
    .QN(_06816_));
 DFF_X1 \registers[11][4]$_SDFFCE_PN0P_  (.D(_00483_),
    .CK(clknet_leaf_38_clk),
    .Q(\registers[11][4] ),
    .QN(_06815_));
 DFF_X1 \registers[11][5]$_SDFFCE_PN0P_  (.D(_00484_),
    .CK(clknet_leaf_38_clk),
    .Q(\registers[11][5] ),
    .QN(_06814_));
 DFF_X1 \registers[11][6]$_SDFFCE_PN0P_  (.D(_00485_),
    .CK(clknet_leaf_30_clk),
    .Q(\registers[11][6] ),
    .QN(_06813_));
 DFF_X1 \registers[11][7]$_SDFFCE_PN0P_  (.D(_00486_),
    .CK(clknet_leaf_30_clk),
    .Q(\registers[11][7] ),
    .QN(_06812_));
 DFF_X1 \registers[11][8]$_SDFFCE_PN0P_  (.D(_00487_),
    .CK(clknet_leaf_3_clk),
    .Q(\registers[11][8] ),
    .QN(_06811_));
 DFF_X1 \registers[11][9]$_SDFFCE_PN0P_  (.D(_00488_),
    .CK(clknet_leaf_5_clk),
    .Q(\registers[11][9] ),
    .QN(_06810_));
 DFF_X1 \registers[12][0]$_SDFFCE_PN0P_  (.D(_00489_),
    .CK(clknet_leaf_2_clk),
    .Q(\registers[12][0] ),
    .QN(_06809_));
 DFF_X1 \registers[12][10]$_SDFFCE_PN0P_  (.D(_00490_),
    .CK(clknet_leaf_157_clk),
    .Q(\registers[12][10] ),
    .QN(_06808_));
 DFF_X1 \registers[12][11]$_SDFFCE_PN0P_  (.D(_00491_),
    .CK(clknet_leaf_156_clk),
    .Q(\registers[12][11] ),
    .QN(_06807_));
 DFF_X1 \registers[12][12]$_SDFFCE_PN0P_  (.D(_00492_),
    .CK(clknet_leaf_156_clk),
    .Q(\registers[12][12] ),
    .QN(_06806_));
 DFF_X1 \registers[12][13]$_SDFFCE_PN0P_  (.D(_00493_),
    .CK(clknet_leaf_2_clk),
    .Q(\registers[12][13] ),
    .QN(_06805_));
 DFF_X1 \registers[12][14]$_SDFFCE_PN0P_  (.D(_00494_),
    .CK(clknet_leaf_158_clk),
    .Q(\registers[12][14] ),
    .QN(_06804_));
 DFF_X1 \registers[12][15]$_SDFFCE_PN0P_  (.D(_00495_),
    .CK(clknet_leaf_158_clk),
    .Q(\registers[12][15] ),
    .QN(_06803_));
 DFF_X1 \registers[12][16]$_SDFFCE_PN0P_  (.D(_00496_),
    .CK(clknet_leaf_1_clk),
    .Q(\registers[12][16] ),
    .QN(_06802_));
 DFF_X1 \registers[12][17]$_SDFFCE_PN0P_  (.D(_00497_),
    .CK(clknet_leaf_4_clk),
    .Q(\registers[12][17] ),
    .QN(_06801_));
 DFF_X1 \registers[12][18]$_SDFFCE_PN0P_  (.D(_00498_),
    .CK(clknet_leaf_3_clk),
    .Q(\registers[12][18] ),
    .QN(_06800_));
 DFF_X1 \registers[12][19]$_SDFFCE_PN0P_  (.D(_00499_),
    .CK(clknet_leaf_8_clk),
    .Q(\registers[12][19] ),
    .QN(_06799_));
 DFF_X1 \registers[12][1]$_SDFFCE_PN0P_  (.D(_00500_),
    .CK(clknet_leaf_8_clk),
    .Q(\registers[12][1] ),
    .QN(_06798_));
 DFF_X1 \registers[12][20]$_SDFFCE_PN0P_  (.D(_00501_),
    .CK(clknet_leaf_8_clk),
    .Q(\registers[12][20] ),
    .QN(_06797_));
 DFF_X1 \registers[12][21]$_SDFFCE_PN0P_  (.D(_00502_),
    .CK(clknet_leaf_8_clk),
    .Q(\registers[12][21] ),
    .QN(_06796_));
 DFF_X1 \registers[12][22]$_SDFFCE_PN0P_  (.D(_00503_),
    .CK(clknet_leaf_25_clk),
    .Q(\registers[12][22] ),
    .QN(_06795_));
 DFF_X1 \registers[12][23]$_SDFFCE_PN0P_  (.D(_00504_),
    .CK(clknet_leaf_25_clk),
    .Q(\registers[12][23] ),
    .QN(_06794_));
 DFF_X1 \registers[12][24]$_SDFFCE_PN0P_  (.D(_00505_),
    .CK(clknet_leaf_28_clk),
    .Q(\registers[12][24] ),
    .QN(_06793_));
 DFF_X1 \registers[12][25]$_SDFFCE_PN0P_  (.D(_00506_),
    .CK(clknet_leaf_25_clk),
    .Q(\registers[12][25] ),
    .QN(_06792_));
 DFF_X1 \registers[12][26]$_SDFFCE_PN0P_  (.D(_00507_),
    .CK(clknet_leaf_28_clk),
    .Q(\registers[12][26] ),
    .QN(_06791_));
 DFF_X1 \registers[12][27]$_SDFFCE_PN0P_  (.D(_00508_),
    .CK(clknet_leaf_31_clk),
    .Q(\registers[12][27] ),
    .QN(_06790_));
 DFF_X1 \registers[12][28]$_SDFFCE_PN0P_  (.D(_00509_),
    .CK(clknet_leaf_34_clk),
    .Q(\registers[12][28] ),
    .QN(_06789_));
 DFF_X1 \registers[12][29]$_SDFFCE_PN0P_  (.D(_00510_),
    .CK(clknet_leaf_38_clk),
    .Q(\registers[12][29] ),
    .QN(_06788_));
 DFF_X1 \registers[12][2]$_SDFFCE_PN0P_  (.D(_00511_),
    .CK(clknet_leaf_39_clk),
    .Q(\registers[12][2] ),
    .QN(_06787_));
 DFF_X1 \registers[12][30]$_SDFFCE_PN0P_  (.D(_00512_),
    .CK(clknet_leaf_33_clk),
    .Q(\registers[12][30] ),
    .QN(_06786_));
 DFF_X1 \registers[12][31]$_SDFFCE_PN0P_  (.D(_00513_),
    .CK(clknet_leaf_40_clk),
    .Q(\registers[12][31] ),
    .QN(_06785_));
 DFF_X1 \registers[12][3]$_SDFFCE_PN0P_  (.D(_00514_),
    .CK(clknet_leaf_40_clk),
    .Q(\registers[12][3] ),
    .QN(_06784_));
 DFF_X1 \registers[12][4]$_SDFFCE_PN0P_  (.D(_00515_),
    .CK(clknet_leaf_39_clk),
    .Q(\registers[12][4] ),
    .QN(_06783_));
 DFF_X1 \registers[12][5]$_SDFFCE_PN0P_  (.D(_00516_),
    .CK(clknet_leaf_39_clk),
    .Q(\registers[12][5] ),
    .QN(_06782_));
 DFF_X1 \registers[12][6]$_SDFFCE_PN0P_  (.D(_00517_),
    .CK(clknet_leaf_32_clk),
    .Q(\registers[12][6] ),
    .QN(_06781_));
 DFF_X1 \registers[12][7]$_SDFFCE_PN0P_  (.D(_00518_),
    .CK(clknet_leaf_31_clk),
    .Q(\registers[12][7] ),
    .QN(_06780_));
 DFF_X1 \registers[12][8]$_SDFFCE_PN0P_  (.D(_00519_),
    .CK(clknet_leaf_11_clk),
    .Q(\registers[12][8] ),
    .QN(_06779_));
 DFF_X1 \registers[12][9]$_SDFFCE_PN0P_  (.D(_00520_),
    .CK(clknet_leaf_11_clk),
    .Q(\registers[12][9] ),
    .QN(_06778_));
 DFF_X1 \registers[13][0]$_SDFFCE_PN0P_  (.D(_00521_),
    .CK(clknet_leaf_155_clk),
    .Q(\registers[13][0] ),
    .QN(_06777_));
 DFF_X1 \registers[13][10]$_SDFFCE_PN0P_  (.D(_00522_),
    .CK(clknet_leaf_152_clk),
    .Q(\registers[13][10] ),
    .QN(_06776_));
 DFF_X1 \registers[13][11]$_SDFFCE_PN0P_  (.D(_00523_),
    .CK(clknet_leaf_157_clk),
    .Q(\registers[13][11] ),
    .QN(_06775_));
 DFF_X1 \registers[13][12]$_SDFFCE_PN0P_  (.D(_00524_),
    .CK(clknet_leaf_157_clk),
    .Q(\registers[13][12] ),
    .QN(_06774_));
 DFF_X1 \registers[13][13]$_SDFFCE_PN0P_  (.D(_00525_),
    .CK(clknet_leaf_2_clk),
    .Q(\registers[13][13] ),
    .QN(_06773_));
 DFF_X1 \registers[13][14]$_SDFFCE_PN0P_  (.D(_00526_),
    .CK(clknet_leaf_158_clk),
    .Q(\registers[13][14] ),
    .QN(_06772_));
 DFF_X1 \registers[13][15]$_SDFFCE_PN0P_  (.D(_00527_),
    .CK(clknet_leaf_156_clk),
    .Q(\registers[13][15] ),
    .QN(_06771_));
 DFF_X1 \registers[13][16]$_SDFFCE_PN0P_  (.D(_00528_),
    .CK(clknet_leaf_2_clk),
    .Q(\registers[13][16] ),
    .QN(_06770_));
 DFF_X1 \registers[13][17]$_SDFFCE_PN0P_  (.D(_00529_),
    .CK(clknet_leaf_2_clk),
    .Q(\registers[13][17] ),
    .QN(_06769_));
 DFF_X1 \registers[13][18]$_SDFFCE_PN0P_  (.D(_00530_),
    .CK(clknet_leaf_3_clk),
    .Q(\registers[13][18] ),
    .QN(_06768_));
 DFF_X1 \registers[13][19]$_SDFFCE_PN0P_  (.D(_00531_),
    .CK(clknet_leaf_9_clk),
    .Q(\registers[13][19] ),
    .QN(_06767_));
 DFF_X1 \registers[13][1]$_SDFFCE_PN0P_  (.D(_00532_),
    .CK(clknet_leaf_10_clk),
    .Q(\registers[13][1] ),
    .QN(_06766_));
 DFF_X1 \registers[13][20]$_SDFFCE_PN0P_  (.D(_00533_),
    .CK(clknet_leaf_9_clk),
    .Q(\registers[13][20] ),
    .QN(_06765_));
 DFF_X1 \registers[13][21]$_SDFFCE_PN0P_  (.D(_00534_),
    .CK(clknet_leaf_9_clk),
    .Q(\registers[13][21] ),
    .QN(_06764_));
 DFF_X1 \registers[13][22]$_SDFFCE_PN0P_  (.D(_00535_),
    .CK(clknet_leaf_24_clk),
    .Q(\registers[13][22] ),
    .QN(_06763_));
 DFF_X1 \registers[13][23]$_SDFFCE_PN0P_  (.D(_00536_),
    .CK(clknet_leaf_24_clk),
    .Q(\registers[13][23] ),
    .QN(_06762_));
 DFF_X1 \registers[13][24]$_SDFFCE_PN0P_  (.D(_00537_),
    .CK(clknet_leaf_23_clk),
    .Q(\registers[13][24] ),
    .QN(_06761_));
 DFF_X1 \registers[13][25]$_SDFFCE_PN0P_  (.D(_00538_),
    .CK(clknet_leaf_23_clk),
    .Q(\registers[13][25] ),
    .QN(_06760_));
 DFF_X1 \registers[13][26]$_SDFFCE_PN0P_  (.D(_00539_),
    .CK(clknet_leaf_31_clk),
    .Q(\registers[13][26] ),
    .QN(_06759_));
 DFF_X1 \registers[13][27]$_SDFFCE_PN0P_  (.D(_00540_),
    .CK(clknet_leaf_31_clk),
    .Q(\registers[13][27] ),
    .QN(_06758_));
 DFF_X1 \registers[13][28]$_SDFFCE_PN0P_  (.D(_00541_),
    .CK(clknet_leaf_31_clk),
    .Q(\registers[13][28] ),
    .QN(_06757_));
 DFF_X1 \registers[13][29]$_SDFFCE_PN0P_  (.D(_00542_),
    .CK(clknet_leaf_33_clk),
    .Q(\registers[13][29] ),
    .QN(_06756_));
 DFF_X1 \registers[13][2]$_SDFFCE_PN0P_  (.D(_00543_),
    .CK(clknet_leaf_40_clk),
    .Q(\registers[13][2] ),
    .QN(_06755_));
 DFF_X1 \registers[13][30]$_SDFFCE_PN0P_  (.D(_00544_),
    .CK(clknet_leaf_32_clk),
    .Q(\registers[13][30] ),
    .QN(_06754_));
 DFF_X1 \registers[13][31]$_SDFFCE_PN0P_  (.D(_00545_),
    .CK(clknet_leaf_40_clk),
    .Q(\registers[13][31] ),
    .QN(_06753_));
 DFF_X1 \registers[13][3]$_SDFFCE_PN0P_  (.D(_00546_),
    .CK(clknet_leaf_40_clk),
    .Q(\registers[13][3] ),
    .QN(_06752_));
 DFF_X1 \registers[13][4]$_SDFFCE_PN0P_  (.D(_00547_),
    .CK(clknet_leaf_32_clk),
    .Q(\registers[13][4] ),
    .QN(_06751_));
 DFF_X1 \registers[13][5]$_SDFFCE_PN0P_  (.D(_00548_),
    .CK(clknet_leaf_32_clk),
    .Q(\registers[13][5] ),
    .QN(_06750_));
 DFF_X1 \registers[13][6]$_SDFFCE_PN0P_  (.D(_00549_),
    .CK(clknet_leaf_32_clk),
    .Q(\registers[13][6] ),
    .QN(_06749_));
 DFF_X1 \registers[13][7]$_SDFFCE_PN0P_  (.D(_00550_),
    .CK(clknet_leaf_22_clk),
    .Q(\registers[13][7] ),
    .QN(_06748_));
 DFF_X1 \registers[13][8]$_SDFFCE_PN0P_  (.D(_00551_),
    .CK(clknet_leaf_11_clk),
    .Q(\registers[13][8] ),
    .QN(_06747_));
 DFF_X1 \registers[13][9]$_SDFFCE_PN0P_  (.D(_00552_),
    .CK(clknet_leaf_10_clk),
    .Q(\registers[13][9] ),
    .QN(_06746_));
 DFF_X1 \registers[14][0]$_SDFFCE_PN0P_  (.D(_00553_),
    .CK(clknet_leaf_155_clk),
    .Q(\registers[14][0] ),
    .QN(_06745_));
 DFF_X1 \registers[14][10]$_SDFFCE_PN0P_  (.D(_00554_),
    .CK(clknet_leaf_157_clk),
    .Q(\registers[14][10] ),
    .QN(_06744_));
 DFF_X1 \registers[14][11]$_SDFFCE_PN0P_  (.D(_00555_),
    .CK(clknet_leaf_156_clk),
    .Q(\registers[14][11] ),
    .QN(_06743_));
 DFF_X1 \registers[14][12]$_SDFFCE_PN0P_  (.D(_00556_),
    .CK(clknet_leaf_157_clk),
    .Q(\registers[14][12] ),
    .QN(_06742_));
 DFF_X1 \registers[14][13]$_SDFFCE_PN0P_  (.D(_00557_),
    .CK(clknet_leaf_1_clk),
    .Q(\registers[14][13] ),
    .QN(_06741_));
 DFF_X1 \registers[14][14]$_SDFFCE_PN0P_  (.D(_00558_),
    .CK(clknet_leaf_1_clk),
    .Q(\registers[14][14] ),
    .QN(_06740_));
 DFF_X1 \registers[14][15]$_SDFFCE_PN0P_  (.D(_00559_),
    .CK(clknet_leaf_156_clk),
    .Q(\registers[14][15] ),
    .QN(_06739_));
 DFF_X1 \registers[14][16]$_SDFFCE_PN0P_  (.D(_00560_),
    .CK(clknet_leaf_1_clk),
    .Q(\registers[14][16] ),
    .QN(_06738_));
 DFF_X1 \registers[14][17]$_SDFFCE_PN0P_  (.D(_00561_),
    .CK(clknet_leaf_3_clk),
    .Q(\registers[14][17] ),
    .QN(_06737_));
 DFF_X1 \registers[14][18]$_SDFFCE_PN0P_  (.D(_00562_),
    .CK(clknet_leaf_3_clk),
    .Q(\registers[14][18] ),
    .QN(_06736_));
 DFF_X1 \registers[14][19]$_SDFFCE_PN0P_  (.D(_00563_),
    .CK(clknet_leaf_8_clk),
    .Q(\registers[14][19] ),
    .QN(_06735_));
 DFF_X1 \registers[14][1]$_SDFFCE_PN0P_  (.D(_00564_),
    .CK(clknet_leaf_8_clk),
    .Q(\registers[14][1] ),
    .QN(_06734_));
 DFF_X1 \registers[14][20]$_SDFFCE_PN0P_  (.D(_00565_),
    .CK(clknet_leaf_8_clk),
    .Q(\registers[14][20] ),
    .QN(_06733_));
 DFF_X1 \registers[14][21]$_SDFFCE_PN0P_  (.D(_00566_),
    .CK(clknet_leaf_8_clk),
    .Q(\registers[14][21] ),
    .QN(_06732_));
 DFF_X1 \registers[14][22]$_SDFFCE_PN0P_  (.D(_00567_),
    .CK(clknet_leaf_25_clk),
    .Q(\registers[14][22] ),
    .QN(_06731_));
 DFF_X1 \registers[14][23]$_SDFFCE_PN0P_  (.D(_00568_),
    .CK(clknet_leaf_24_clk),
    .Q(\registers[14][23] ),
    .QN(_06730_));
 DFF_X1 \registers[14][24]$_SDFFCE_PN0P_  (.D(_00569_),
    .CK(clknet_leaf_25_clk),
    .Q(\registers[14][24] ),
    .QN(_06729_));
 DFF_X1 \registers[14][25]$_SDFFCE_PN0P_  (.D(_00570_),
    .CK(clknet_leaf_24_clk),
    .Q(\registers[14][25] ),
    .QN(_06728_));
 DFF_X1 \registers[14][26]$_SDFFCE_PN0P_  (.D(_00571_),
    .CK(clknet_leaf_30_clk),
    .Q(\registers[14][26] ),
    .QN(_06727_));
 DFF_X1 \registers[14][27]$_SDFFCE_PN0P_  (.D(_00572_),
    .CK(clknet_leaf_31_clk),
    .Q(\registers[14][27] ),
    .QN(_06726_));
 DFF_X1 \registers[14][28]$_SDFFCE_PN0P_  (.D(_00573_),
    .CK(clknet_leaf_34_clk),
    .Q(\registers[14][28] ),
    .QN(_06725_));
 DFF_X1 \registers[14][29]$_SDFFCE_PN0P_  (.D(_00574_),
    .CK(clknet_leaf_33_clk),
    .Q(\registers[14][29] ),
    .QN(_06724_));
 DFF_X1 \registers[14][2]$_SDFFCE_PN0P_  (.D(_00575_),
    .CK(clknet_leaf_33_clk),
    .Q(\registers[14][2] ),
    .QN(_06723_));
 DFF_X1 \registers[14][30]$_SDFFCE_PN0P_  (.D(_00576_),
    .CK(clknet_leaf_33_clk),
    .Q(\registers[14][30] ),
    .QN(_06722_));
 DFF_X1 \registers[14][31]$_SDFFCE_PN0P_  (.D(_00577_),
    .CK(clknet_leaf_39_clk),
    .Q(\registers[14][31] ),
    .QN(_06721_));
 DFF_X1 \registers[14][3]$_SDFFCE_PN0P_  (.D(_00578_),
    .CK(clknet_leaf_44_clk),
    .Q(\registers[14][3] ),
    .QN(_06720_));
 DFF_X1 \registers[14][4]$_SDFFCE_PN0P_  (.D(_00579_),
    .CK(clknet_leaf_39_clk),
    .Q(\registers[14][4] ),
    .QN(_06719_));
 DFF_X1 \registers[14][5]$_SDFFCE_PN0P_  (.D(_00580_),
    .CK(clknet_leaf_39_clk),
    .Q(\registers[14][5] ),
    .QN(_06718_));
 DFF_X1 \registers[14][6]$_SDFFCE_PN0P_  (.D(_00581_),
    .CK(clknet_leaf_40_clk),
    .Q(\registers[14][6] ),
    .QN(_06717_));
 DFF_X1 \registers[14][7]$_SDFFCE_PN0P_  (.D(_00582_),
    .CK(clknet_leaf_39_clk),
    .Q(\registers[14][7] ),
    .QN(_06716_));
 DFF_X1 \registers[14][8]$_SDFFCE_PN0P_  (.D(_00583_),
    .CK(clknet_leaf_11_clk),
    .Q(\registers[14][8] ),
    .QN(_06715_));
 DFF_X1 \registers[14][9]$_SDFFCE_PN0P_  (.D(_00584_),
    .CK(clknet_leaf_11_clk),
    .Q(\registers[14][9] ),
    .QN(_06714_));
 DFF_X1 \registers[15][0]$_SDFFCE_PN0P_  (.D(_00585_),
    .CK(clknet_leaf_144_clk),
    .Q(\registers[15][0] ),
    .QN(_06713_));
 DFF_X1 \registers[15][10]$_SDFFCE_PN0P_  (.D(_00586_),
    .CK(clknet_leaf_152_clk),
    .Q(\registers[15][10] ),
    .QN(_06712_));
 DFF_X1 \registers[15][11]$_SDFFCE_PN0P_  (.D(_00587_),
    .CK(clknet_leaf_152_clk),
    .Q(\registers[15][11] ),
    .QN(_06711_));
 DFF_X1 \registers[15][12]$_SDFFCE_PN0P_  (.D(_00588_),
    .CK(clknet_leaf_152_clk),
    .Q(\registers[15][12] ),
    .QN(_06710_));
 DFF_X1 \registers[15][13]$_SDFFCE_PN0P_  (.D(_00589_),
    .CK(clknet_leaf_144_clk),
    .Q(\registers[15][13] ),
    .QN(_06709_));
 DFF_X1 \registers[15][14]$_SDFFCE_PN0P_  (.D(_00590_),
    .CK(clknet_leaf_153_clk),
    .Q(\registers[15][14] ),
    .QN(_06708_));
 DFF_X1 \registers[15][15]$_SDFFCE_PN0P_  (.D(_00591_),
    .CK(clknet_leaf_153_clk),
    .Q(\registers[15][15] ),
    .QN(_06707_));
 DFF_X1 \registers[15][16]$_SDFFCE_PN0P_  (.D(_00592_),
    .CK(clknet_leaf_154_clk),
    .Q(\registers[15][16] ),
    .QN(_06706_));
 DFF_X1 \registers[15][17]$_SDFFCE_PN0P_  (.D(_00593_),
    .CK(clknet_leaf_12_clk),
    .Q(\registers[15][17] ),
    .QN(_06705_));
 DFF_X1 \registers[15][18]$_SDFFCE_PN0P_  (.D(_00594_),
    .CK(clknet_leaf_12_clk),
    .Q(\registers[15][18] ),
    .QN(_06704_));
 DFF_X1 \registers[15][19]$_SDFFCE_PN0P_  (.D(_00595_),
    .CK(clknet_leaf_10_clk),
    .Q(\registers[15][19] ),
    .QN(_06703_));
 DFF_X1 \registers[15][1]$_SDFFCE_PN0P_  (.D(_00596_),
    .CK(clknet_leaf_10_clk),
    .Q(\registers[15][1] ),
    .QN(_06702_));
 DFF_X1 \registers[15][20]$_SDFFCE_PN0P_  (.D(_00597_),
    .CK(clknet_leaf_9_clk),
    .Q(\registers[15][20] ),
    .QN(_06701_));
 DFF_X1 \registers[15][21]$_SDFFCE_PN0P_  (.D(_00598_),
    .CK(clknet_leaf_9_clk),
    .Q(\registers[15][21] ),
    .QN(_06700_));
 DFF_X1 \registers[15][22]$_SDFFCE_PN0P_  (.D(_00599_),
    .CK(clknet_leaf_24_clk),
    .Q(\registers[15][22] ),
    .QN(_06699_));
 DFF_X1 \registers[15][23]$_SDFFCE_PN0P_  (.D(_00600_),
    .CK(clknet_leaf_23_clk),
    .Q(\registers[15][23] ),
    .QN(_06698_));
 DFF_X1 \registers[15][24]$_SDFFCE_PN0P_  (.D(_00601_),
    .CK(clknet_leaf_23_clk),
    .Q(\registers[15][24] ),
    .QN(_06697_));
 DFF_X1 \registers[15][25]$_SDFFCE_PN0P_  (.D(_00602_),
    .CK(clknet_leaf_23_clk),
    .Q(\registers[15][25] ),
    .QN(_06696_));
 DFF_X1 \registers[15][26]$_SDFFCE_PN0P_  (.D(_00603_),
    .CK(clknet_leaf_22_clk),
    .Q(\registers[15][26] ),
    .QN(_06695_));
 DFF_X1 \registers[15][27]$_SDFFCE_PN0P_  (.D(_00604_),
    .CK(clknet_leaf_22_clk),
    .Q(\registers[15][27] ),
    .QN(_06694_));
 DFF_X1 \registers[15][28]$_SDFFCE_PN0P_  (.D(_00605_),
    .CK(clknet_leaf_32_clk),
    .Q(\registers[15][28] ),
    .QN(_06693_));
 DFF_X1 \registers[15][29]$_SDFFCE_PN0P_  (.D(_00606_),
    .CK(clknet_leaf_32_clk),
    .Q(\registers[15][29] ),
    .QN(_06692_));
 DFF_X1 \registers[15][2]$_SDFFCE_PN0P_  (.D(_00607_),
    .CK(clknet_leaf_41_clk),
    .Q(\registers[15][2] ),
    .QN(_06691_));
 DFF_X1 \registers[15][30]$_SDFFCE_PN0P_  (.D(_00608_),
    .CK(clknet_leaf_41_clk),
    .Q(\registers[15][30] ),
    .QN(_06690_));
 DFF_X1 \registers[15][31]$_SDFFCE_PN0P_  (.D(_00609_),
    .CK(clknet_leaf_41_clk),
    .Q(\registers[15][31] ),
    .QN(_06689_));
 DFF_X1 \registers[15][3]$_SDFFCE_PN0P_  (.D(_00610_),
    .CK(clknet_leaf_40_clk),
    .Q(\registers[15][3] ),
    .QN(_06688_));
 DFF_X1 \registers[15][4]$_SDFFCE_PN0P_  (.D(_00611_),
    .CK(clknet_leaf_41_clk),
    .Q(\registers[15][4] ),
    .QN(_06687_));
 DFF_X1 \registers[15][5]$_SDFFCE_PN0P_  (.D(_00612_),
    .CK(clknet_leaf_41_clk),
    .Q(\registers[15][5] ),
    .QN(_06686_));
 DFF_X1 \registers[15][6]$_SDFFCE_PN0P_  (.D(_00613_),
    .CK(clknet_leaf_32_clk),
    .Q(\registers[15][6] ),
    .QN(_06685_));
 DFF_X1 \registers[15][7]$_SDFFCE_PN0P_  (.D(_00614_),
    .CK(clknet_leaf_22_clk),
    .Q(\registers[15][7] ),
    .QN(_06684_));
 DFF_X1 \registers[15][8]$_SDFFCE_PN0P_  (.D(_00615_),
    .CK(clknet_leaf_12_clk),
    .Q(\registers[15][8] ),
    .QN(_06683_));
 DFF_X1 \registers[15][9]$_SDFFCE_PN0P_  (.D(_00616_),
    .CK(clknet_leaf_11_clk),
    .Q(\registers[15][9] ),
    .QN(_06682_));
 DFF_X1 \registers[16][0]$_SDFFCE_PN0P_  (.D(_00617_),
    .CK(clknet_leaf_112_clk),
    .Q(\registers[16][0] ),
    .QN(_06681_));
 DFF_X1 \registers[16][10]$_SDFFCE_PN0P_  (.D(_00618_),
    .CK(clknet_leaf_119_clk),
    .Q(\registers[16][10] ),
    .QN(_06680_));
 DFF_X1 \registers[16][11]$_SDFFCE_PN0P_  (.D(_00619_),
    .CK(clknet_leaf_118_clk),
    .Q(\registers[16][11] ),
    .QN(_06679_));
 DFF_X1 \registers[16][12]$_SDFFCE_PN0P_  (.D(_00620_),
    .CK(clknet_leaf_118_clk),
    .Q(\registers[16][12] ),
    .QN(_06678_));
 DFF_X1 \registers[16][13]$_SDFFCE_PN0P_  (.D(_00621_),
    .CK(clknet_leaf_118_clk),
    .Q(\registers[16][13] ),
    .QN(_06677_));
 DFF_X1 \registers[16][14]$_SDFFCE_PN0P_  (.D(_00622_),
    .CK(clknet_leaf_119_clk),
    .Q(\registers[16][14] ),
    .QN(_06676_));
 DFF_X1 \registers[16][15]$_SDFFCE_PN0P_  (.D(_00623_),
    .CK(clknet_leaf_120_clk),
    .Q(\registers[16][15] ),
    .QN(_06675_));
 DFF_X1 \registers[16][16]$_SDFFCE_PN0P_  (.D(_00624_),
    .CK(clknet_leaf_120_clk),
    .Q(\registers[16][16] ),
    .QN(_06674_));
 DFF_X1 \registers[16][17]$_SDFFCE_PN0P_  (.D(_00625_),
    .CK(clknet_leaf_111_clk),
    .Q(\registers[16][17] ),
    .QN(_06673_));
 DFF_X1 \registers[16][18]$_SDFFCE_PN0P_  (.D(_00626_),
    .CK(clknet_leaf_111_clk),
    .Q(\registers[16][18] ),
    .QN(_06672_));
 DFF_X1 \registers[16][19]$_SDFFCE_PN0P_  (.D(_00627_),
    .CK(clknet_leaf_106_clk),
    .Q(\registers[16][19] ),
    .QN(_06671_));
 DFF_X1 \registers[16][1]$_SDFFCE_PN0P_  (.D(_00628_),
    .CK(clknet_leaf_106_clk),
    .Q(\registers[16][1] ),
    .QN(_06670_));
 DFF_X1 \registers[16][20]$_SDFFCE_PN0P_  (.D(_00629_),
    .CK(clknet_leaf_106_clk),
    .Q(\registers[16][20] ),
    .QN(_06669_));
 DFF_X1 \registers[16][21]$_SDFFCE_PN0P_  (.D(_00630_),
    .CK(clknet_leaf_105_clk),
    .Q(\registers[16][21] ),
    .QN(_06668_));
 DFF_X1 \registers[16][22]$_SDFFCE_PN0P_  (.D(_00631_),
    .CK(clknet_leaf_88_clk),
    .Q(\registers[16][22] ),
    .QN(_06667_));
 DFF_X1 \registers[16][23]$_SDFFCE_PN0P_  (.D(_00632_),
    .CK(clknet_leaf_88_clk),
    .Q(\registers[16][23] ),
    .QN(_06666_));
 DFF_X1 \registers[16][24]$_SDFFCE_PN0P_  (.D(_00633_),
    .CK(clknet_leaf_88_clk),
    .Q(\registers[16][24] ),
    .QN(_06665_));
 DFF_X1 \registers[16][25]$_SDFFCE_PN0P_  (.D(_00634_),
    .CK(clknet_leaf_88_clk),
    .Q(\registers[16][25] ),
    .QN(_06664_));
 DFF_X1 \registers[16][26]$_SDFFCE_PN0P_  (.D(_00635_),
    .CK(clknet_leaf_82_clk),
    .Q(\registers[16][26] ),
    .QN(_06663_));
 DFF_X1 \registers[16][27]$_SDFFCE_PN0P_  (.D(_00636_),
    .CK(clknet_leaf_83_clk),
    .Q(\registers[16][27] ),
    .QN(_06662_));
 DFF_X1 \registers[16][28]$_SDFFCE_PN0P_  (.D(_00637_),
    .CK(clknet_leaf_72_clk),
    .Q(\registers[16][28] ),
    .QN(_06661_));
 DFF_X1 \registers[16][29]$_SDFFCE_PN0P_  (.D(_00638_),
    .CK(clknet_leaf_74_clk),
    .Q(\registers[16][29] ),
    .QN(_06660_));
 DFF_X1 \registers[16][2]$_SDFFCE_PN0P_  (.D(_00639_),
    .CK(clknet_leaf_74_clk),
    .Q(\registers[16][2] ),
    .QN(_06659_));
 DFF_X1 \registers[16][30]$_SDFFCE_PN0P_  (.D(_00640_),
    .CK(clknet_leaf_75_clk),
    .Q(\registers[16][30] ),
    .QN(_06658_));
 DFF_X1 \registers[16][31]$_SDFFCE_PN0P_  (.D(_00641_),
    .CK(clknet_leaf_75_clk),
    .Q(\registers[16][31] ),
    .QN(_06657_));
 DFF_X1 \registers[16][3]$_SDFFCE_PN0P_  (.D(_00642_),
    .CK(clknet_leaf_75_clk),
    .Q(\registers[16][3] ),
    .QN(_06656_));
 DFF_X1 \registers[16][4]$_SDFFCE_PN0P_  (.D(_00643_),
    .CK(clknet_leaf_72_clk),
    .Q(\registers[16][4] ),
    .QN(_06655_));
 DFF_X1 \registers[16][5]$_SDFFCE_PN0P_  (.D(_00644_),
    .CK(clknet_leaf_74_clk),
    .Q(\registers[16][5] ),
    .QN(_06654_));
 DFF_X1 \registers[16][6]$_SDFFCE_PN0P_  (.D(_00645_),
    .CK(clknet_leaf_82_clk),
    .Q(\registers[16][6] ),
    .QN(_06653_));
 DFF_X1 \registers[16][7]$_SDFFCE_PN0P_  (.D(_00646_),
    .CK(clknet_leaf_82_clk),
    .Q(\registers[16][7] ),
    .QN(_06652_));
 DFF_X1 \registers[16][8]$_SDFFCE_PN0P_  (.D(_00647_),
    .CK(clknet_leaf_112_clk),
    .Q(\registers[16][8] ),
    .QN(_06651_));
 DFF_X1 \registers[16][9]$_SDFFCE_PN0P_  (.D(_00648_),
    .CK(clknet_leaf_102_clk),
    .Q(\registers[16][9] ),
    .QN(_06650_));
 DFF_X1 \registers[17][0]$_SDFFCE_PN0P_  (.D(_00649_),
    .CK(clknet_leaf_112_clk),
    .Q(\registers[17][0] ),
    .QN(_06649_));
 DFF_X1 \registers[17][10]$_SDFFCE_PN0P_  (.D(_00650_),
    .CK(clknet_leaf_119_clk),
    .Q(\registers[17][10] ),
    .QN(_06648_));
 DFF_X1 \registers[17][11]$_SDFFCE_PN0P_  (.D(_00651_),
    .CK(clknet_leaf_118_clk),
    .Q(\registers[17][11] ),
    .QN(_06647_));
 DFF_X1 \registers[17][12]$_SDFFCE_PN0P_  (.D(_00652_),
    .CK(clknet_leaf_118_clk),
    .Q(\registers[17][12] ),
    .QN(_06646_));
 DFF_X1 \registers[17][13]$_SDFFCE_PN0P_  (.D(_00653_),
    .CK(clknet_leaf_118_clk),
    .Q(\registers[17][13] ),
    .QN(_06645_));
 DFF_X1 \registers[17][14]$_SDFFCE_PN0P_  (.D(_00654_),
    .CK(clknet_leaf_120_clk),
    .Q(\registers[17][14] ),
    .QN(_06644_));
 DFF_X1 \registers[17][15]$_SDFFCE_PN0P_  (.D(_00655_),
    .CK(clknet_leaf_120_clk),
    .Q(\registers[17][15] ),
    .QN(_06643_));
 DFF_X1 \registers[17][16]$_SDFFCE_PN0P_  (.D(_00656_),
    .CK(clknet_leaf_120_clk),
    .Q(\registers[17][16] ),
    .QN(_06642_));
 DFF_X1 \registers[17][17]$_SDFFCE_PN0P_  (.D(_00657_),
    .CK(clknet_leaf_111_clk),
    .Q(\registers[17][17] ),
    .QN(_06641_));
 DFF_X1 \registers[17][18]$_SDFFCE_PN0P_  (.D(_00658_),
    .CK(clknet_leaf_111_clk),
    .Q(\registers[17][18] ),
    .QN(_06640_));
 DFF_X1 \registers[17][19]$_SDFFCE_PN0P_  (.D(_00659_),
    .CK(clknet_leaf_103_clk),
    .Q(\registers[17][19] ),
    .QN(_06639_));
 DFF_X1 \registers[17][1]$_SDFFCE_PN0P_  (.D(_00660_),
    .CK(clknet_leaf_106_clk),
    .Q(\registers[17][1] ),
    .QN(_06638_));
 DFF_X1 \registers[17][20]$_SDFFCE_PN0P_  (.D(_00661_),
    .CK(clknet_leaf_105_clk),
    .Q(\registers[17][20] ),
    .QN(_06637_));
 DFF_X1 \registers[17][21]$_SDFFCE_PN0P_  (.D(_00662_),
    .CK(clknet_leaf_89_clk),
    .Q(\registers[17][21] ),
    .QN(_06636_));
 DFF_X1 \registers[17][22]$_SDFFCE_PN0P_  (.D(_00663_),
    .CK(clknet_leaf_87_clk),
    .Q(\registers[17][22] ),
    .QN(_06635_));
 DFF_X1 \registers[17][23]$_SDFFCE_PN0P_  (.D(_00664_),
    .CK(clknet_leaf_88_clk),
    .Q(\registers[17][23] ),
    .QN(_06634_));
 DFF_X1 \registers[17][24]$_SDFFCE_PN0P_  (.D(_00665_),
    .CK(clknet_leaf_88_clk),
    .Q(\registers[17][24] ),
    .QN(_06633_));
 DFF_X1 \registers[17][25]$_SDFFCE_PN0P_  (.D(_00666_),
    .CK(clknet_leaf_91_clk),
    .Q(\registers[17][25] ),
    .QN(_06632_));
 DFF_X1 \registers[17][26]$_SDFFCE_PN0P_  (.D(_00667_),
    .CK(clknet_leaf_82_clk),
    .Q(\registers[17][26] ),
    .QN(_06631_));
 DFF_X1 \registers[17][27]$_SDFFCE_PN0P_  (.D(_00668_),
    .CK(clknet_leaf_82_clk),
    .Q(\registers[17][27] ),
    .QN(_06630_));
 DFF_X1 \registers[17][28]$_SDFFCE_PN0P_  (.D(_00669_),
    .CK(clknet_leaf_75_clk),
    .Q(\registers[17][28] ),
    .QN(_06629_));
 DFF_X1 \registers[17][29]$_SDFFCE_PN0P_  (.D(_00670_),
    .CK(clknet_leaf_73_clk),
    .Q(\registers[17][29] ),
    .QN(_06628_));
 DFF_X1 \registers[17][2]$_SDFFCE_PN0P_  (.D(_00671_),
    .CK(clknet_leaf_74_clk),
    .Q(\registers[17][2] ),
    .QN(_06627_));
 DFF_X1 \registers[17][30]$_SDFFCE_PN0P_  (.D(_00672_),
    .CK(clknet_leaf_75_clk),
    .Q(\registers[17][30] ),
    .QN(_06626_));
 DFF_X1 \registers[17][31]$_SDFFCE_PN0P_  (.D(_00673_),
    .CK(clknet_leaf_75_clk),
    .Q(\registers[17][31] ),
    .QN(_06625_));
 DFF_X1 \registers[17][3]$_SDFFCE_PN0P_  (.D(_00674_),
    .CK(clknet_leaf_75_clk),
    .Q(\registers[17][3] ),
    .QN(_06624_));
 DFF_X1 \registers[17][4]$_SDFFCE_PN0P_  (.D(_00675_),
    .CK(clknet_leaf_80_clk),
    .Q(\registers[17][4] ),
    .QN(_06623_));
 DFF_X1 \registers[17][5]$_SDFFCE_PN0P_  (.D(_00676_),
    .CK(clknet_leaf_72_clk),
    .Q(\registers[17][5] ),
    .QN(_06622_));
 DFF_X1 \registers[17][6]$_SDFFCE_PN0P_  (.D(_00677_),
    .CK(clknet_leaf_80_clk),
    .Q(\registers[17][6] ),
    .QN(_06621_));
 DFF_X1 \registers[17][7]$_SDFFCE_PN0P_  (.D(_00678_),
    .CK(clknet_leaf_82_clk),
    .Q(\registers[17][7] ),
    .QN(_06620_));
 DFF_X1 \registers[17][8]$_SDFFCE_PN0P_  (.D(_00679_),
    .CK(clknet_leaf_111_clk),
    .Q(\registers[17][8] ),
    .QN(_06619_));
 DFF_X1 \registers[17][9]$_SDFFCE_PN0P_  (.D(_00680_),
    .CK(clknet_leaf_102_clk),
    .Q(\registers[17][9] ),
    .QN(_06618_));
 DFF_X1 \registers[18][0]$_SDFFCE_PN0P_  (.D(_00681_),
    .CK(clknet_leaf_114_clk),
    .Q(\registers[18][0] ),
    .QN(_06617_));
 DFF_X1 \registers[18][10]$_SDFFCE_PN0P_  (.D(_00682_),
    .CK(clknet_leaf_114_clk),
    .Q(\registers[18][10] ),
    .QN(_06616_));
 DFF_X1 \registers[18][11]$_SDFFCE_PN0P_  (.D(_00683_),
    .CK(clknet_leaf_117_clk),
    .Q(\registers[18][11] ),
    .QN(_06615_));
 DFF_X1 \registers[18][12]$_SDFFCE_PN0P_  (.D(_00684_),
    .CK(clknet_leaf_116_clk),
    .Q(\registers[18][12] ),
    .QN(_06614_));
 DFF_X1 \registers[18][13]$_SDFFCE_PN0P_  (.D(_00685_),
    .CK(clknet_leaf_115_clk),
    .Q(\registers[18][13] ),
    .QN(_06613_));
 DFF_X1 \registers[18][14]$_SDFFCE_PN0P_  (.D(_00686_),
    .CK(clknet_leaf_116_clk),
    .Q(\registers[18][14] ),
    .QN(_06612_));
 DFF_X1 \registers[18][15]$_SDFFCE_PN0P_  (.D(_00687_),
    .CK(clknet_leaf_115_clk),
    .Q(\registers[18][15] ),
    .QN(_06611_));
 DFF_X1 \registers[18][16]$_SDFFCE_PN0P_  (.D(_00688_),
    .CK(clknet_leaf_115_clk),
    .Q(\registers[18][16] ),
    .QN(_06610_));
 DFF_X1 \registers[18][17]$_SDFFCE_PN0P_  (.D(_00689_),
    .CK(clknet_leaf_109_clk),
    .Q(\registers[18][17] ),
    .QN(_06609_));
 DFF_X1 \registers[18][18]$_SDFFCE_PN0P_  (.D(_00690_),
    .CK(clknet_leaf_110_clk),
    .Q(\registers[18][18] ),
    .QN(_06608_));
 DFF_X1 \registers[18][19]$_SDFFCE_PN0P_  (.D(_00691_),
    .CK(clknet_leaf_108_clk),
    .Q(\registers[18][19] ),
    .QN(_06607_));
 DFF_X1 \registers[18][1]$_SDFFCE_PN0P_  (.D(_00692_),
    .CK(clknet_leaf_108_clk),
    .Q(\registers[18][1] ),
    .QN(_06606_));
 DFF_X1 \registers[18][20]$_SDFFCE_PN0P_  (.D(_00693_),
    .CK(clknet_leaf_107_clk),
    .Q(\registers[18][20] ),
    .QN(_06605_));
 DFF_X1 \registers[18][21]$_SDFFCE_PN0P_  (.D(_00694_),
    .CK(clknet_leaf_107_clk),
    .Q(\registers[18][21] ),
    .QN(_06604_));
 DFF_X1 \registers[18][22]$_SDFFCE_PN0P_  (.D(_00695_),
    .CK(clknet_leaf_87_clk),
    .Q(\registers[18][22] ),
    .QN(_06603_));
 DFF_X1 \registers[18][23]$_SDFFCE_PN0P_  (.D(_00696_),
    .CK(clknet_leaf_86_clk),
    .Q(\registers[18][23] ),
    .QN(_06602_));
 DFF_X1 \registers[18][24]$_SDFFCE_PN0P_  (.D(_00697_),
    .CK(clknet_leaf_86_clk),
    .Q(\registers[18][24] ),
    .QN(_06601_));
 DFF_X1 \registers[18][25]$_SDFFCE_PN0P_  (.D(_00698_),
    .CK(clknet_leaf_86_clk),
    .Q(\registers[18][25] ),
    .QN(_06600_));
 DFF_X1 \registers[18][26]$_SDFFCE_PN0P_  (.D(_00699_),
    .CK(clknet_leaf_84_clk),
    .Q(\registers[18][26] ),
    .QN(_06599_));
 DFF_X1 \registers[18][27]$_SDFFCE_PN0P_  (.D(_00700_),
    .CK(clknet_leaf_84_clk),
    .Q(\registers[18][27] ),
    .QN(_06598_));
 DFF_X1 \registers[18][28]$_SDFFCE_PN0P_  (.D(_00701_),
    .CK(clknet_leaf_79_clk),
    .Q(\registers[18][28] ),
    .QN(_06597_));
 DFF_X1 \registers[18][29]$_SDFFCE_PN0P_  (.D(_00702_),
    .CK(clknet_leaf_79_clk),
    .Q(\registers[18][29] ),
    .QN(_06596_));
 DFF_X1 \registers[18][2]$_SDFFCE_PN0P_  (.D(_00703_),
    .CK(clknet_leaf_78_clk),
    .Q(\registers[18][2] ),
    .QN(_06595_));
 DFF_X1 \registers[18][30]$_SDFFCE_PN0P_  (.D(_00704_),
    .CK(clknet_leaf_83_clk),
    .Q(\registers[18][30] ),
    .QN(_06594_));
 DFF_X1 \registers[18][31]$_SDFFCE_PN0P_  (.D(_00705_),
    .CK(clknet_leaf_78_clk),
    .Q(\registers[18][31] ),
    .QN(_06593_));
 DFF_X1 \registers[18][3]$_SDFFCE_PN0P_  (.D(_00706_),
    .CK(clknet_leaf_79_clk),
    .Q(\registers[18][3] ),
    .QN(_06592_));
 DFF_X1 \registers[18][4]$_SDFFCE_PN0P_  (.D(_00707_),
    .CK(clknet_leaf_78_clk),
    .Q(\registers[18][4] ),
    .QN(_06591_));
 DFF_X1 \registers[18][5]$_SDFFCE_PN0P_  (.D(_00708_),
    .CK(clknet_leaf_80_clk),
    .Q(\registers[18][5] ),
    .QN(_06590_));
 DFF_X1 \registers[18][6]$_SDFFCE_PN0P_  (.D(_00709_),
    .CK(clknet_leaf_84_clk),
    .Q(\registers[18][6] ),
    .QN(_06589_));
 DFF_X1 \registers[18][7]$_SDFFCE_PN0P_  (.D(_00710_),
    .CK(clknet_leaf_84_clk),
    .Q(\registers[18][7] ),
    .QN(_06588_));
 DFF_X1 \registers[18][8]$_SDFFCE_PN0P_  (.D(_00711_),
    .CK(clknet_leaf_110_clk),
    .Q(\registers[18][8] ),
    .QN(_06587_));
 DFF_X1 \registers[18][9]$_SDFFCE_PN0P_  (.D(_00712_),
    .CK(clknet_leaf_110_clk),
    .Q(\registers[18][9] ),
    .QN(_06586_));
 DFF_X1 \registers[19][0]$_SDFFCE_PN0P_  (.D(_00713_),
    .CK(clknet_leaf_114_clk),
    .Q(\registers[19][0] ),
    .QN(_06585_));
 DFF_X1 \registers[19][10]$_SDFFCE_PN0P_  (.D(_00714_),
    .CK(clknet_leaf_114_clk),
    .Q(\registers[19][10] ),
    .QN(_06584_));
 DFF_X1 \registers[19][11]$_SDFFCE_PN0P_  (.D(_00715_),
    .CK(clknet_leaf_115_clk),
    .Q(\registers[19][11] ),
    .QN(_06583_));
 DFF_X1 \registers[19][12]$_SDFFCE_PN0P_  (.D(_00716_),
    .CK(clknet_leaf_115_clk),
    .Q(\registers[19][12] ),
    .QN(_06582_));
 DFF_X1 \registers[19][13]$_SDFFCE_PN0P_  (.D(_00717_),
    .CK(clknet_leaf_115_clk),
    .Q(\registers[19][13] ),
    .QN(_06581_));
 DFF_X1 \registers[19][14]$_SDFFCE_PN0P_  (.D(_00718_),
    .CK(clknet_leaf_116_clk),
    .Q(\registers[19][14] ),
    .QN(_06580_));
 DFF_X1 \registers[19][15]$_SDFFCE_PN0P_  (.D(_00719_),
    .CK(clknet_leaf_116_clk),
    .Q(\registers[19][15] ),
    .QN(_06579_));
 DFF_X1 \registers[19][16]$_SDFFCE_PN0P_  (.D(_00720_),
    .CK(clknet_leaf_115_clk),
    .Q(\registers[19][16] ),
    .QN(_06578_));
 DFF_X1 \registers[19][17]$_SDFFCE_PN0P_  (.D(_00721_),
    .CK(clknet_leaf_109_clk),
    .Q(\registers[19][17] ),
    .QN(_06577_));
 DFF_X1 \registers[19][18]$_SDFFCE_PN0P_  (.D(_00722_),
    .CK(clknet_leaf_109_clk),
    .Q(\registers[19][18] ),
    .QN(_06576_));
 DFF_X1 \registers[19][19]$_SDFFCE_PN0P_  (.D(_00723_),
    .CK(clknet_leaf_108_clk),
    .Q(\registers[19][19] ),
    .QN(_06575_));
 DFF_X1 \registers[19][1]$_SDFFCE_PN0P_  (.D(_00724_),
    .CK(clknet_leaf_108_clk),
    .Q(\registers[19][1] ),
    .QN(_06574_));
 DFF_X1 \registers[19][20]$_SDFFCE_PN0P_  (.D(_00725_),
    .CK(clknet_leaf_107_clk),
    .Q(\registers[19][20] ),
    .QN(_06573_));
 DFF_X1 \registers[19][21]$_SDFFCE_PN0P_  (.D(_00726_),
    .CK(clknet_leaf_107_clk),
    .Q(\registers[19][21] ),
    .QN(_06572_));
 DFF_X1 \registers[19][22]$_SDFFCE_PN0P_  (.D(_00727_),
    .CK(clknet_leaf_87_clk),
    .Q(\registers[19][22] ),
    .QN(_06571_));
 DFF_X1 \registers[19][23]$_SDFFCE_PN0P_  (.D(_00728_),
    .CK(clknet_leaf_86_clk),
    .Q(\registers[19][23] ),
    .QN(_06570_));
 DFF_X1 \registers[19][24]$_SDFFCE_PN0P_  (.D(_00729_),
    .CK(clknet_leaf_86_clk),
    .Q(\registers[19][24] ),
    .QN(_06569_));
 DFF_X1 \registers[19][25]$_SDFFCE_PN0P_  (.D(_00730_),
    .CK(clknet_leaf_86_clk),
    .Q(\registers[19][25] ),
    .QN(_06568_));
 DFF_X1 \registers[19][26]$_SDFFCE_PN0P_  (.D(_00731_),
    .CK(clknet_leaf_84_clk),
    .Q(\registers[19][26] ),
    .QN(_06567_));
 DFF_X1 \registers[19][27]$_SDFFCE_PN0P_  (.D(_00732_),
    .CK(clknet_leaf_84_clk),
    .Q(\registers[19][27] ),
    .QN(_06566_));
 DFF_X1 \registers[19][28]$_SDFFCE_PN0P_  (.D(_00733_),
    .CK(clknet_leaf_79_clk),
    .Q(\registers[19][28] ),
    .QN(_06565_));
 DFF_X1 \registers[19][29]$_SDFFCE_PN0P_  (.D(_00734_),
    .CK(clknet_leaf_79_clk),
    .Q(\registers[19][29] ),
    .QN(_06564_));
 DFF_X1 \registers[19][2]$_SDFFCE_PN0P_  (.D(_00735_),
    .CK(clknet_leaf_77_clk),
    .Q(\registers[19][2] ),
    .QN(_06563_));
 DFF_X1 \registers[19][30]$_SDFFCE_PN0P_  (.D(_00736_),
    .CK(clknet_leaf_84_clk),
    .Q(\registers[19][30] ),
    .QN(_06562_));
 DFF_X1 \registers[19][31]$_SDFFCE_PN0P_  (.D(_00737_),
    .CK(clknet_leaf_77_clk),
    .Q(\registers[19][31] ),
    .QN(_06561_));
 DFF_X1 \registers[19][3]$_SDFFCE_PN0P_  (.D(_00738_),
    .CK(clknet_leaf_79_clk),
    .Q(\registers[19][3] ),
    .QN(_06560_));
 DFF_X1 \registers[19][4]$_SDFFCE_PN0P_  (.D(_00739_),
    .CK(clknet_leaf_78_clk),
    .Q(\registers[19][4] ),
    .QN(_06559_));
 DFF_X1 \registers[19][5]$_SDFFCE_PN0P_  (.D(_00740_),
    .CK(clknet_leaf_79_clk),
    .Q(\registers[19][5] ),
    .QN(_06558_));
 DFF_X1 \registers[19][6]$_SDFFCE_PN0P_  (.D(_00741_),
    .CK(clknet_leaf_83_clk),
    .Q(\registers[19][6] ),
    .QN(_06557_));
 DFF_X1 \registers[19][7]$_SDFFCE_PN0P_  (.D(_00742_),
    .CK(clknet_leaf_83_clk),
    .Q(\registers[19][7] ),
    .QN(_06556_));
 DFF_X1 \registers[19][8]$_SDFFCE_PN0P_  (.D(_00743_),
    .CK(clknet_leaf_110_clk),
    .Q(\registers[19][8] ),
    .QN(_06555_));
 DFF_X1 \registers[19][9]$_SDFFCE_PN0P_  (.D(_00744_),
    .CK(clknet_leaf_109_clk),
    .Q(\registers[19][9] ),
    .QN(_06554_));
 DFF_X1 \registers[1][0]$_SDFFCE_PN0P_  (.D(_00745_),
    .CK(clknet_leaf_132_clk),
    .Q(\registers[1][0] ),
    .QN(_06553_));
 DFF_X1 \registers[1][10]$_SDFFCE_PN0P_  (.D(_00746_),
    .CK(clknet_leaf_125_clk),
    .Q(\registers[1][10] ),
    .QN(_06552_));
 DFF_X1 \registers[1][11]$_SDFFCE_PN0P_  (.D(_00747_),
    .CK(clknet_leaf_125_clk),
    .Q(\registers[1][11] ),
    .QN(_06551_));
 DFF_X1 \registers[1][12]$_SDFFCE_PN0P_  (.D(_00748_),
    .CK(clknet_leaf_125_clk),
    .Q(\registers[1][12] ),
    .QN(_06550_));
 DFF_X1 \registers[1][13]$_SDFFCE_PN0P_  (.D(_00749_),
    .CK(clknet_leaf_127_clk),
    .Q(\registers[1][13] ),
    .QN(_06549_));
 DFF_X1 \registers[1][14]$_SDFFCE_PN0P_  (.D(_00750_),
    .CK(clknet_leaf_127_clk),
    .Q(\registers[1][14] ),
    .QN(_06548_));
 DFF_X1 \registers[1][15]$_SDFFCE_PN0P_  (.D(_00751_),
    .CK(clknet_leaf_129_clk),
    .Q(\registers[1][15] ),
    .QN(_06547_));
 DFF_X1 \registers[1][16]$_SDFFCE_PN0P_  (.D(_00752_),
    .CK(clknet_leaf_132_clk),
    .Q(\registers[1][16] ),
    .QN(_06546_));
 DFF_X1 \registers[1][17]$_SDFFCE_PN0P_  (.D(_00753_),
    .CK(clknet_leaf_135_clk),
    .Q(\registers[1][17] ),
    .QN(_06545_));
 DFF_X1 \registers[1][18]$_SDFFCE_PN0P_  (.D(_00754_),
    .CK(clknet_leaf_135_clk),
    .Q(\registers[1][18] ),
    .QN(_06544_));
 DFF_X1 \registers[1][19]$_SDFFCE_PN0P_  (.D(_00755_),
    .CK(clknet_leaf_98_clk),
    .Q(\registers[1][19] ),
    .QN(_06543_));
 DFF_X1 \registers[1][1]$_SDFFCE_PN0P_  (.D(_00756_),
    .CK(clknet_leaf_138_clk),
    .Q(\registers[1][1] ),
    .QN(_06542_));
 DFF_X1 \registers[1][20]$_SDFFCE_PN0P_  (.D(_00757_),
    .CK(clknet_leaf_98_clk),
    .Q(\registers[1][20] ),
    .QN(_06541_));
 DFF_X1 \registers[1][21]$_SDFFCE_PN0P_  (.D(_00758_),
    .CK(clknet_leaf_98_clk),
    .Q(\registers[1][21] ),
    .QN(_06540_));
 DFF_X1 \registers[1][22]$_SDFFCE_PN0P_  (.D(_00759_),
    .CK(clknet_leaf_96_clk),
    .Q(\registers[1][22] ),
    .QN(_06539_));
 DFF_X1 \registers[1][23]$_SDFFCE_PN0P_  (.D(_00760_),
    .CK(clknet_leaf_96_clk),
    .Q(\registers[1][23] ),
    .QN(_06538_));
 DFF_X1 \registers[1][24]$_SDFFCE_PN0P_  (.D(_00761_),
    .CK(clknet_leaf_96_clk),
    .Q(\registers[1][24] ),
    .QN(_06537_));
 DFF_X1 \registers[1][25]$_SDFFCE_PN0P_  (.D(_00762_),
    .CK(clknet_leaf_56_clk),
    .Q(\registers[1][25] ),
    .QN(_06536_));
 DFF_X1 \registers[1][26]$_SDFFCE_PN0P_  (.D(_00763_),
    .CK(clknet_leaf_59_clk),
    .Q(\registers[1][26] ),
    .QN(_06535_));
 DFF_X1 \registers[1][27]$_SDFFCE_PN0P_  (.D(_00764_),
    .CK(clknet_leaf_59_clk),
    .Q(\registers[1][27] ),
    .QN(_06534_));
 DFF_X1 \registers[1][28]$_SDFFCE_PN0P_  (.D(_00765_),
    .CK(clknet_leaf_66_clk),
    .Q(\registers[1][28] ),
    .QN(_06533_));
 DFF_X1 \registers[1][29]$_SDFFCE_PN0P_  (.D(_00766_),
    .CK(clknet_leaf_66_clk),
    .Q(\registers[1][29] ),
    .QN(_06532_));
 DFF_X1 \registers[1][2]$_SDFFCE_PN0P_  (.D(_00767_),
    .CK(clknet_leaf_66_clk),
    .Q(\registers[1][2] ),
    .QN(_06531_));
 DFF_X1 \registers[1][30]$_SDFFCE_PN0P_  (.D(_00768_),
    .CK(clknet_leaf_66_clk),
    .Q(\registers[1][30] ),
    .QN(_06530_));
 DFF_X1 \registers[1][31]$_SDFFCE_PN0P_  (.D(_00769_),
    .CK(clknet_leaf_66_clk),
    .Q(\registers[1][31] ),
    .QN(_06529_));
 DFF_X1 \registers[1][3]$_SDFFCE_PN0P_  (.D(_00770_),
    .CK(clknet_leaf_66_clk),
    .Q(\registers[1][3] ),
    .QN(_06528_));
 DFF_X1 \registers[1][4]$_SDFFCE_PN0P_  (.D(_00771_),
    .CK(clknet_leaf_61_clk),
    .Q(\registers[1][4] ),
    .QN(_06527_));
 DFF_X1 \registers[1][5]$_SDFFCE_PN0P_  (.D(_00772_),
    .CK(clknet_leaf_61_clk),
    .Q(\registers[1][5] ),
    .QN(_06526_));
 DFF_X1 \registers[1][6]$_SDFFCE_PN0P_  (.D(_00773_),
    .CK(clknet_leaf_59_clk),
    .Q(\registers[1][6] ),
    .QN(_06525_));
 DFF_X1 \registers[1][7]$_SDFFCE_PN0P_  (.D(_00774_),
    .CK(clknet_leaf_59_clk),
    .Q(\registers[1][7] ),
    .QN(_06524_));
 DFF_X1 \registers[1][8]$_SDFFCE_PN0P_  (.D(_00775_),
    .CK(clknet_leaf_135_clk),
    .Q(\registers[1][8] ),
    .QN(_06523_));
 DFF_X1 \registers[1][9]$_SDFFCE_PN0P_  (.D(_00776_),
    .CK(clknet_leaf_135_clk),
    .Q(\registers[1][9] ),
    .QN(_06522_));
 DFF_X1 \registers[20][0]$_SDFFCE_PN0P_  (.D(_00777_),
    .CK(clknet_leaf_112_clk),
    .Q(\registers[20][0] ),
    .QN(_06521_));
 DFF_X1 \registers[20][10]$_SDFFCE_PN0P_  (.D(_00778_),
    .CK(clknet_leaf_122_clk),
    .Q(\registers[20][10] ),
    .QN(_06520_));
 DFF_X1 \registers[20][11]$_SDFFCE_PN0P_  (.D(_00779_),
    .CK(clknet_leaf_113_clk),
    .Q(\registers[20][11] ),
    .QN(_06519_));
 DFF_X1 \registers[20][12]$_SDFFCE_PN0P_  (.D(_00780_),
    .CK(clknet_leaf_113_clk),
    .Q(\registers[20][12] ),
    .QN(_06518_));
 DFF_X1 \registers[20][13]$_SDFFCE_PN0P_  (.D(_00781_),
    .CK(clknet_leaf_122_clk),
    .Q(\registers[20][13] ),
    .QN(_06517_));
 DFF_X1 \registers[20][14]$_SDFFCE_PN0P_  (.D(_00782_),
    .CK(clknet_leaf_121_clk),
    .Q(\registers[20][14] ),
    .QN(_06516_));
 DFF_X1 \registers[20][15]$_SDFFCE_PN0P_  (.D(_00783_),
    .CK(clknet_leaf_121_clk),
    .Q(\registers[20][15] ),
    .QN(_06515_));
 DFF_X1 \registers[20][16]$_SDFFCE_PN0P_  (.D(_00784_),
    .CK(clknet_leaf_112_clk),
    .Q(\registers[20][16] ),
    .QN(_06514_));
 DFF_X1 \registers[20][17]$_SDFFCE_PN0P_  (.D(_00785_),
    .CK(clknet_leaf_102_clk),
    .Q(\registers[20][17] ),
    .QN(_06513_));
 DFF_X1 \registers[20][18]$_SDFFCE_PN0P_  (.D(_00786_),
    .CK(clknet_leaf_102_clk),
    .Q(\registers[20][18] ),
    .QN(_06512_));
 DFF_X1 \registers[20][19]$_SDFFCE_PN0P_  (.D(_00787_),
    .CK(clknet_leaf_103_clk),
    .Q(\registers[20][19] ),
    .QN(_06511_));
 DFF_X1 \registers[20][1]$_SDFFCE_PN0P_  (.D(_00788_),
    .CK(clknet_leaf_103_clk),
    .Q(\registers[20][1] ),
    .QN(_06510_));
 DFF_X1 \registers[20][20]$_SDFFCE_PN0P_  (.D(_00789_),
    .CK(clknet_leaf_105_clk),
    .Q(\registers[20][20] ),
    .QN(_06509_));
 DFF_X1 \registers[20][21]$_SDFFCE_PN0P_  (.D(_00790_),
    .CK(clknet_leaf_105_clk),
    .Q(\registers[20][21] ),
    .QN(_06508_));
 DFF_X1 \registers[20][22]$_SDFFCE_PN0P_  (.D(_00791_),
    .CK(clknet_leaf_105_clk),
    .Q(\registers[20][22] ),
    .QN(_06507_));
 DFF_X1 \registers[20][23]$_SDFFCE_PN0P_  (.D(_00792_),
    .CK(clknet_leaf_89_clk),
    .Q(\registers[20][23] ),
    .QN(_06506_));
 DFF_X1 \registers[20][24]$_SDFFCE_PN0P_  (.D(_00793_),
    .CK(clknet_leaf_90_clk),
    .Q(\registers[20][24] ),
    .QN(_06505_));
 DFF_X1 \registers[20][25]$_SDFFCE_PN0P_  (.D(_00794_),
    .CK(clknet_leaf_89_clk),
    .Q(\registers[20][25] ),
    .QN(_06504_));
 DFF_X1 \registers[20][26]$_SDFFCE_PN0P_  (.D(_00795_),
    .CK(clknet_leaf_91_clk),
    .Q(\registers[20][26] ),
    .QN(_06503_));
 DFF_X1 \registers[20][27]$_SDFFCE_PN0P_  (.D(_00796_),
    .CK(clknet_leaf_91_clk),
    .Q(\registers[20][27] ),
    .QN(_06502_));
 DFF_X1 \registers[20][28]$_SDFFCE_PN0P_  (.D(_00797_),
    .CK(clknet_leaf_81_clk),
    .Q(\registers[20][28] ),
    .QN(_06501_));
 DFF_X1 \registers[20][29]$_SDFFCE_PN0P_  (.D(_00798_),
    .CK(clknet_leaf_71_clk),
    .Q(\registers[20][29] ),
    .QN(_06500_));
 DFF_X1 \registers[20][2]$_SDFFCE_PN0P_  (.D(_00799_),
    .CK(clknet_leaf_73_clk),
    .Q(\registers[20][2] ),
    .QN(_06499_));
 DFF_X1 \registers[20][30]$_SDFFCE_PN0P_  (.D(_00800_),
    .CK(clknet_leaf_81_clk),
    .Q(\registers[20][30] ),
    .QN(_06498_));
 DFF_X1 \registers[20][31]$_SDFFCE_PN0P_  (.D(_00801_),
    .CK(clknet_leaf_73_clk),
    .Q(\registers[20][31] ),
    .QN(_06497_));
 DFF_X1 \registers[20][3]$_SDFFCE_PN0P_  (.D(_00802_),
    .CK(clknet_leaf_72_clk),
    .Q(\registers[20][3] ),
    .QN(_06496_));
 DFF_X1 \registers[20][4]$_SDFFCE_PN0P_  (.D(_00803_),
    .CK(clknet_leaf_73_clk),
    .Q(\registers[20][4] ),
    .QN(_06495_));
 DFF_X1 \registers[20][5]$_SDFFCE_PN0P_  (.D(_00804_),
    .CK(clknet_leaf_73_clk),
    .Q(\registers[20][5] ),
    .QN(_06494_));
 DFF_X1 \registers[20][6]$_SDFFCE_PN0P_  (.D(_00805_),
    .CK(clknet_leaf_92_clk),
    .Q(\registers[20][6] ),
    .QN(_06493_));
 DFF_X1 \registers[20][7]$_SDFFCE_PN0P_  (.D(_00806_),
    .CK(clknet_leaf_81_clk),
    .Q(\registers[20][7] ),
    .QN(_06492_));
 DFF_X1 \registers[20][8]$_SDFFCE_PN0P_  (.D(_00807_),
    .CK(clknet_leaf_112_clk),
    .Q(\registers[20][8] ),
    .QN(_06491_));
 DFF_X1 \registers[20][9]$_SDFFCE_PN0P_  (.D(_00808_),
    .CK(clknet_leaf_101_clk),
    .Q(\registers[20][9] ),
    .QN(_06490_));
 DFF_X1 \registers[21][0]$_SDFFCE_PN0P_  (.D(_00809_),
    .CK(clknet_leaf_122_clk),
    .Q(\registers[21][0] ),
    .QN(_06489_));
 DFF_X1 \registers[21][10]$_SDFFCE_PN0P_  (.D(_00810_),
    .CK(clknet_leaf_122_clk),
    .Q(\registers[21][10] ),
    .QN(_06488_));
 DFF_X1 \registers[21][11]$_SDFFCE_PN0P_  (.D(_00811_),
    .CK(clknet_leaf_113_clk),
    .Q(\registers[21][11] ),
    .QN(_06487_));
 DFF_X1 \registers[21][12]$_SDFFCE_PN0P_  (.D(_00812_),
    .CK(clknet_leaf_113_clk),
    .Q(\registers[21][12] ),
    .QN(_06486_));
 DFF_X1 \registers[21][13]$_SDFFCE_PN0P_  (.D(_00813_),
    .CK(clknet_leaf_121_clk),
    .Q(\registers[21][13] ),
    .QN(_06485_));
 DFF_X1 \registers[21][14]$_SDFFCE_PN0P_  (.D(_00814_),
    .CK(clknet_leaf_121_clk),
    .Q(\registers[21][14] ),
    .QN(_06484_));
 DFF_X1 \registers[21][15]$_SDFFCE_PN0P_  (.D(_00815_),
    .CK(clknet_leaf_121_clk),
    .Q(\registers[21][15] ),
    .QN(_06483_));
 DFF_X1 \registers[21][16]$_SDFFCE_PN0P_  (.D(_00816_),
    .CK(clknet_leaf_122_clk),
    .Q(\registers[21][16] ),
    .QN(_06482_));
 DFF_X1 \registers[21][17]$_SDFFCE_PN0P_  (.D(_00817_),
    .CK(clknet_leaf_102_clk),
    .Q(\registers[21][17] ),
    .QN(_06481_));
 DFF_X1 \registers[21][18]$_SDFFCE_PN0P_  (.D(_00818_),
    .CK(clknet_leaf_103_clk),
    .Q(\registers[21][18] ),
    .QN(_06480_));
 DFF_X1 \registers[21][19]$_SDFFCE_PN0P_  (.D(_00819_),
    .CK(clknet_leaf_103_clk),
    .Q(\registers[21][19] ),
    .QN(_06479_));
 DFF_X1 \registers[21][1]$_SDFFCE_PN0P_  (.D(_00820_),
    .CK(clknet_leaf_103_clk),
    .Q(\registers[21][1] ),
    .QN(_06478_));
 DFF_X1 \registers[21][20]$_SDFFCE_PN0P_  (.D(_00821_),
    .CK(clknet_leaf_105_clk),
    .Q(\registers[21][20] ),
    .QN(_06477_));
 DFF_X1 \registers[21][21]$_SDFFCE_PN0P_  (.D(_00822_),
    .CK(clknet_leaf_105_clk),
    .Q(\registers[21][21] ),
    .QN(_06476_));
 DFF_X1 \registers[21][22]$_SDFFCE_PN0P_  (.D(_00823_),
    .CK(clknet_leaf_89_clk),
    .Q(\registers[21][22] ),
    .QN(_06475_));
 DFF_X1 \registers[21][23]$_SDFFCE_PN0P_  (.D(_00824_),
    .CK(clknet_leaf_89_clk),
    .Q(\registers[21][23] ),
    .QN(_06474_));
 DFF_X1 \registers[21][24]$_SDFFCE_PN0P_  (.D(_00825_),
    .CK(clknet_leaf_90_clk),
    .Q(\registers[21][24] ),
    .QN(_06473_));
 DFF_X1 \registers[21][25]$_SDFFCE_PN0P_  (.D(_00826_),
    .CK(clknet_leaf_88_clk),
    .Q(\registers[21][25] ),
    .QN(_06472_));
 DFF_X1 \registers[21][26]$_SDFFCE_PN0P_  (.D(_00827_),
    .CK(clknet_leaf_91_clk),
    .Q(\registers[21][26] ),
    .QN(_06471_));
 DFF_X1 \registers[21][27]$_SDFFCE_PN0P_  (.D(_00828_),
    .CK(clknet_leaf_91_clk),
    .Q(\registers[21][27] ),
    .QN(_06470_));
 DFF_X1 \registers[21][28]$_SDFFCE_PN0P_  (.D(_00829_),
    .CK(clknet_leaf_81_clk),
    .Q(\registers[21][28] ),
    .QN(_06469_));
 DFF_X1 \registers[21][29]$_SDFFCE_PN0P_  (.D(_00830_),
    .CK(clknet_leaf_80_clk),
    .Q(\registers[21][29] ),
    .QN(_06468_));
 DFF_X1 \registers[21][2]$_SDFFCE_PN0P_  (.D(_00831_),
    .CK(clknet_leaf_73_clk),
    .Q(\registers[21][2] ),
    .QN(_06467_));
 DFF_X1 \registers[21][30]$_SDFFCE_PN0P_  (.D(_00832_),
    .CK(clknet_leaf_80_clk),
    .Q(\registers[21][30] ),
    .QN(_06466_));
 DFF_X1 \registers[21][31]$_SDFFCE_PN0P_  (.D(_00833_),
    .CK(clknet_leaf_72_clk),
    .Q(\registers[21][31] ),
    .QN(_06465_));
 DFF_X1 \registers[21][3]$_SDFFCE_PN0P_  (.D(_00834_),
    .CK(clknet_leaf_80_clk),
    .Q(\registers[21][3] ),
    .QN(_06464_));
 DFF_X1 \registers[21][4]$_SDFFCE_PN0P_  (.D(_00835_),
    .CK(clknet_leaf_72_clk),
    .Q(\registers[21][4] ),
    .QN(_06463_));
 DFF_X1 \registers[21][5]$_SDFFCE_PN0P_  (.D(_00836_),
    .CK(clknet_leaf_72_clk),
    .Q(\registers[21][5] ),
    .QN(_06462_));
 DFF_X1 \registers[21][6]$_SDFFCE_PN0P_  (.D(_00837_),
    .CK(clknet_leaf_81_clk),
    .Q(\registers[21][6] ),
    .QN(_06461_));
 DFF_X1 \registers[21][7]$_SDFFCE_PN0P_  (.D(_00838_),
    .CK(clknet_leaf_81_clk),
    .Q(\registers[21][7] ),
    .QN(_06460_));
 DFF_X1 \registers[21][8]$_SDFFCE_PN0P_  (.D(_00839_),
    .CK(clknet_leaf_113_clk),
    .Q(\registers[21][8] ),
    .QN(_06459_));
 DFF_X1 \registers[21][9]$_SDFFCE_PN0P_  (.D(_00840_),
    .CK(clknet_leaf_112_clk),
    .Q(\registers[21][9] ),
    .QN(_06458_));
 DFF_X1 \registers[22][0]$_SDFFCE_PN0P_  (.D(_00841_),
    .CK(clknet_leaf_114_clk),
    .Q(\registers[22][0] ),
    .QN(_06457_));
 DFF_X1 \registers[22][10]$_SDFFCE_PN0P_  (.D(_00842_),
    .CK(clknet_leaf_113_clk),
    .Q(\registers[22][10] ),
    .QN(_06456_));
 DFF_X1 \registers[22][11]$_SDFFCE_PN0P_  (.D(_00843_),
    .CK(clknet_leaf_117_clk),
    .Q(\registers[22][11] ),
    .QN(_06455_));
 DFF_X1 \registers[22][12]$_SDFFCE_PN0P_  (.D(_00844_),
    .CK(clknet_leaf_117_clk),
    .Q(\registers[22][12] ),
    .QN(_06454_));
 DFF_X1 \registers[22][13]$_SDFFCE_PN0P_  (.D(_00845_),
    .CK(clknet_leaf_118_clk),
    .Q(\registers[22][13] ),
    .QN(_06453_));
 DFF_X1 \registers[22][14]$_SDFFCE_PN0P_  (.D(_00846_),
    .CK(clknet_leaf_117_clk),
    .Q(\registers[22][14] ),
    .QN(_06452_));
 DFF_X1 \registers[22][15]$_SDFFCE_PN0P_  (.D(_00847_),
    .CK(clknet_leaf_118_clk),
    .Q(\registers[22][15] ),
    .QN(_06451_));
 DFF_X1 \registers[22][16]$_SDFFCE_PN0P_  (.D(_00848_),
    .CK(clknet_leaf_113_clk),
    .Q(\registers[22][16] ),
    .QN(_06450_));
 DFF_X1 \registers[22][17]$_SDFFCE_PN0P_  (.D(_00849_),
    .CK(clknet_leaf_111_clk),
    .Q(\registers[22][17] ),
    .QN(_06449_));
 DFF_X1 \registers[22][18]$_SDFFCE_PN0P_  (.D(_00850_),
    .CK(clknet_leaf_109_clk),
    .Q(\registers[22][18] ),
    .QN(_06448_));
 DFF_X1 \registers[22][19]$_SDFFCE_PN0P_  (.D(_00851_),
    .CK(clknet_leaf_108_clk),
    .Q(\registers[22][19] ),
    .QN(_06447_));
 DFF_X1 \registers[22][1]$_SDFFCE_PN0P_  (.D(_00852_),
    .CK(clknet_leaf_106_clk),
    .Q(\registers[22][1] ),
    .QN(_06446_));
 DFF_X1 \registers[22][20]$_SDFFCE_PN0P_  (.D(_00853_),
    .CK(clknet_leaf_107_clk),
    .Q(\registers[22][20] ),
    .QN(_06445_));
 DFF_X1 \registers[22][21]$_SDFFCE_PN0P_  (.D(_00854_),
    .CK(clknet_leaf_106_clk),
    .Q(\registers[22][21] ),
    .QN(_06444_));
 DFF_X1 \registers[22][22]$_SDFFCE_PN0P_  (.D(_00855_),
    .CK(clknet_leaf_87_clk),
    .Q(\registers[22][22] ),
    .QN(_06443_));
 DFF_X1 \registers[22][23]$_SDFFCE_PN0P_  (.D(_00856_),
    .CK(clknet_leaf_85_clk),
    .Q(\registers[22][23] ),
    .QN(_06442_));
 DFF_X1 \registers[22][24]$_SDFFCE_PN0P_  (.D(_00857_),
    .CK(clknet_leaf_85_clk),
    .Q(\registers[22][24] ),
    .QN(_06441_));
 DFF_X1 \registers[22][25]$_SDFFCE_PN0P_  (.D(_00858_),
    .CK(clknet_leaf_87_clk),
    .Q(\registers[22][25] ),
    .QN(_06440_));
 DFF_X1 \registers[22][26]$_SDFFCE_PN0P_  (.D(_00859_),
    .CK(clknet_leaf_83_clk),
    .Q(\registers[22][26] ),
    .QN(_06439_));
 DFF_X1 \registers[22][27]$_SDFFCE_PN0P_  (.D(_00860_),
    .CK(clknet_leaf_85_clk),
    .Q(\registers[22][27] ),
    .QN(_06438_));
 DFF_X1 \registers[22][28]$_SDFFCE_PN0P_  (.D(_00861_),
    .CK(clknet_leaf_76_clk),
    .Q(\registers[22][28] ),
    .QN(_06437_));
 DFF_X1 \registers[22][29]$_SDFFCE_PN0P_  (.D(_00862_),
    .CK(clknet_leaf_77_clk),
    .Q(\registers[22][29] ),
    .QN(_06436_));
 DFF_X1 \registers[22][2]$_SDFFCE_PN0P_  (.D(_00863_),
    .CK(clknet_leaf_76_clk),
    .Q(\registers[22][2] ),
    .QN(_06435_));
 DFF_X1 \registers[22][30]$_SDFFCE_PN0P_  (.D(_00864_),
    .CK(clknet_leaf_78_clk),
    .Q(\registers[22][30] ),
    .QN(_06434_));
 DFF_X1 \registers[22][31]$_SDFFCE_PN0P_  (.D(_00865_),
    .CK(clknet_leaf_76_clk),
    .Q(\registers[22][31] ),
    .QN(_06433_));
 DFF_X1 \registers[22][3]$_SDFFCE_PN0P_  (.D(_00866_),
    .CK(clknet_leaf_80_clk),
    .Q(\registers[22][3] ),
    .QN(_06432_));
 DFF_X1 \registers[22][4]$_SDFFCE_PN0P_  (.D(_00867_),
    .CK(clknet_leaf_76_clk),
    .Q(\registers[22][4] ),
    .QN(_06431_));
 DFF_X1 \registers[22][5]$_SDFFCE_PN0P_  (.D(_00868_),
    .CK(clknet_leaf_78_clk),
    .Q(\registers[22][5] ),
    .QN(_06430_));
 DFF_X1 \registers[22][6]$_SDFFCE_PN0P_  (.D(_00869_),
    .CK(clknet_leaf_83_clk),
    .Q(\registers[22][6] ),
    .QN(_06429_));
 DFF_X1 \registers[22][7]$_SDFFCE_PN0P_  (.D(_00870_),
    .CK(clknet_leaf_83_clk),
    .Q(\registers[22][7] ),
    .QN(_06428_));
 DFF_X1 \registers[22][8]$_SDFFCE_PN0P_  (.D(_00871_),
    .CK(clknet_leaf_111_clk),
    .Q(\registers[22][8] ),
    .QN(_06427_));
 DFF_X1 \registers[22][9]$_SDFFCE_PN0P_  (.D(_00872_),
    .CK(clknet_leaf_110_clk),
    .Q(\registers[22][9] ),
    .QN(_06426_));
 DFF_X1 \registers[23][0]$_SDFFCE_PN0P_  (.D(_00873_),
    .CK(clknet_leaf_114_clk),
    .Q(\registers[23][0] ),
    .QN(_06425_));
 DFF_X1 \registers[23][10]$_SDFFCE_PN0P_  (.D(_00874_),
    .CK(clknet_leaf_114_clk),
    .Q(\registers[23][10] ),
    .QN(_06424_));
 DFF_X1 \registers[23][11]$_SDFFCE_PN0P_  (.D(_00875_),
    .CK(clknet_leaf_116_clk),
    .Q(\registers[23][11] ),
    .QN(_06423_));
 DFF_X1 \registers[23][12]$_SDFFCE_PN0P_  (.D(_00876_),
    .CK(clknet_leaf_116_clk),
    .Q(\registers[23][12] ),
    .QN(_06422_));
 DFF_X1 \registers[23][13]$_SDFFCE_PN0P_  (.D(_00877_),
    .CK(clknet_leaf_117_clk),
    .Q(\registers[23][13] ),
    .QN(_06421_));
 DFF_X1 \registers[23][14]$_SDFFCE_PN0P_  (.D(_00878_),
    .CK(clknet_leaf_116_clk),
    .Q(\registers[23][14] ),
    .QN(_06420_));
 DFF_X1 \registers[23][15]$_SDFFCE_PN0P_  (.D(_00879_),
    .CK(clknet_leaf_117_clk),
    .Q(\registers[23][15] ),
    .QN(_06419_));
 DFF_X1 \registers[23][16]$_SDFFCE_PN0P_  (.D(_00880_),
    .CK(clknet_leaf_113_clk),
    .Q(\registers[23][16] ),
    .QN(_06418_));
 DFF_X1 \registers[23][17]$_SDFFCE_PN0P_  (.D(_00881_),
    .CK(clknet_leaf_109_clk),
    .Q(\registers[23][17] ),
    .QN(_06417_));
 DFF_X1 \registers[23][18]$_SDFFCE_PN0P_  (.D(_00882_),
    .CK(clknet_leaf_109_clk),
    .Q(\registers[23][18] ),
    .QN(_06416_));
 DFF_X1 \registers[23][19]$_SDFFCE_PN0P_  (.D(_00883_),
    .CK(clknet_leaf_108_clk),
    .Q(\registers[23][19] ),
    .QN(_06415_));
 DFF_X1 \registers[23][1]$_SDFFCE_PN0P_  (.D(_00884_),
    .CK(clknet_leaf_107_clk),
    .Q(\registers[23][1] ),
    .QN(_06414_));
 DFF_X1 \registers[23][20]$_SDFFCE_PN0P_  (.D(_00885_),
    .CK(clknet_leaf_107_clk),
    .Q(\registers[23][20] ),
    .QN(_06413_));
 DFF_X1 \registers[23][21]$_SDFFCE_PN0P_  (.D(_00886_),
    .CK(clknet_leaf_107_clk),
    .Q(\registers[23][21] ),
    .QN(_06412_));
 DFF_X1 \registers[23][22]$_SDFFCE_PN0P_  (.D(_00887_),
    .CK(clknet_leaf_87_clk),
    .Q(\registers[23][22] ),
    .QN(_06411_));
 DFF_X1 \registers[23][23]$_SDFFCE_PN0P_  (.D(_00888_),
    .CK(clknet_leaf_85_clk),
    .Q(\registers[23][23] ),
    .QN(_06410_));
 DFF_X1 \registers[23][24]$_SDFFCE_PN0P_  (.D(_00889_),
    .CK(clknet_leaf_85_clk),
    .Q(\registers[23][24] ),
    .QN(_06409_));
 DFF_X1 \registers[23][25]$_SDFFCE_PN0P_  (.D(_00890_),
    .CK(clknet_leaf_86_clk),
    .Q(\registers[23][25] ),
    .QN(_06408_));
 DFF_X1 \registers[23][26]$_SDFFCE_PN0P_  (.D(_00891_),
    .CK(clknet_leaf_85_clk),
    .Q(\registers[23][26] ),
    .QN(_06407_));
 DFF_X1 \registers[23][27]$_SDFFCE_PN0P_  (.D(_00892_),
    .CK(clknet_leaf_85_clk),
    .Q(\registers[23][27] ),
    .QN(_06406_));
 DFF_X1 \registers[23][28]$_SDFFCE_PN0P_  (.D(_00893_),
    .CK(clknet_leaf_76_clk),
    .Q(\registers[23][28] ),
    .QN(_06405_));
 DFF_X1 \registers[23][29]$_SDFFCE_PN0P_  (.D(_00894_),
    .CK(clknet_leaf_77_clk),
    .Q(\registers[23][29] ),
    .QN(_06404_));
 DFF_X1 \registers[23][2]$_SDFFCE_PN0P_  (.D(_00895_),
    .CK(clknet_leaf_77_clk),
    .Q(\registers[23][2] ),
    .QN(_06403_));
 DFF_X1 \registers[23][30]$_SDFFCE_PN0P_  (.D(_00896_),
    .CK(clknet_leaf_77_clk),
    .Q(\registers[23][30] ),
    .QN(_06402_));
 DFF_X1 \registers[23][31]$_SDFFCE_PN0P_  (.D(_00897_),
    .CK(clknet_leaf_76_clk),
    .Q(\registers[23][31] ),
    .QN(_06401_));
 DFF_X1 \registers[23][3]$_SDFFCE_PN0P_  (.D(_00898_),
    .CK(clknet_leaf_77_clk),
    .Q(\registers[23][3] ),
    .QN(_06400_));
 DFF_X1 \registers[23][4]$_SDFFCE_PN0P_  (.D(_00899_),
    .CK(clknet_leaf_76_clk),
    .Q(\registers[23][4] ),
    .QN(_06399_));
 DFF_X1 \registers[23][5]$_SDFFCE_PN0P_  (.D(_00900_),
    .CK(clknet_leaf_77_clk),
    .Q(\registers[23][5] ),
    .QN(_06398_));
 DFF_X1 \registers[23][6]$_SDFFCE_PN0P_  (.D(_00901_),
    .CK(clknet_leaf_78_clk),
    .Q(\registers[23][6] ),
    .QN(_06397_));
 DFF_X1 \registers[23][7]$_SDFFCE_PN0P_  (.D(_00902_),
    .CK(clknet_leaf_78_clk),
    .Q(\registers[23][7] ),
    .QN(_06396_));
 DFF_X1 \registers[23][8]$_SDFFCE_PN0P_  (.D(_00903_),
    .CK(clknet_leaf_110_clk),
    .Q(\registers[23][8] ),
    .QN(_06395_));
 DFF_X1 \registers[23][9]$_SDFFCE_PN0P_  (.D(_00904_),
    .CK(clknet_leaf_110_clk),
    .Q(\registers[23][9] ),
    .QN(_06394_));
 DFF_X1 \registers[24][0]$_SDFFCE_PN0P_  (.D(_00905_),
    .CK(clknet_leaf_146_clk),
    .Q(\registers[24][0] ),
    .QN(_06393_));
 DFF_X1 \registers[24][10]$_SDFFCE_PN0P_  (.D(_00906_),
    .CK(clknet_leaf_147_clk),
    .Q(\registers[24][10] ),
    .QN(_06392_));
 DFF_X1 \registers[24][11]$_SDFFCE_PN0P_  (.D(_00907_),
    .CK(clknet_leaf_147_clk),
    .Q(\registers[24][11] ),
    .QN(_06391_));
 DFF_X1 \registers[24][12]$_SDFFCE_PN0P_  (.D(_00908_),
    .CK(clknet_leaf_147_clk),
    .Q(\registers[24][12] ),
    .QN(_06390_));
 DFF_X1 \registers[24][13]$_SDFFCE_PN0P_  (.D(_00909_),
    .CK(clknet_leaf_145_clk),
    .Q(\registers[24][13] ),
    .QN(_06389_));
 DFF_X1 \registers[24][14]$_SDFFCE_PN0P_  (.D(_00910_),
    .CK(clknet_leaf_145_clk),
    .Q(\registers[24][14] ),
    .QN(_06388_));
 DFF_X1 \registers[24][15]$_SDFFCE_PN0P_  (.D(_00911_),
    .CK(clknet_leaf_145_clk),
    .Q(\registers[24][15] ),
    .QN(_06387_));
 DFF_X1 \registers[24][16]$_SDFFCE_PN0P_  (.D(_00912_),
    .CK(clknet_leaf_144_clk),
    .Q(\registers[24][16] ),
    .QN(_06386_));
 DFF_X1 \registers[24][17]$_SDFFCE_PN0P_  (.D(_00913_),
    .CK(clknet_leaf_143_clk),
    .Q(\registers[24][17] ),
    .QN(_06385_));
 DFF_X1 \registers[24][18]$_SDFFCE_PN0P_  (.D(_00914_),
    .CK(clknet_leaf_143_clk),
    .Q(\registers[24][18] ),
    .QN(_06384_));
 DFF_X1 \registers[24][19]$_SDFFCE_PN0P_  (.D(_00915_),
    .CK(clknet_leaf_140_clk),
    .Q(\registers[24][19] ),
    .QN(_06383_));
 DFF_X1 \registers[24][1]$_SDFFCE_PN0P_  (.D(_00916_),
    .CK(clknet_leaf_16_clk),
    .Q(\registers[24][1] ),
    .QN(_06382_));
 DFF_X1 \registers[24][20]$_SDFFCE_PN0P_  (.D(_00917_),
    .CK(clknet_leaf_17_clk),
    .Q(\registers[24][20] ),
    .QN(_06381_));
 DFF_X1 \registers[24][21]$_SDFFCE_PN0P_  (.D(_00918_),
    .CK(clknet_leaf_17_clk),
    .Q(\registers[24][21] ),
    .QN(_06380_));
 DFF_X1 \registers[24][22]$_SDFFCE_PN0P_  (.D(_00919_),
    .CK(clknet_leaf_15_clk),
    .Q(\registers[24][22] ),
    .QN(_06379_));
 DFF_X1 \registers[24][23]$_SDFFCE_PN0P_  (.D(_00920_),
    .CK(clknet_leaf_18_clk),
    .Q(\registers[24][23] ),
    .QN(_06378_));
 DFF_X1 \registers[24][24]$_SDFFCE_PN0P_  (.D(_00921_),
    .CK(clknet_leaf_18_clk),
    .Q(\registers[24][24] ),
    .QN(_06377_));
 DFF_X1 \registers[24][25]$_SDFFCE_PN0P_  (.D(_00922_),
    .CK(clknet_leaf_54_clk),
    .Q(\registers[24][25] ),
    .QN(_06376_));
 DFF_X1 \registers[24][26]$_SDFFCE_PN0P_  (.D(_00923_),
    .CK(clknet_leaf_52_clk),
    .Q(\registers[24][26] ),
    .QN(_06375_));
 DFF_X1 \registers[24][27]$_SDFFCE_PN0P_  (.D(_00924_),
    .CK(clknet_leaf_54_clk),
    .Q(\registers[24][27] ),
    .QN(_06374_));
 DFF_X1 \registers[24][28]$_SDFFCE_PN0P_  (.D(_00925_),
    .CK(clknet_leaf_45_clk),
    .Q(\registers[24][28] ),
    .QN(_06373_));
 DFF_X1 \registers[24][29]$_SDFFCE_PN0P_  (.D(_00926_),
    .CK(clknet_leaf_43_clk),
    .Q(\registers[24][29] ),
    .QN(_06372_));
 DFF_X1 \registers[24][2]$_SDFFCE_PN0P_  (.D(_00927_),
    .CK(clknet_leaf_44_clk),
    .Q(\registers[24][2] ),
    .QN(_06371_));
 DFF_X1 \registers[24][30]$_SDFFCE_PN0P_  (.D(_00928_),
    .CK(clknet_leaf_46_clk),
    .Q(\registers[24][30] ),
    .QN(_06370_));
 DFF_X1 \registers[24][31]$_SDFFCE_PN0P_  (.D(_00929_),
    .CK(clknet_leaf_45_clk),
    .Q(\registers[24][31] ),
    .QN(_06369_));
 DFF_X1 \registers[24][3]$_SDFFCE_PN0P_  (.D(_00930_),
    .CK(clknet_leaf_46_clk),
    .Q(\registers[24][3] ),
    .QN(_06368_));
 DFF_X1 \registers[24][4]$_SDFFCE_PN0P_  (.D(_00931_),
    .CK(clknet_leaf_45_clk),
    .Q(\registers[24][4] ),
    .QN(_06367_));
 DFF_X1 \registers[24][5]$_SDFFCE_PN0P_  (.D(_00932_),
    .CK(clknet_leaf_47_clk),
    .Q(\registers[24][5] ),
    .QN(_06366_));
 DFF_X1 \registers[24][6]$_SDFFCE_PN0P_  (.D(_00933_),
    .CK(clknet_leaf_47_clk),
    .Q(\registers[24][6] ),
    .QN(_06365_));
 DFF_X1 \registers[24][7]$_SDFFCE_PN0P_  (.D(_00934_),
    .CK(clknet_leaf_48_clk),
    .Q(\registers[24][7] ),
    .QN(_06364_));
 DFF_X1 \registers[24][8]$_SDFFCE_PN0P_  (.D(_00935_),
    .CK(clknet_leaf_141_clk),
    .Q(\registers[24][8] ),
    .QN(_06363_));
 DFF_X1 \registers[24][9]$_SDFFCE_PN0P_  (.D(_00936_),
    .CK(clknet_leaf_142_clk),
    .Q(\registers[24][9] ),
    .QN(_06362_));
 DFF_X1 \registers[25][0]$_SDFFCE_PN0P_  (.D(_00937_),
    .CK(clknet_leaf_146_clk),
    .Q(\registers[25][0] ),
    .QN(_06361_));
 DFF_X1 \registers[25][10]$_SDFFCE_PN0P_  (.D(_00938_),
    .CK(clknet_leaf_149_clk),
    .Q(\registers[25][10] ),
    .QN(_06360_));
 DFF_X1 \registers[25][11]$_SDFFCE_PN0P_  (.D(_00939_),
    .CK(clknet_leaf_148_clk),
    .Q(\registers[25][11] ),
    .QN(_06359_));
 DFF_X1 \registers[25][12]$_SDFFCE_PN0P_  (.D(_00940_),
    .CK(clknet_leaf_148_clk),
    .Q(\registers[25][12] ),
    .QN(_06358_));
 DFF_X1 \registers[25][13]$_SDFFCE_PN0P_  (.D(_00941_),
    .CK(clknet_leaf_150_clk),
    .Q(\registers[25][13] ),
    .QN(_06357_));
 DFF_X1 \registers[25][14]$_SDFFCE_PN0P_  (.D(_00942_),
    .CK(clknet_leaf_153_clk),
    .Q(\registers[25][14] ),
    .QN(_06356_));
 DFF_X1 \registers[25][15]$_SDFFCE_PN0P_  (.D(_00943_),
    .CK(clknet_leaf_148_clk),
    .Q(\registers[25][15] ),
    .QN(_06355_));
 DFF_X1 \registers[25][16]$_SDFFCE_PN0P_  (.D(_00944_),
    .CK(clknet_leaf_144_clk),
    .Q(\registers[25][16] ),
    .QN(_06354_));
 DFF_X1 \registers[25][17]$_SDFFCE_PN0P_  (.D(_00945_),
    .CK(clknet_leaf_13_clk),
    .Q(\registers[25][17] ),
    .QN(_06353_));
 DFF_X1 \registers[25][18]$_SDFFCE_PN0P_  (.D(_00946_),
    .CK(clknet_leaf_140_clk),
    .Q(\registers[25][18] ),
    .QN(_06352_));
 DFF_X1 \registers[25][19]$_SDFFCE_PN0P_  (.D(_00947_),
    .CK(clknet_leaf_140_clk),
    .Q(\registers[25][19] ),
    .QN(_06351_));
 DFF_X1 \registers[25][1]$_SDFFCE_PN0P_  (.D(_00948_),
    .CK(clknet_leaf_16_clk),
    .Q(\registers[25][1] ),
    .QN(_06350_));
 DFF_X1 \registers[25][20]$_SDFFCE_PN0P_  (.D(_00949_),
    .CK(clknet_leaf_16_clk),
    .Q(\registers[25][20] ),
    .QN(_06349_));
 DFF_X1 \registers[25][21]$_SDFFCE_PN0P_  (.D(_00950_),
    .CK(clknet_leaf_17_clk),
    .Q(\registers[25][21] ),
    .QN(_06348_));
 DFF_X1 \registers[25][22]$_SDFFCE_PN0P_  (.D(_00951_),
    .CK(clknet_leaf_19_clk),
    .Q(\registers[25][22] ),
    .QN(_06347_));
 DFF_X1 \registers[25][23]$_SDFFCE_PN0P_  (.D(_00952_),
    .CK(clknet_leaf_18_clk),
    .Q(\registers[25][23] ),
    .QN(_06346_));
 DFF_X1 \registers[25][24]$_SDFFCE_PN0P_  (.D(_00953_),
    .CK(clknet_leaf_18_clk),
    .Q(\registers[25][24] ),
    .QN(_06345_));
 DFF_X1 \registers[25][25]$_SDFFCE_PN0P_  (.D(_00954_),
    .CK(clknet_leaf_55_clk),
    .Q(\registers[25][25] ),
    .QN(_06344_));
 DFF_X1 \registers[25][26]$_SDFFCE_PN0P_  (.D(_00955_),
    .CK(clknet_leaf_52_clk),
    .Q(\registers[25][26] ),
    .QN(_06343_));
 DFF_X1 \registers[25][27]$_SDFFCE_PN0P_  (.D(_00956_),
    .CK(clknet_leaf_53_clk),
    .Q(\registers[25][27] ),
    .QN(_06342_));
 DFF_X1 \registers[25][28]$_SDFFCE_PN0P_  (.D(_00957_),
    .CK(clknet_leaf_44_clk),
    .Q(\registers[25][28] ),
    .QN(_06341_));
 DFF_X1 \registers[25][29]$_SDFFCE_PN0P_  (.D(_00958_),
    .CK(clknet_leaf_44_clk),
    .Q(\registers[25][29] ),
    .QN(_06340_));
 DFF_X1 \registers[25][2]$_SDFFCE_PN0P_  (.D(_00959_),
    .CK(clknet_leaf_44_clk),
    .Q(\registers[25][2] ),
    .QN(_06339_));
 DFF_X1 \registers[25][30]$_SDFFCE_PN0P_  (.D(_00960_),
    .CK(clknet_leaf_46_clk),
    .Q(\registers[25][30] ),
    .QN(_06338_));
 DFF_X1 \registers[25][31]$_SDFFCE_PN0P_  (.D(_00961_),
    .CK(clknet_leaf_45_clk),
    .Q(\registers[25][31] ),
    .QN(_06337_));
 DFF_X1 \registers[25][3]$_SDFFCE_PN0P_  (.D(_00962_),
    .CK(clknet_leaf_46_clk),
    .Q(\registers[25][3] ),
    .QN(_06336_));
 DFF_X1 \registers[25][4]$_SDFFCE_PN0P_  (.D(_00963_),
    .CK(clknet_leaf_45_clk),
    .Q(\registers[25][4] ),
    .QN(_06335_));
 DFF_X1 \registers[25][5]$_SDFFCE_PN0P_  (.D(_00964_),
    .CK(clknet_leaf_47_clk),
    .Q(\registers[25][5] ),
    .QN(_06334_));
 DFF_X1 \registers[25][6]$_SDFFCE_PN0P_  (.D(_00965_),
    .CK(clknet_leaf_49_clk),
    .Q(\registers[25][6] ),
    .QN(_06333_));
 DFF_X1 \registers[25][7]$_SDFFCE_PN0P_  (.D(_00966_),
    .CK(clknet_leaf_47_clk),
    .Q(\registers[25][7] ),
    .QN(_06332_));
 DFF_X1 \registers[25][8]$_SDFFCE_PN0P_  (.D(_00967_),
    .CK(clknet_leaf_141_clk),
    .Q(\registers[25][8] ),
    .QN(_06331_));
 DFF_X1 \registers[25][9]$_SDFFCE_PN0P_  (.D(_00968_),
    .CK(clknet_leaf_142_clk),
    .Q(\registers[25][9] ),
    .QN(_06330_));
 DFF_X1 \registers[26][0]$_SDFFCE_PN0P_  (.D(_00969_),
    .CK(clknet_leaf_146_clk),
    .Q(\registers[26][0] ),
    .QN(_06329_));
 DFF_X1 \registers[26][10]$_SDFFCE_PN0P_  (.D(_00970_),
    .CK(clknet_leaf_146_clk),
    .Q(\registers[26][10] ),
    .QN(_06328_));
 DFF_X1 \registers[26][11]$_SDFFCE_PN0P_  (.D(_00971_),
    .CK(clknet_leaf_147_clk),
    .Q(\registers[26][11] ),
    .QN(_06327_));
 DFF_X1 \registers[26][12]$_SDFFCE_PN0P_  (.D(_00972_),
    .CK(clknet_leaf_147_clk),
    .Q(\registers[26][12] ),
    .QN(_06326_));
 DFF_X1 \registers[26][13]$_SDFFCE_PN0P_  (.D(_00973_),
    .CK(clknet_leaf_145_clk),
    .Q(\registers[26][13] ),
    .QN(_06325_));
 DFF_X1 \registers[26][14]$_SDFFCE_PN0P_  (.D(_00974_),
    .CK(clknet_leaf_145_clk),
    .Q(\registers[26][14] ),
    .QN(_06324_));
 DFF_X1 \registers[26][15]$_SDFFCE_PN0P_  (.D(_00975_),
    .CK(clknet_leaf_145_clk),
    .Q(\registers[26][15] ),
    .QN(_06323_));
 DFF_X1 \registers[26][16]$_SDFFCE_PN0P_  (.D(_00976_),
    .CK(clknet_leaf_146_clk),
    .Q(\registers[26][16] ),
    .QN(_06322_));
 DFF_X1 \registers[26][17]$_SDFFCE_PN0P_  (.D(_00977_),
    .CK(clknet_leaf_142_clk),
    .Q(\registers[26][17] ),
    .QN(_06321_));
 DFF_X1 \registers[26][18]$_SDFFCE_PN0P_  (.D(_00978_),
    .CK(clknet_leaf_142_clk),
    .Q(\registers[26][18] ),
    .QN(_06320_));
 DFF_X1 \registers[26][19]$_SDFFCE_PN0P_  (.D(_00979_),
    .CK(clknet_leaf_140_clk),
    .Q(\registers[26][19] ),
    .QN(_06319_));
 DFF_X1 \registers[26][1]$_SDFFCE_PN0P_  (.D(_00980_),
    .CK(clknet_leaf_16_clk),
    .Q(\registers[26][1] ),
    .QN(_06318_));
 DFF_X1 \registers[26][20]$_SDFFCE_PN0P_  (.D(_00981_),
    .CK(clknet_leaf_139_clk),
    .Q(\registers[26][20] ),
    .QN(_06317_));
 DFF_X1 \registers[26][21]$_SDFFCE_PN0P_  (.D(_00982_),
    .CK(clknet_leaf_17_clk),
    .Q(\registers[26][21] ),
    .QN(_06316_));
 DFF_X1 \registers[26][22]$_SDFFCE_PN0P_  (.D(_00983_),
    .CK(clknet_leaf_17_clk),
    .Q(\registers[26][22] ),
    .QN(_06315_));
 DFF_X1 \registers[26][23]$_SDFFCE_PN0P_  (.D(_00984_),
    .CK(clknet_leaf_17_clk),
    .Q(\registers[26][23] ),
    .QN(_06314_));
 DFF_X1 \registers[26][24]$_SDFFCE_PN0P_  (.D(_00985_),
    .CK(clknet_leaf_54_clk),
    .Q(\registers[26][24] ),
    .QN(_06313_));
 DFF_X1 \registers[26][25]$_SDFFCE_PN0P_  (.D(_00986_),
    .CK(clknet_leaf_55_clk),
    .Q(\registers[26][25] ),
    .QN(_06312_));
 DFF_X1 \registers[26][26]$_SDFFCE_PN0P_  (.D(_00987_),
    .CK(clknet_leaf_52_clk),
    .Q(\registers[26][26] ),
    .QN(_06311_));
 DFF_X1 \registers[26][27]$_SDFFCE_PN0P_  (.D(_00988_),
    .CK(clknet_leaf_54_clk),
    .Q(\registers[26][27] ),
    .QN(_06310_));
 DFF_X1 \registers[26][28]$_SDFFCE_PN0P_  (.D(_00989_),
    .CK(clknet_leaf_44_clk),
    .Q(\registers[26][28] ),
    .QN(_06309_));
 DFF_X1 \registers[26][29]$_SDFFCE_PN0P_  (.D(_00990_),
    .CK(clknet_leaf_44_clk),
    .Q(\registers[26][29] ),
    .QN(_06308_));
 DFF_X1 \registers[26][2]$_SDFFCE_PN0P_  (.D(_00991_),
    .CK(clknet_leaf_44_clk),
    .Q(\registers[26][2] ),
    .QN(_06307_));
 DFF_X1 \registers[26][30]$_SDFFCE_PN0P_  (.D(_00992_),
    .CK(clknet_leaf_46_clk),
    .Q(\registers[26][30] ),
    .QN(_06306_));
 DFF_X1 \registers[26][31]$_SDFFCE_PN0P_  (.D(_00993_),
    .CK(clknet_leaf_46_clk),
    .Q(\registers[26][31] ),
    .QN(_06305_));
 DFF_X1 \registers[26][3]$_SDFFCE_PN0P_  (.D(_00994_),
    .CK(clknet_leaf_46_clk),
    .Q(\registers[26][3] ),
    .QN(_06304_));
 DFF_X1 \registers[26][4]$_SDFFCE_PN0P_  (.D(_00995_),
    .CK(clknet_leaf_47_clk),
    .Q(\registers[26][4] ),
    .QN(_06303_));
 DFF_X1 \registers[26][5]$_SDFFCE_PN0P_  (.D(_00996_),
    .CK(clknet_leaf_47_clk),
    .Q(\registers[26][5] ),
    .QN(_06302_));
 DFF_X1 \registers[26][6]$_SDFFCE_PN0P_  (.D(_00997_),
    .CK(clknet_leaf_47_clk),
    .Q(\registers[26][6] ),
    .QN(_06301_));
 DFF_X1 \registers[26][7]$_SDFFCE_PN0P_  (.D(_00998_),
    .CK(clknet_leaf_48_clk),
    .Q(\registers[26][7] ),
    .QN(_06300_));
 DFF_X1 \registers[26][8]$_SDFFCE_PN0P_  (.D(_00999_),
    .CK(clknet_leaf_141_clk),
    .Q(\registers[26][8] ),
    .QN(_06299_));
 DFF_X1 \registers[26][9]$_SDFFCE_PN0P_  (.D(_01000_),
    .CK(clknet_leaf_142_clk),
    .Q(\registers[26][9] ),
    .QN(_06298_));
 DFF_X1 \registers[27][0]$_SDFFCE_PN0P_  (.D(_01001_),
    .CK(clknet_leaf_131_clk),
    .Q(\registers[27][0] ),
    .QN(_06297_));
 DFF_X1 \registers[27][10]$_SDFFCE_PN0P_  (.D(_01002_),
    .CK(clknet_leaf_130_clk),
    .Q(\registers[27][10] ),
    .QN(_06296_));
 DFF_X1 \registers[27][11]$_SDFFCE_PN0P_  (.D(_01003_),
    .CK(clknet_leaf_128_clk),
    .Q(\registers[27][11] ),
    .QN(_06295_));
 DFF_X1 \registers[27][12]$_SDFFCE_PN0P_  (.D(_01004_),
    .CK(clknet_leaf_129_clk),
    .Q(\registers[27][12] ),
    .QN(_06294_));
 DFF_X1 \registers[27][13]$_SDFFCE_PN0P_  (.D(_01005_),
    .CK(clknet_leaf_148_clk),
    .Q(\registers[27][13] ),
    .QN(_06293_));
 DFF_X1 \registers[27][14]$_SDFFCE_PN0P_  (.D(_01006_),
    .CK(clknet_leaf_153_clk),
    .Q(\registers[27][14] ),
    .QN(_06292_));
 DFF_X1 \registers[27][15]$_SDFFCE_PN0P_  (.D(_01007_),
    .CK(clknet_leaf_148_clk),
    .Q(\registers[27][15] ),
    .QN(_06291_));
 DFF_X1 \registers[27][16]$_SDFFCE_PN0P_  (.D(_01008_),
    .CK(clknet_leaf_144_clk),
    .Q(\registers[27][16] ),
    .QN(_06290_));
 DFF_X1 \registers[27][17]$_SDFFCE_PN0P_  (.D(_01009_),
    .CK(clknet_leaf_13_clk),
    .Q(\registers[27][17] ),
    .QN(_06289_));
 DFF_X1 \registers[27][18]$_SDFFCE_PN0P_  (.D(_01010_),
    .CK(clknet_leaf_140_clk),
    .Q(\registers[27][18] ),
    .QN(_06288_));
 DFF_X1 \registers[27][19]$_SDFFCE_PN0P_  (.D(_01011_),
    .CK(clknet_leaf_140_clk),
    .Q(\registers[27][19] ),
    .QN(_06287_));
 DFF_X1 \registers[27][1]$_SDFFCE_PN0P_  (.D(_01012_),
    .CK(clknet_leaf_16_clk),
    .Q(\registers[27][1] ),
    .QN(_06286_));
 DFF_X1 \registers[27][20]$_SDFFCE_PN0P_  (.D(_01013_),
    .CK(clknet_leaf_15_clk),
    .Q(\registers[27][20] ),
    .QN(_06285_));
 DFF_X1 \registers[27][21]$_SDFFCE_PN0P_  (.D(_01014_),
    .CK(clknet_leaf_16_clk),
    .Q(\registers[27][21] ),
    .QN(_06284_));
 DFF_X1 \registers[27][22]$_SDFFCE_PN0P_  (.D(_01015_),
    .CK(clknet_leaf_19_clk),
    .Q(\registers[27][22] ),
    .QN(_06283_));
 DFF_X1 \registers[27][23]$_SDFFCE_PN0P_  (.D(_01016_),
    .CK(clknet_leaf_18_clk),
    .Q(\registers[27][23] ),
    .QN(_06282_));
 DFF_X1 \registers[27][24]$_SDFFCE_PN0P_  (.D(_01017_),
    .CK(clknet_leaf_18_clk),
    .Q(\registers[27][24] ),
    .QN(_06281_));
 DFF_X1 \registers[27][25]$_SDFFCE_PN0P_  (.D(_01018_),
    .CK(clknet_leaf_18_clk),
    .Q(\registers[27][25] ),
    .QN(_06280_));
 DFF_X1 \registers[27][26]$_SDFFCE_PN0P_  (.D(_01019_),
    .CK(clknet_leaf_52_clk),
    .Q(\registers[27][26] ),
    .QN(_06279_));
 DFF_X1 \registers[27][27]$_SDFFCE_PN0P_  (.D(_01020_),
    .CK(clknet_leaf_53_clk),
    .Q(\registers[27][27] ),
    .QN(_06278_));
 DFF_X1 \registers[27][28]$_SDFFCE_PN0P_  (.D(_01021_),
    .CK(clknet_leaf_45_clk),
    .Q(\registers[27][28] ),
    .QN(_06277_));
 DFF_X1 \registers[27][29]$_SDFFCE_PN0P_  (.D(_01022_),
    .CK(clknet_leaf_45_clk),
    .Q(\registers[27][29] ),
    .QN(_06276_));
 DFF_X1 \registers[27][2]$_SDFFCE_PN0P_  (.D(_01023_),
    .CK(clknet_leaf_43_clk),
    .Q(\registers[27][2] ),
    .QN(_06275_));
 DFF_X1 \registers[27][30]$_SDFFCE_PN0P_  (.D(_01024_),
    .CK(clknet_leaf_43_clk),
    .Q(\registers[27][30] ),
    .QN(_06274_));
 DFF_X1 \registers[27][31]$_SDFFCE_PN0P_  (.D(_01025_),
    .CK(clknet_leaf_43_clk),
    .Q(\registers[27][31] ),
    .QN(_06273_));
 DFF_X1 \registers[27][3]$_SDFFCE_PN0P_  (.D(_01026_),
    .CK(clknet_leaf_43_clk),
    .Q(\registers[27][3] ),
    .QN(_06272_));
 DFF_X1 \registers[27][4]$_SDFFCE_PN0P_  (.D(_01027_),
    .CK(clknet_leaf_43_clk),
    .Q(\registers[27][4] ),
    .QN(_06271_));
 DFF_X1 \registers[27][5]$_SDFFCE_PN0P_  (.D(_01028_),
    .CK(clknet_leaf_42_clk),
    .Q(\registers[27][5] ),
    .QN(_06270_));
 DFF_X1 \registers[27][6]$_SDFFCE_PN0P_  (.D(_01029_),
    .CK(clknet_leaf_49_clk),
    .Q(\registers[27][6] ),
    .QN(_06269_));
 DFF_X1 \registers[27][7]$_SDFFCE_PN0P_  (.D(_01030_),
    .CK(clknet_leaf_42_clk),
    .Q(\registers[27][7] ),
    .QN(_06268_));
 DFF_X1 \registers[27][8]$_SDFFCE_PN0P_  (.D(_01031_),
    .CK(clknet_leaf_142_clk),
    .Q(\registers[27][8] ),
    .QN(_06267_));
 DFF_X1 \registers[27][9]$_SDFFCE_PN0P_  (.D(_01032_),
    .CK(clknet_leaf_143_clk),
    .Q(\registers[27][9] ),
    .QN(_06266_));
 DFF_X1 \registers[28][0]$_SDFFCE_PN0P_  (.D(_01033_),
    .CK(clknet_leaf_146_clk),
    .Q(\registers[28][0] ),
    .QN(_06265_));
 DFF_X1 \registers[28][10]$_SDFFCE_PN0P_  (.D(_01034_),
    .CK(clknet_leaf_148_clk),
    .Q(\registers[28][10] ),
    .QN(_06264_));
 DFF_X1 \registers[28][11]$_SDFFCE_PN0P_  (.D(_01035_),
    .CK(clknet_leaf_150_clk),
    .Q(\registers[28][11] ),
    .QN(_06263_));
 DFF_X1 \registers[28][12]$_SDFFCE_PN0P_  (.D(_01036_),
    .CK(clknet_leaf_150_clk),
    .Q(\registers[28][12] ),
    .QN(_06262_));
 DFF_X1 \registers[28][13]$_SDFFCE_PN0P_  (.D(_01037_),
    .CK(clknet_leaf_151_clk),
    .Q(\registers[28][13] ),
    .QN(_06261_));
 DFF_X1 \registers[28][14]$_SDFFCE_PN0P_  (.D(_01038_),
    .CK(clknet_leaf_151_clk),
    .Q(\registers[28][14] ),
    .QN(_06260_));
 DFF_X1 \registers[28][15]$_SDFFCE_PN0P_  (.D(_01039_),
    .CK(clknet_leaf_150_clk),
    .Q(\registers[28][15] ),
    .QN(_06259_));
 DFF_X1 \registers[28][16]$_SDFFCE_PN0P_  (.D(_01040_),
    .CK(clknet_leaf_153_clk),
    .Q(\registers[28][16] ),
    .QN(_06258_));
 DFF_X1 \registers[28][17]$_SDFFCE_PN0P_  (.D(_01041_),
    .CK(clknet_leaf_12_clk),
    .Q(\registers[28][17] ),
    .QN(_06257_));
 DFF_X1 \registers[28][18]$_SDFFCE_PN0P_  (.D(_01042_),
    .CK(clknet_leaf_12_clk),
    .Q(\registers[28][18] ),
    .QN(_06256_));
 DFF_X1 \registers[28][19]$_SDFFCE_PN0P_  (.D(_01043_),
    .CK(clknet_leaf_10_clk),
    .Q(\registers[28][19] ),
    .QN(_06255_));
 DFF_X1 \registers[28][1]$_SDFFCE_PN0P_  (.D(_01044_),
    .CK(clknet_leaf_14_clk),
    .Q(\registers[28][1] ),
    .QN(_06254_));
 DFF_X1 \registers[28][20]$_SDFFCE_PN0P_  (.D(_01045_),
    .CK(clknet_leaf_14_clk),
    .Q(\registers[28][20] ),
    .QN(_06253_));
 DFF_X1 \registers[28][21]$_SDFFCE_PN0P_  (.D(_01046_),
    .CK(clknet_leaf_14_clk),
    .Q(\registers[28][21] ),
    .QN(_06252_));
 DFF_X1 \registers[28][22]$_SDFFCE_PN0P_  (.D(_01047_),
    .CK(clknet_leaf_19_clk),
    .Q(\registers[28][22] ),
    .QN(_06251_));
 DFF_X1 \registers[28][23]$_SDFFCE_PN0P_  (.D(_01048_),
    .CK(clknet_leaf_20_clk),
    .Q(\registers[28][23] ),
    .QN(_06250_));
 DFF_X1 \registers[28][24]$_SDFFCE_PN0P_  (.D(_01049_),
    .CK(clknet_leaf_20_clk),
    .Q(\registers[28][24] ),
    .QN(_06249_));
 DFF_X1 \registers[28][25]$_SDFFCE_PN0P_  (.D(_01050_),
    .CK(clknet_leaf_20_clk),
    .Q(\registers[28][25] ),
    .QN(_06248_));
 DFF_X1 \registers[28][26]$_SDFFCE_PN0P_  (.D(_01051_),
    .CK(clknet_leaf_21_clk),
    .Q(\registers[28][26] ),
    .QN(_06247_));
 DFF_X1 \registers[28][27]$_SDFFCE_PN0P_  (.D(_01052_),
    .CK(clknet_leaf_21_clk),
    .Q(\registers[28][27] ),
    .QN(_06246_));
 DFF_X1 \registers[28][28]$_SDFFCE_PN0P_  (.D(_01053_),
    .CK(clknet_leaf_51_clk),
    .Q(\registers[28][28] ),
    .QN(_06245_));
 DFF_X1 \registers[28][29]$_SDFFCE_PN0P_  (.D(_01054_),
    .CK(clknet_leaf_50_clk),
    .Q(\registers[28][29] ),
    .QN(_06244_));
 DFF_X1 \registers[28][2]$_SDFFCE_PN0P_  (.D(_01055_),
    .CK(clknet_leaf_42_clk),
    .Q(\registers[28][2] ),
    .QN(_06243_));
 DFF_X1 \registers[28][30]$_SDFFCE_PN0P_  (.D(_01056_),
    .CK(clknet_leaf_51_clk),
    .Q(\registers[28][30] ),
    .QN(_06242_));
 DFF_X1 \registers[28][31]$_SDFFCE_PN0P_  (.D(_01057_),
    .CK(clknet_leaf_42_clk),
    .Q(\registers[28][31] ),
    .QN(_06241_));
 DFF_X1 \registers[28][3]$_SDFFCE_PN0P_  (.D(_01058_),
    .CK(clknet_leaf_41_clk),
    .Q(\registers[28][3] ),
    .QN(_06240_));
 DFF_X1 \registers[28][4]$_SDFFCE_PN0P_  (.D(_01059_),
    .CK(clknet_leaf_42_clk),
    .Q(\registers[28][4] ),
    .QN(_06239_));
 DFF_X1 \registers[28][5]$_SDFFCE_PN0P_  (.D(_01060_),
    .CK(clknet_leaf_42_clk),
    .Q(\registers[28][5] ),
    .QN(_06238_));
 DFF_X1 \registers[28][6]$_SDFFCE_PN0P_  (.D(_01061_),
    .CK(clknet_leaf_51_clk),
    .Q(\registers[28][6] ),
    .QN(_06237_));
 DFF_X1 \registers[28][7]$_SDFFCE_PN0P_  (.D(_01062_),
    .CK(clknet_leaf_51_clk),
    .Q(\registers[28][7] ),
    .QN(_06236_));
 DFF_X1 \registers[28][8]$_SDFFCE_PN0P_  (.D(_01063_),
    .CK(clknet_leaf_143_clk),
    .Q(\registers[28][8] ),
    .QN(_06235_));
 DFF_X1 \registers[28][9]$_SDFFCE_PN0P_  (.D(_01064_),
    .CK(clknet_leaf_143_clk),
    .Q(\registers[28][9] ),
    .QN(_06234_));
 DFF_X1 \registers[29][0]$_SDFFCE_PN0P_  (.D(_01065_),
    .CK(clknet_leaf_149_clk),
    .Q(\registers[29][0] ),
    .QN(_06233_));
 DFF_X1 \registers[29][10]$_SDFFCE_PN0P_  (.D(_01066_),
    .CK(clknet_leaf_149_clk),
    .Q(\registers[29][10] ),
    .QN(_06232_));
 DFF_X1 \registers[29][11]$_SDFFCE_PN0P_  (.D(_01067_),
    .CK(clknet_leaf_149_clk),
    .Q(\registers[29][11] ),
    .QN(_06231_));
 DFF_X1 \registers[29][12]$_SDFFCE_PN0P_  (.D(_01068_),
    .CK(clknet_leaf_149_clk),
    .Q(\registers[29][12] ),
    .QN(_06230_));
 DFF_X1 \registers[29][13]$_SDFFCE_PN0P_  (.D(_01069_),
    .CK(clknet_leaf_151_clk),
    .Q(\registers[29][13] ),
    .QN(_06229_));
 DFF_X1 \registers[29][14]$_SDFFCE_PN0P_  (.D(_01070_),
    .CK(clknet_leaf_151_clk),
    .Q(\registers[29][14] ),
    .QN(_06228_));
 DFF_X1 \registers[29][15]$_SDFFCE_PN0P_  (.D(_01071_),
    .CK(clknet_leaf_150_clk),
    .Q(\registers[29][15] ),
    .QN(_06227_));
 DFF_X1 \registers[29][16]$_SDFFCE_PN0P_  (.D(_01072_),
    .CK(clknet_leaf_151_clk),
    .Q(\registers[29][16] ),
    .QN(_06226_));
 DFF_X1 \registers[29][17]$_SDFFCE_PN0P_  (.D(_01073_),
    .CK(clknet_leaf_152_clk),
    .Q(\registers[29][17] ),
    .QN(_06225_));
 DFF_X1 \registers[29][18]$_SDFFCE_PN0P_  (.D(_01074_),
    .CK(clknet_leaf_152_clk),
    .Q(\registers[29][18] ),
    .QN(_06224_));
 DFF_X1 \registers[29][19]$_SDFFCE_PN0P_  (.D(_01075_),
    .CK(clknet_leaf_14_clk),
    .Q(\registers[29][19] ),
    .QN(_06223_));
 DFF_X1 \registers[29][1]$_SDFFCE_PN0P_  (.D(_01076_),
    .CK(clknet_leaf_14_clk),
    .Q(\registers[29][1] ),
    .QN(_06222_));
 DFF_X1 \registers[29][20]$_SDFFCE_PN0P_  (.D(_01077_),
    .CK(clknet_leaf_9_clk),
    .Q(\registers[29][20] ),
    .QN(_06221_));
 DFF_X1 \registers[29][21]$_SDFFCE_PN0P_  (.D(_01078_),
    .CK(clknet_leaf_9_clk),
    .Q(\registers[29][21] ),
    .QN(_06220_));
 DFF_X1 \registers[29][22]$_SDFFCE_PN0P_  (.D(_01079_),
    .CK(clknet_leaf_15_clk),
    .Q(\registers[29][22] ),
    .QN(_06219_));
 DFF_X1 \registers[29][23]$_SDFFCE_PN0P_  (.D(_01080_),
    .CK(clknet_leaf_24_clk),
    .Q(\registers[29][23] ),
    .QN(_06218_));
 DFF_X1 \registers[29][24]$_SDFFCE_PN0P_  (.D(_01081_),
    .CK(clknet_leaf_23_clk),
    .Q(\registers[29][24] ),
    .QN(_06217_));
 DFF_X1 \registers[29][25]$_SDFFCE_PN0P_  (.D(_01082_),
    .CK(clknet_leaf_23_clk),
    .Q(\registers[29][25] ),
    .QN(_06216_));
 DFF_X1 \registers[29][26]$_SDFFCE_PN0P_  (.D(_01083_),
    .CK(clknet_leaf_22_clk),
    .Q(\registers[29][26] ),
    .QN(_06215_));
 DFF_X1 \registers[29][27]$_SDFFCE_PN0P_  (.D(_01084_),
    .CK(clknet_leaf_21_clk),
    .Q(\registers[29][27] ),
    .QN(_06214_));
 DFF_X1 \registers[29][28]$_SDFFCE_PN0P_  (.D(_01085_),
    .CK(clknet_leaf_22_clk),
    .Q(\registers[29][28] ),
    .QN(_06213_));
 DFF_X1 \registers[29][29]$_SDFFCE_PN0P_  (.D(_01086_),
    .CK(clknet_leaf_22_clk),
    .Q(\registers[29][29] ),
    .QN(_06212_));
 DFF_X1 \registers[29][2]$_SDFFCE_PN0P_  (.D(_01087_),
    .CK(clknet_leaf_51_clk),
    .Q(\registers[29][2] ),
    .QN(_06211_));
 DFF_X1 \registers[29][30]$_SDFFCE_PN0P_  (.D(_00000_),
    .CK(clknet_leaf_53_clk),
    .Q(\registers[29][30] ),
    .QN(_06210_));
 DFF_X1 \registers[29][31]$_SDFFCE_PN0P_  (.D(_00001_),
    .CK(clknet_leaf_49_clk),
    .Q(\registers[29][31] ),
    .QN(_06209_));
 DFF_X1 \registers[29][3]$_SDFFCE_PN0P_  (.D(_00002_),
    .CK(clknet_leaf_48_clk),
    .Q(\registers[29][3] ),
    .QN(_06208_));
 DFF_X1 \registers[29][4]$_SDFFCE_PN0P_  (.D(_00003_),
    .CK(clknet_leaf_48_clk),
    .Q(\registers[29][4] ),
    .QN(_06207_));
 DFF_X1 \registers[29][5]$_SDFFCE_PN0P_  (.D(_00004_),
    .CK(clknet_leaf_48_clk),
    .Q(\registers[29][5] ),
    .QN(_06206_));
 DFF_X1 \registers[29][6]$_SDFFCE_PN0P_  (.D(_00005_),
    .CK(clknet_leaf_53_clk),
    .Q(\registers[29][6] ),
    .QN(_06205_));
 DFF_X1 \registers[29][7]$_SDFFCE_PN0P_  (.D(_00006_),
    .CK(clknet_leaf_53_clk),
    .Q(\registers[29][7] ),
    .QN(_06204_));
 DFF_X1 \registers[29][8]$_SDFFCE_PN0P_  (.D(_00007_),
    .CK(clknet_leaf_141_clk),
    .Q(\registers[29][8] ),
    .QN(_06203_));
 DFF_X1 \registers[29][9]$_SDFFCE_PN0P_  (.D(_00008_),
    .CK(clknet_leaf_140_clk),
    .Q(\registers[29][9] ),
    .QN(_06202_));
 DFF_X1 \registers[2][0]$_SDFFCE_PN0P_  (.D(_00009_),
    .CK(clknet_leaf_131_clk),
    .Q(\registers[2][0] ),
    .QN(_06201_));
 DFF_X1 \registers[2][10]$_SDFFCE_PN0P_  (.D(_00010_),
    .CK(clknet_leaf_129_clk),
    .Q(\registers[2][10] ),
    .QN(_06200_));
 DFF_X1 \registers[2][11]$_SDFFCE_PN0P_  (.D(_00011_),
    .CK(clknet_leaf_126_clk),
    .Q(\registers[2][11] ),
    .QN(_06199_));
 DFF_X1 \registers[2][12]$_SDFFCE_PN0P_  (.D(_00012_),
    .CK(clknet_leaf_129_clk),
    .Q(\registers[2][12] ),
    .QN(_06198_));
 DFF_X1 \registers[2][13]$_SDFFCE_PN0P_  (.D(_00013_),
    .CK(clknet_leaf_131_clk),
    .Q(\registers[2][13] ),
    .QN(_06197_));
 DFF_X1 \registers[2][14]$_SDFFCE_PN0P_  (.D(_00014_),
    .CK(clknet_leaf_129_clk),
    .Q(\registers[2][14] ),
    .QN(_06196_));
 DFF_X1 \registers[2][15]$_SDFFCE_PN0P_  (.D(_00015_),
    .CK(clknet_leaf_129_clk),
    .Q(\registers[2][15] ),
    .QN(_06195_));
 DFF_X1 \registers[2][16]$_SDFFCE_PN0P_  (.D(_00016_),
    .CK(clknet_leaf_130_clk),
    .Q(\registers[2][16] ),
    .QN(_06194_));
 DFF_X1 \registers[2][17]$_SDFFCE_PN0P_  (.D(_00017_),
    .CK(clknet_leaf_135_clk),
    .Q(\registers[2][17] ),
    .QN(_06193_));
 DFF_X1 \registers[2][18]$_SDFFCE_PN0P_  (.D(_00018_),
    .CK(clknet_leaf_137_clk),
    .Q(\registers[2][18] ),
    .QN(_06192_));
 DFF_X1 \registers[2][19]$_SDFFCE_PN0P_  (.D(_00019_),
    .CK(clknet_leaf_138_clk),
    .Q(\registers[2][19] ),
    .QN(_06191_));
 DFF_X1 \registers[2][1]$_SDFFCE_PN0P_  (.D(_00020_),
    .CK(clknet_leaf_138_clk),
    .Q(\registers[2][1] ),
    .QN(_06190_));
 DFF_X1 \registers[2][20]$_SDFFCE_PN0P_  (.D(_00021_),
    .CK(clknet_leaf_97_clk),
    .Q(\registers[2][20] ),
    .QN(_06189_));
 DFF_X1 \registers[2][21]$_SDFFCE_PN0P_  (.D(_00022_),
    .CK(clknet_leaf_97_clk),
    .Q(\registers[2][21] ),
    .QN(_06188_));
 DFF_X1 \registers[2][22]$_SDFFCE_PN0P_  (.D(_00023_),
    .CK(clknet_leaf_96_clk),
    .Q(\registers[2][22] ),
    .QN(_06187_));
 DFF_X1 \registers[2][23]$_SDFFCE_PN0P_  (.D(_00024_),
    .CK(clknet_leaf_96_clk),
    .Q(\registers[2][23] ),
    .QN(_06186_));
 DFF_X1 \registers[2][24]$_SDFFCE_PN0P_  (.D(_00025_),
    .CK(clknet_leaf_56_clk),
    .Q(\registers[2][24] ),
    .QN(_06185_));
 DFF_X1 \registers[2][25]$_SDFFCE_PN0P_  (.D(_00026_),
    .CK(clknet_leaf_56_clk),
    .Q(\registers[2][25] ),
    .QN(_06184_));
 DFF_X1 \registers[2][26]$_SDFFCE_PN0P_  (.D(_00027_),
    .CK(clknet_leaf_57_clk),
    .Q(\registers[2][26] ),
    .QN(_06183_));
 DFF_X1 \registers[2][27]$_SDFFCE_PN0P_  (.D(_00028_),
    .CK(clknet_leaf_56_clk),
    .Q(\registers[2][27] ),
    .QN(_06182_));
 DFF_X1 \registers[2][28]$_SDFFCE_PN0P_  (.D(_00029_),
    .CK(clknet_leaf_64_clk),
    .Q(\registers[2][28] ),
    .QN(_06181_));
 DFF_X1 \registers[2][29]$_SDFFCE_PN0P_  (.D(_00030_),
    .CK(clknet_leaf_63_clk),
    .Q(\registers[2][29] ),
    .QN(_06180_));
 DFF_X1 \registers[2][2]$_SDFFCE_PN0P_  (.D(_00031_),
    .CK(clknet_leaf_64_clk),
    .Q(\registers[2][2] ),
    .QN(_06179_));
 DFF_X1 \registers[2][30]$_SDFFCE_PN0P_  (.D(_00032_),
    .CK(clknet_leaf_67_clk),
    .Q(\registers[2][30] ),
    .QN(_06178_));
 DFF_X1 \registers[2][31]$_SDFFCE_PN0P_  (.D(_00033_),
    .CK(clknet_leaf_64_clk),
    .Q(\registers[2][31] ),
    .QN(_06177_));
 DFF_X1 \registers[2][3]$_SDFFCE_PN0P_  (.D(_00034_),
    .CK(clknet_leaf_64_clk),
    .Q(\registers[2][3] ),
    .QN(_06176_));
 DFF_X1 \registers[2][4]$_SDFFCE_PN0P_  (.D(_00035_),
    .CK(clknet_leaf_63_clk),
    .Q(\registers[2][4] ),
    .QN(_06175_));
 DFF_X1 \registers[2][5]$_SDFFCE_PN0P_  (.D(_00036_),
    .CK(clknet_leaf_61_clk),
    .Q(\registers[2][5] ),
    .QN(_06174_));
 DFF_X1 \registers[2][6]$_SDFFCE_PN0P_  (.D(_00037_),
    .CK(clknet_leaf_61_clk),
    .Q(\registers[2][6] ),
    .QN(_06173_));
 DFF_X1 \registers[2][7]$_SDFFCE_PN0P_  (.D(_00038_),
    .CK(clknet_leaf_58_clk),
    .Q(\registers[2][7] ),
    .QN(_06172_));
 DFF_X1 \registers[2][8]$_SDFFCE_PN0P_  (.D(_00039_),
    .CK(clknet_leaf_137_clk),
    .Q(\registers[2][8] ),
    .QN(_06171_));
 DFF_X1 \registers[2][9]$_SDFFCE_PN0P_  (.D(_00040_),
    .CK(clknet_leaf_137_clk),
    .Q(\registers[2][9] ),
    .QN(_06170_));
 DFF_X1 \registers[30][0]$_SDFFCE_PN0P_  (.D(_00041_),
    .CK(clknet_leaf_146_clk),
    .Q(\registers[30][0] ),
    .QN(_06169_));
 DFF_X1 \registers[30][10]$_SDFFCE_PN0P_  (.D(_00042_),
    .CK(clknet_leaf_148_clk),
    .Q(\registers[30][10] ),
    .QN(_06168_));
 DFF_X1 \registers[30][11]$_SDFFCE_PN0P_  (.D(_00043_),
    .CK(clknet_leaf_149_clk),
    .Q(\registers[30][11] ),
    .QN(_06167_));
 DFF_X1 \registers[30][12]$_SDFFCE_PN0P_  (.D(_00044_),
    .CK(clknet_leaf_149_clk),
    .Q(\registers[30][12] ),
    .QN(_06166_));
 DFF_X1 \registers[30][13]$_SDFFCE_PN0P_  (.D(_00045_),
    .CK(clknet_leaf_151_clk),
    .Q(\registers[30][13] ),
    .QN(_06165_));
 DFF_X1 \registers[30][14]$_SDFFCE_PN0P_  (.D(_00046_),
    .CK(clknet_leaf_152_clk),
    .Q(\registers[30][14] ),
    .QN(_06164_));
 DFF_X1 \registers[30][15]$_SDFFCE_PN0P_  (.D(_00047_),
    .CK(clknet_leaf_150_clk),
    .Q(\registers[30][15] ),
    .QN(_06163_));
 DFF_X1 \registers[30][16]$_SDFFCE_PN0P_  (.D(_00048_),
    .CK(clknet_leaf_145_clk),
    .Q(\registers[30][16] ),
    .QN(_06162_));
 DFF_X1 \registers[30][17]$_SDFFCE_PN0P_  (.D(_00049_),
    .CK(clknet_leaf_144_clk),
    .Q(\registers[30][17] ),
    .QN(_06161_));
 DFF_X1 \registers[30][18]$_SDFFCE_PN0P_  (.D(_00050_),
    .CK(clknet_leaf_143_clk),
    .Q(\registers[30][18] ),
    .QN(_06160_));
 DFF_X1 \registers[30][19]$_SDFFCE_PN0P_  (.D(_00051_),
    .CK(clknet_leaf_13_clk),
    .Q(\registers[30][19] ),
    .QN(_06159_));
 DFF_X1 \registers[30][1]$_SDFFCE_PN0P_  (.D(_00052_),
    .CK(clknet_leaf_14_clk),
    .Q(\registers[30][1] ),
    .QN(_06158_));
 DFF_X1 \registers[30][20]$_SDFFCE_PN0P_  (.D(_00053_),
    .CK(clknet_leaf_14_clk),
    .Q(\registers[30][20] ),
    .QN(_06157_));
 DFF_X1 \registers[30][21]$_SDFFCE_PN0P_  (.D(_00054_),
    .CK(clknet_leaf_15_clk),
    .Q(\registers[30][21] ),
    .QN(_06156_));
 DFF_X1 \registers[30][22]$_SDFFCE_PN0P_  (.D(_00055_),
    .CK(clknet_leaf_19_clk),
    .Q(\registers[30][22] ),
    .QN(_06155_));
 DFF_X1 \registers[30][23]$_SDFFCE_PN0P_  (.D(_00056_),
    .CK(clknet_leaf_20_clk),
    .Q(\registers[30][23] ),
    .QN(_06154_));
 DFF_X1 \registers[30][24]$_SDFFCE_PN0P_  (.D(_00057_),
    .CK(clknet_leaf_20_clk),
    .Q(\registers[30][24] ),
    .QN(_06153_));
 DFF_X1 \registers[30][25]$_SDFFCE_PN0P_  (.D(_00058_),
    .CK(clknet_leaf_20_clk),
    .Q(\registers[30][25] ),
    .QN(_06152_));
 DFF_X1 \registers[30][26]$_SDFFCE_PN0P_  (.D(_00059_),
    .CK(clknet_leaf_21_clk),
    .Q(\registers[30][26] ),
    .QN(_06151_));
 DFF_X1 \registers[30][27]$_SDFFCE_PN0P_  (.D(_00060_),
    .CK(clknet_leaf_21_clk),
    .Q(\registers[30][27] ),
    .QN(_06150_));
 DFF_X1 \registers[30][28]$_SDFFCE_PN0P_  (.D(_00061_),
    .CK(clknet_leaf_51_clk),
    .Q(\registers[30][28] ),
    .QN(_06149_));
 DFF_X1 \registers[30][29]$_SDFFCE_PN0P_  (.D(_00062_),
    .CK(clknet_leaf_50_clk),
    .Q(\registers[30][29] ),
    .QN(_06148_));
 DFF_X1 \registers[30][2]$_SDFFCE_PN0P_  (.D(_00063_),
    .CK(clknet_leaf_50_clk),
    .Q(\registers[30][2] ),
    .QN(_06147_));
 DFF_X1 \registers[30][30]$_SDFFCE_PN0P_  (.D(_00064_),
    .CK(clknet_leaf_51_clk),
    .Q(\registers[30][30] ),
    .QN(_06146_));
 DFF_X1 \registers[30][31]$_SDFFCE_PN0P_  (.D(_00065_),
    .CK(clknet_leaf_49_clk),
    .Q(\registers[30][31] ),
    .QN(_06145_));
 DFF_X1 \registers[30][3]$_SDFFCE_PN0P_  (.D(_00066_),
    .CK(clknet_leaf_50_clk),
    .Q(\registers[30][3] ),
    .QN(_06144_));
 DFF_X1 \registers[30][4]$_SDFFCE_PN0P_  (.D(_00067_),
    .CK(clknet_leaf_49_clk),
    .Q(\registers[30][4] ),
    .QN(_06143_));
 DFF_X1 \registers[30][5]$_SDFFCE_PN0P_  (.D(_00068_),
    .CK(clknet_leaf_50_clk),
    .Q(\registers[30][5] ),
    .QN(_06142_));
 DFF_X1 \registers[30][6]$_SDFFCE_PN0P_  (.D(_00069_),
    .CK(clknet_leaf_52_clk),
    .Q(\registers[30][6] ),
    .QN(_06141_));
 DFF_X1 \registers[30][7]$_SDFFCE_PN0P_  (.D(_00070_),
    .CK(clknet_leaf_52_clk),
    .Q(\registers[30][7] ),
    .QN(_06140_));
 DFF_X1 \registers[30][8]$_SDFFCE_PN0P_  (.D(_00071_),
    .CK(clknet_leaf_142_clk),
    .Q(\registers[30][8] ),
    .QN(_06139_));
 DFF_X1 \registers[30][9]$_SDFFCE_PN0P_  (.D(_00072_),
    .CK(clknet_leaf_143_clk),
    .Q(\registers[30][9] ),
    .QN(_06138_));
 DFF_X1 \registers[31][0]$_SDFFCE_PN0P_  (.D(_00073_),
    .CK(clknet_leaf_141_clk),
    .Q(\registers[31][0] ),
    .QN(_06137_));
 DFF_X1 \registers[31][10]$_SDFFCE_PN0P_  (.D(_00074_),
    .CK(clknet_leaf_128_clk),
    .Q(\registers[31][10] ),
    .QN(_06136_));
 DFF_X1 \registers[31][11]$_SDFFCE_PN0P_  (.D(_00075_),
    .CK(clknet_leaf_149_clk),
    .Q(\registers[31][11] ),
    .QN(_06135_));
 DFF_X1 \registers[31][12]$_SDFFCE_PN0P_  (.D(_00076_),
    .CK(clknet_leaf_128_clk),
    .Q(\registers[31][12] ),
    .QN(_06134_));
 DFF_X1 \registers[31][13]$_SDFFCE_PN0P_  (.D(_00077_),
    .CK(clknet_leaf_151_clk),
    .Q(\registers[31][13] ),
    .QN(_06133_));
 DFF_X1 \registers[31][14]$_SDFFCE_PN0P_  (.D(_00078_),
    .CK(clknet_leaf_153_clk),
    .Q(\registers[31][14] ),
    .QN(_06132_));
 DFF_X1 \registers[31][15]$_SDFFCE_PN0P_  (.D(_00079_),
    .CK(clknet_leaf_150_clk),
    .Q(\registers[31][15] ),
    .QN(_06131_));
 DFF_X1 \registers[31][16]$_SDFFCE_PN0P_  (.D(_00080_),
    .CK(clknet_leaf_144_clk),
    .Q(\registers[31][16] ),
    .QN(_06130_));
 DFF_X1 \registers[31][17]$_SDFFCE_PN0P_  (.D(_00081_),
    .CK(clknet_leaf_13_clk),
    .Q(\registers[31][17] ),
    .QN(_06129_));
 DFF_X1 \registers[31][18]$_SDFFCE_PN0P_  (.D(_00082_),
    .CK(clknet_leaf_13_clk),
    .Q(\registers[31][18] ),
    .QN(_06128_));
 DFF_X1 \registers[31][19]$_SDFFCE_PN0P_  (.D(_00083_),
    .CK(clknet_leaf_13_clk),
    .Q(\registers[31][19] ),
    .QN(_06127_));
 DFF_X1 \registers[31][1]$_SDFFCE_PN0P_  (.D(_00084_),
    .CK(clknet_leaf_13_clk),
    .Q(\registers[31][1] ),
    .QN(_06126_));
 DFF_X1 \registers[31][20]$_SDFFCE_PN0P_  (.D(_00085_),
    .CK(clknet_leaf_15_clk),
    .Q(\registers[31][20] ),
    .QN(_06125_));
 DFF_X1 \registers[31][21]$_SDFFCE_PN0P_  (.D(_00086_),
    .CK(clknet_leaf_15_clk),
    .Q(\registers[31][21] ),
    .QN(_06124_));
 DFF_X1 \registers[31][22]$_SDFFCE_PN0P_  (.D(_00087_),
    .CK(clknet_leaf_19_clk),
    .Q(\registers[31][22] ),
    .QN(_06123_));
 DFF_X1 \registers[31][23]$_SDFFCE_PN0P_  (.D(_00088_),
    .CK(clknet_leaf_19_clk),
    .Q(\registers[31][23] ),
    .QN(_06122_));
 DFF_X1 \registers[31][24]$_SDFFCE_PN0P_  (.D(_00089_),
    .CK(clknet_leaf_20_clk),
    .Q(\registers[31][24] ),
    .QN(_06121_));
 DFF_X1 \registers[31][25]$_SDFFCE_PN0P_  (.D(_00090_),
    .CK(clknet_leaf_20_clk),
    .Q(\registers[31][25] ),
    .QN(_06120_));
 DFF_X1 \registers[31][26]$_SDFFCE_PN0P_  (.D(_00091_),
    .CK(clknet_leaf_21_clk),
    .Q(\registers[31][26] ),
    .QN(_06119_));
 DFF_X1 \registers[31][27]$_SDFFCE_PN0P_  (.D(_00092_),
    .CK(clknet_leaf_21_clk),
    .Q(\registers[31][27] ),
    .QN(_06118_));
 DFF_X1 \registers[31][28]$_SDFFCE_PN0P_  (.D(_00093_),
    .CK(clknet_leaf_52_clk),
    .Q(\registers[31][28] ),
    .QN(_06117_));
 DFF_X1 \registers[31][29]$_SDFFCE_PN0P_  (.D(_00094_),
    .CK(clknet_leaf_50_clk),
    .Q(\registers[31][29] ),
    .QN(_06116_));
 DFF_X1 \registers[31][2]$_SDFFCE_PN0P_  (.D(_00095_),
    .CK(clknet_leaf_41_clk),
    .Q(\registers[31][2] ),
    .QN(_06115_));
 DFF_X1 \registers[31][30]$_SDFFCE_PN0P_  (.D(_00096_),
    .CK(clknet_leaf_53_clk),
    .Q(\registers[31][30] ),
    .QN(_06114_));
 DFF_X1 \registers[31][31]$_SDFFCE_PN0P_  (.D(_00097_),
    .CK(clknet_leaf_49_clk),
    .Q(\registers[31][31] ),
    .QN(_06113_));
 DFF_X1 \registers[31][3]$_SDFFCE_PN0P_  (.D(_00098_),
    .CK(clknet_leaf_48_clk),
    .Q(\registers[31][3] ),
    .QN(_06112_));
 DFF_X1 \registers[31][4]$_SDFFCE_PN0P_  (.D(_00099_),
    .CK(clknet_leaf_49_clk),
    .Q(\registers[31][4] ),
    .QN(_06111_));
 DFF_X1 \registers[31][5]$_SDFFCE_PN0P_  (.D(_00100_),
    .CK(clknet_leaf_54_clk),
    .Q(\registers[31][5] ),
    .QN(_06110_));
 DFF_X1 \registers[31][6]$_SDFFCE_PN0P_  (.D(_00101_),
    .CK(clknet_leaf_53_clk),
    .Q(\registers[31][6] ),
    .QN(_06109_));
 DFF_X1 \registers[31][7]$_SDFFCE_PN0P_  (.D(_00102_),
    .CK(clknet_leaf_54_clk),
    .Q(\registers[31][7] ),
    .QN(_06108_));
 DFF_X1 \registers[31][8]$_SDFFCE_PN0P_  (.D(_00103_),
    .CK(clknet_leaf_141_clk),
    .Q(\registers[31][8] ),
    .QN(_06107_));
 DFF_X1 \registers[31][9]$_SDFFCE_PN0P_  (.D(_00104_),
    .CK(clknet_leaf_141_clk),
    .Q(\registers[31][9] ),
    .QN(_06106_));
 DFF_X1 \registers[3][0]$_SDFFCE_PN0P_  (.D(_00105_),
    .CK(clknet_leaf_132_clk),
    .Q(\registers[3][0] ),
    .QN(_06105_));
 DFF_X1 \registers[3][10]$_SDFFCE_PN0P_  (.D(_00106_),
    .CK(clknet_leaf_126_clk),
    .Q(\registers[3][10] ),
    .QN(_06104_));
 DFF_X1 \registers[3][11]$_SDFFCE_PN0P_  (.D(_00107_),
    .CK(clknet_leaf_126_clk),
    .Q(\registers[3][11] ),
    .QN(_06103_));
 DFF_X1 \registers[3][12]$_SDFFCE_PN0P_  (.D(_00108_),
    .CK(clknet_leaf_126_clk),
    .Q(\registers[3][12] ),
    .QN(_06102_));
 DFF_X1 \registers[3][13]$_SDFFCE_PN0P_  (.D(_00109_),
    .CK(clknet_leaf_133_clk),
    .Q(\registers[3][13] ),
    .QN(_06101_));
 DFF_X1 \registers[3][14]$_SDFFCE_PN0P_  (.D(_00110_),
    .CK(clknet_leaf_124_clk),
    .Q(\registers[3][14] ),
    .QN(_06100_));
 DFF_X1 \registers[3][15]$_SDFFCE_PN0P_  (.D(_00111_),
    .CK(clknet_leaf_124_clk),
    .Q(\registers[3][15] ),
    .QN(_06099_));
 DFF_X1 \registers[3][16]$_SDFFCE_PN0P_  (.D(_00112_),
    .CK(clknet_leaf_132_clk),
    .Q(\registers[3][16] ),
    .QN(_06098_));
 DFF_X1 \registers[3][17]$_SDFFCE_PN0P_  (.D(_00113_),
    .CK(clknet_leaf_134_clk),
    .Q(\registers[3][17] ),
    .QN(_06097_));
 DFF_X1 \registers[3][18]$_SDFFCE_PN0P_  (.D(_00114_),
    .CK(clknet_leaf_134_clk),
    .Q(\registers[3][18] ),
    .QN(_06096_));
 DFF_X1 \registers[3][19]$_SDFFCE_PN0P_  (.D(_00115_),
    .CK(clknet_leaf_98_clk),
    .Q(\registers[3][19] ),
    .QN(_06095_));
 DFF_X1 \registers[3][1]$_SDFFCE_PN0P_  (.D(_00116_),
    .CK(clknet_leaf_98_clk),
    .Q(\registers[3][1] ),
    .QN(_06094_));
 DFF_X1 \registers[3][20]$_SDFFCE_PN0P_  (.D(_00117_),
    .CK(clknet_leaf_98_clk),
    .Q(\registers[3][20] ),
    .QN(_06093_));
 DFF_X1 \registers[3][21]$_SDFFCE_PN0P_  (.D(_00118_),
    .CK(clknet_leaf_98_clk),
    .Q(\registers[3][21] ),
    .QN(_06092_));
 DFF_X1 \registers[3][22]$_SDFFCE_PN0P_  (.D(_00119_),
    .CK(clknet_leaf_95_clk),
    .Q(\registers[3][22] ),
    .QN(_06091_));
 DFF_X1 \registers[3][23]$_SDFFCE_PN0P_  (.D(_00120_),
    .CK(clknet_leaf_95_clk),
    .Q(\registers[3][23] ),
    .QN(_06090_));
 DFF_X1 \registers[3][24]$_SDFFCE_PN0P_  (.D(_00121_),
    .CK(clknet_leaf_95_clk),
    .Q(\registers[3][24] ),
    .QN(_06089_));
 DFF_X1 \registers[3][25]$_SDFFCE_PN0P_  (.D(_00122_),
    .CK(clknet_leaf_95_clk),
    .Q(\registers[3][25] ),
    .QN(_06088_));
 DFF_X1 \registers[3][26]$_SDFFCE_PN0P_  (.D(_00123_),
    .CK(clknet_leaf_59_clk),
    .Q(\registers[3][26] ),
    .QN(_06087_));
 DFF_X1 \registers[3][27]$_SDFFCE_PN0P_  (.D(_00124_),
    .CK(clknet_leaf_93_clk),
    .Q(\registers[3][27] ),
    .QN(_06086_));
 DFF_X1 \registers[3][28]$_SDFFCE_PN0P_  (.D(_00125_),
    .CK(clknet_leaf_67_clk),
    .Q(\registers[3][28] ),
    .QN(_06085_));
 DFF_X1 \registers[3][29]$_SDFFCE_PN0P_  (.D(_00126_),
    .CK(clknet_leaf_68_clk),
    .Q(\registers[3][29] ),
    .QN(_06084_));
 DFF_X1 \registers[3][2]$_SDFFCE_PN0P_  (.D(_00127_),
    .CK(clknet_leaf_67_clk),
    .Q(\registers[3][2] ),
    .QN(_06083_));
 DFF_X1 \registers[3][30]$_SDFFCE_PN0P_  (.D(_00128_),
    .CK(clknet_leaf_68_clk),
    .Q(\registers[3][30] ),
    .QN(_06082_));
 DFF_X1 \registers[3][31]$_SDFFCE_PN0P_  (.D(_00129_),
    .CK(clknet_leaf_68_clk),
    .Q(\registers[3][31] ),
    .QN(_06081_));
 DFF_X1 \registers[3][3]$_SDFFCE_PN0P_  (.D(_00130_),
    .CK(clknet_leaf_67_clk),
    .Q(\registers[3][3] ),
    .QN(_06080_));
 DFF_X1 \registers[3][4]$_SDFFCE_PN0P_  (.D(_00131_),
    .CK(clknet_leaf_67_clk),
    .Q(\registers[3][4] ),
    .QN(_06079_));
 DFF_X1 \registers[3][5]$_SDFFCE_PN0P_  (.D(_00132_),
    .CK(clknet_leaf_68_clk),
    .Q(\registers[3][5] ),
    .QN(_06078_));
 DFF_X1 \registers[3][6]$_SDFFCE_PN0P_  (.D(_00133_),
    .CK(clknet_leaf_61_clk),
    .Q(\registers[3][6] ),
    .QN(_06077_));
 DFF_X1 \registers[3][7]$_SDFFCE_PN0P_  (.D(_00134_),
    .CK(clknet_leaf_59_clk),
    .Q(\registers[3][7] ),
    .QN(_06076_));
 DFF_X1 \registers[3][8]$_SDFFCE_PN0P_  (.D(_00135_),
    .CK(clknet_leaf_134_clk),
    .Q(\registers[3][8] ),
    .QN(_06075_));
 DFF_X1 \registers[3][9]$_SDFFCE_PN0P_  (.D(_00136_),
    .CK(clknet_leaf_134_clk),
    .Q(\registers[3][9] ),
    .QN(_06074_));
 DFF_X1 \registers[4][0]$_SDFFCE_PN0P_  (.D(_00137_),
    .CK(clknet_leaf_134_clk),
    .Q(\registers[4][0] ),
    .QN(_06073_));
 DFF_X1 \registers[4][10]$_SDFFCE_PN0P_  (.D(_00138_),
    .CK(clknet_leaf_125_clk),
    .Q(\registers[4][10] ),
    .QN(_06072_));
 DFF_X1 \registers[4][11]$_SDFFCE_PN0P_  (.D(_00139_),
    .CK(clknet_leaf_125_clk),
    .Q(\registers[4][11] ),
    .QN(_06071_));
 DFF_X1 \registers[4][12]$_SDFFCE_PN0P_  (.D(_00140_),
    .CK(clknet_leaf_119_clk),
    .Q(\registers[4][12] ),
    .QN(_06070_));
 DFF_X1 \registers[4][13]$_SDFFCE_PN0P_  (.D(_00141_),
    .CK(clknet_leaf_133_clk),
    .Q(\registers[4][13] ),
    .QN(_06069_));
 DFF_X1 \registers[4][14]$_SDFFCE_PN0P_  (.D(_00142_),
    .CK(clknet_leaf_125_clk),
    .Q(\registers[4][14] ),
    .QN(_06068_));
 DFF_X1 \registers[4][15]$_SDFFCE_PN0P_  (.D(_00143_),
    .CK(clknet_leaf_119_clk),
    .Q(\registers[4][15] ),
    .QN(_06067_));
 DFF_X1 \registers[4][16]$_SDFFCE_PN0P_  (.D(_00144_),
    .CK(clknet_leaf_124_clk),
    .Q(\registers[4][16] ),
    .QN(_06066_));
 DFF_X1 \registers[4][17]$_SDFFCE_PN0P_  (.D(_00145_),
    .CK(clknet_leaf_101_clk),
    .Q(\registers[4][17] ),
    .QN(_06065_));
 DFF_X1 \registers[4][18]$_SDFFCE_PN0P_  (.D(_00146_),
    .CK(clknet_leaf_101_clk),
    .Q(\registers[4][18] ),
    .QN(_06064_));
 DFF_X1 \registers[4][19]$_SDFFCE_PN0P_  (.D(_00147_),
    .CK(clknet_leaf_99_clk),
    .Q(\registers[4][19] ),
    .QN(_06063_));
 DFF_X1 \registers[4][1]$_SDFFCE_PN0P_  (.D(_00148_),
    .CK(clknet_leaf_100_clk),
    .Q(\registers[4][1] ),
    .QN(_06062_));
 DFF_X1 \registers[4][20]$_SDFFCE_PN0P_  (.D(_00149_),
    .CK(clknet_leaf_99_clk),
    .Q(\registers[4][20] ),
    .QN(_06061_));
 DFF_X1 \registers[4][21]$_SDFFCE_PN0P_  (.D(_00150_),
    .CK(clknet_leaf_99_clk),
    .Q(\registers[4][21] ),
    .QN(_06060_));
 DFF_X1 \registers[4][22]$_SDFFCE_PN0P_  (.D(_00151_),
    .CK(clknet_leaf_94_clk),
    .Q(\registers[4][22] ),
    .QN(_06059_));
 DFF_X1 \registers[4][23]$_SDFFCE_PN0P_  (.D(_00152_),
    .CK(clknet_leaf_94_clk),
    .Q(\registers[4][23] ),
    .QN(_06058_));
 DFF_X1 \registers[4][24]$_SDFFCE_PN0P_  (.D(_00153_),
    .CK(clknet_leaf_94_clk),
    .Q(\registers[4][24] ),
    .QN(_06057_));
 DFF_X1 \registers[4][25]$_SDFFCE_PN0P_  (.D(_00154_),
    .CK(clknet_leaf_94_clk),
    .Q(\registers[4][25] ),
    .QN(_06056_));
 DFF_X1 \registers[4][26]$_SDFFCE_PN0P_  (.D(_00155_),
    .CK(clknet_leaf_92_clk),
    .Q(\registers[4][26] ),
    .QN(_06055_));
 DFF_X1 \registers[4][27]$_SDFFCE_PN0P_  (.D(_00156_),
    .CK(clknet_leaf_92_clk),
    .Q(\registers[4][27] ),
    .QN(_06054_));
 DFF_X1 \registers[4][28]$_SDFFCE_PN0P_  (.D(_00157_),
    .CK(clknet_leaf_69_clk),
    .Q(\registers[4][28] ),
    .QN(_06053_));
 DFF_X1 \registers[4][29]$_SDFFCE_PN0P_  (.D(_00158_),
    .CK(clknet_leaf_69_clk),
    .Q(\registers[4][29] ),
    .QN(_06052_));
 DFF_X1 \registers[4][2]$_SDFFCE_PN0P_  (.D(_00159_),
    .CK(clknet_leaf_68_clk),
    .Q(\registers[4][2] ),
    .QN(_06051_));
 DFF_X1 \registers[4][30]$_SDFFCE_PN0P_  (.D(_00160_),
    .CK(clknet_leaf_74_clk),
    .Q(\registers[4][30] ),
    .QN(_06050_));
 DFF_X1 \registers[4][31]$_SDFFCE_PN0P_  (.D(_00161_),
    .CK(clknet_leaf_68_clk),
    .Q(\registers[4][31] ),
    .QN(_06049_));
 DFF_X1 \registers[4][3]$_SDFFCE_PN0P_  (.D(_00162_),
    .CK(clknet_leaf_69_clk),
    .Q(\registers[4][3] ),
    .QN(_06048_));
 DFF_X1 \registers[4][4]$_SDFFCE_PN0P_  (.D(_00163_),
    .CK(clknet_leaf_68_clk),
    .Q(\registers[4][4] ),
    .QN(_06047_));
 DFF_X1 \registers[4][5]$_SDFFCE_PN0P_  (.D(_00164_),
    .CK(clknet_leaf_68_clk),
    .Q(\registers[4][5] ),
    .QN(_06046_));
 DFF_X1 \registers[4][6]$_SDFFCE_PN0P_  (.D(_00165_),
    .CK(clknet_leaf_60_clk),
    .Q(\registers[4][6] ),
    .QN(_06045_));
 DFF_X1 \registers[4][7]$_SDFFCE_PN0P_  (.D(_00166_),
    .CK(clknet_leaf_92_clk),
    .Q(\registers[4][7] ),
    .QN(_06044_));
 DFF_X1 \registers[4][8]$_SDFFCE_PN0P_  (.D(_00167_),
    .CK(clknet_leaf_100_clk),
    .Q(\registers[4][8] ),
    .QN(_06043_));
 DFF_X1 \registers[4][9]$_SDFFCE_PN0P_  (.D(_00168_),
    .CK(clknet_leaf_100_clk),
    .Q(\registers[4][9] ),
    .QN(_06042_));
 DFF_X1 \registers[5][0]$_SDFFCE_PN0P_  (.D(_00169_),
    .CK(clknet_leaf_133_clk),
    .Q(\registers[5][0] ),
    .QN(_06041_));
 DFF_X1 \registers[5][10]$_SDFFCE_PN0P_  (.D(_00170_),
    .CK(clknet_leaf_124_clk),
    .Q(\registers[5][10] ),
    .QN(_06040_));
 DFF_X1 \registers[5][11]$_SDFFCE_PN0P_  (.D(_00171_),
    .CK(clknet_leaf_125_clk),
    .Q(\registers[5][11] ),
    .QN(_06039_));
 DFF_X1 \registers[5][12]$_SDFFCE_PN0P_  (.D(_00172_),
    .CK(clknet_leaf_119_clk),
    .Q(\registers[5][12] ),
    .QN(_06038_));
 DFF_X1 \registers[5][13]$_SDFFCE_PN0P_  (.D(_00173_),
    .CK(clknet_leaf_133_clk),
    .Q(\registers[5][13] ),
    .QN(_06037_));
 DFF_X1 \registers[5][14]$_SDFFCE_PN0P_  (.D(_00174_),
    .CK(clknet_leaf_124_clk),
    .Q(\registers[5][14] ),
    .QN(_06036_));
 DFF_X1 \registers[5][15]$_SDFFCE_PN0P_  (.D(_00175_),
    .CK(clknet_leaf_119_clk),
    .Q(\registers[5][15] ),
    .QN(_06035_));
 DFF_X1 \registers[5][16]$_SDFFCE_PN0P_  (.D(_00176_),
    .CK(clknet_leaf_124_clk),
    .Q(\registers[5][16] ),
    .QN(_06034_));
 DFF_X1 \registers[5][17]$_SDFFCE_PN0P_  (.D(_00177_),
    .CK(clknet_leaf_101_clk),
    .Q(\registers[5][17] ),
    .QN(_06033_));
 DFF_X1 \registers[5][18]$_SDFFCE_PN0P_  (.D(_00178_),
    .CK(clknet_leaf_101_clk),
    .Q(\registers[5][18] ),
    .QN(_06032_));
 DFF_X1 \registers[5][19]$_SDFFCE_PN0P_  (.D(_00179_),
    .CK(clknet_leaf_104_clk),
    .Q(\registers[5][19] ),
    .QN(_06031_));
 DFF_X1 \registers[5][1]$_SDFFCE_PN0P_  (.D(_00180_),
    .CK(clknet_leaf_100_clk),
    .Q(\registers[5][1] ),
    .QN(_06030_));
 DFF_X1 \registers[5][20]$_SDFFCE_PN0P_  (.D(_00181_),
    .CK(clknet_leaf_104_clk),
    .Q(\registers[5][20] ),
    .QN(_06029_));
 DFF_X1 \registers[5][21]$_SDFFCE_PN0P_  (.D(_00182_),
    .CK(clknet_leaf_90_clk),
    .Q(\registers[5][21] ),
    .QN(_06028_));
 DFF_X1 \registers[5][22]$_SDFFCE_PN0P_  (.D(_00183_),
    .CK(clknet_leaf_94_clk),
    .Q(\registers[5][22] ),
    .QN(_06027_));
 DFF_X1 \registers[5][23]$_SDFFCE_PN0P_  (.D(_00184_),
    .CK(clknet_leaf_94_clk),
    .Q(\registers[5][23] ),
    .QN(_06026_));
 DFF_X1 \registers[5][24]$_SDFFCE_PN0P_  (.D(_00185_),
    .CK(clknet_leaf_93_clk),
    .Q(\registers[5][24] ),
    .QN(_06025_));
 DFF_X1 \registers[5][25]$_SDFFCE_PN0P_  (.D(_00186_),
    .CK(clknet_leaf_94_clk),
    .Q(\registers[5][25] ),
    .QN(_06024_));
 DFF_X1 \registers[5][26]$_SDFFCE_PN0P_  (.D(_00187_),
    .CK(clknet_leaf_92_clk),
    .Q(\registers[5][26] ),
    .QN(_06023_));
 DFF_X1 \registers[5][27]$_SDFFCE_PN0P_  (.D(_00188_),
    .CK(clknet_leaf_92_clk),
    .Q(\registers[5][27] ),
    .QN(_06022_));
 DFF_X1 \registers[5][28]$_SDFFCE_PN0P_  (.D(_00189_),
    .CK(clknet_leaf_69_clk),
    .Q(\registers[5][28] ),
    .QN(_06021_));
 DFF_X1 \registers[5][29]$_SDFFCE_PN0P_  (.D(_00190_),
    .CK(clknet_leaf_69_clk),
    .Q(\registers[5][29] ),
    .QN(_06020_));
 DFF_X1 \registers[5][2]$_SDFFCE_PN0P_  (.D(_00191_),
    .CK(clknet_leaf_69_clk),
    .Q(\registers[5][2] ),
    .QN(_06019_));
 DFF_X1 \registers[5][30]$_SDFFCE_PN0P_  (.D(_00192_),
    .CK(clknet_leaf_73_clk),
    .Q(\registers[5][30] ),
    .QN(_06018_));
 DFF_X1 \registers[5][31]$_SDFFCE_PN0P_  (.D(_00193_),
    .CK(clknet_leaf_69_clk),
    .Q(\registers[5][31] ),
    .QN(_06017_));
 DFF_X1 \registers[5][3]$_SDFFCE_PN0P_  (.D(_00194_),
    .CK(clknet_leaf_74_clk),
    .Q(\registers[5][3] ),
    .QN(_06016_));
 DFF_X1 \registers[5][4]$_SDFFCE_PN0P_  (.D(_00195_),
    .CK(clknet_leaf_70_clk),
    .Q(\registers[5][4] ),
    .QN(_06015_));
 DFF_X1 \registers[5][5]$_SDFFCE_PN0P_  (.D(_00196_),
    .CK(clknet_leaf_70_clk),
    .Q(\registers[5][5] ),
    .QN(_06014_));
 DFF_X1 \registers[5][6]$_SDFFCE_PN0P_  (.D(_00197_),
    .CK(clknet_leaf_60_clk),
    .Q(\registers[5][6] ),
    .QN(_06013_));
 DFF_X1 \registers[5][7]$_SDFFCE_PN0P_  (.D(_00198_),
    .CK(clknet_leaf_60_clk),
    .Q(\registers[5][7] ),
    .QN(_06012_));
 DFF_X1 \registers[5][8]$_SDFFCE_PN0P_  (.D(_00199_),
    .CK(clknet_leaf_101_clk),
    .Q(\registers[5][8] ),
    .QN(_06011_));
 DFF_X1 \registers[5][9]$_SDFFCE_PN0P_  (.D(_00200_),
    .CK(clknet_leaf_133_clk),
    .Q(\registers[5][9] ),
    .QN(_06010_));
 DFF_X1 \registers[6][0]$_SDFFCE_PN0P_  (.D(_00201_),
    .CK(clknet_leaf_131_clk),
    .Q(\registers[6][0] ),
    .QN(_06009_));
 DFF_X1 \registers[6][10]$_SDFFCE_PN0P_  (.D(_00202_),
    .CK(clknet_leaf_128_clk),
    .Q(\registers[6][10] ),
    .QN(_06008_));
 DFF_X1 \registers[6][11]$_SDFFCE_PN0P_  (.D(_00203_),
    .CK(clknet_leaf_128_clk),
    .Q(\registers[6][11] ),
    .QN(_06007_));
 DFF_X1 \registers[6][12]$_SDFFCE_PN0P_  (.D(_00204_),
    .CK(clknet_leaf_128_clk),
    .Q(\registers[6][12] ),
    .QN(_06006_));
 DFF_X1 \registers[6][13]$_SDFFCE_PN0P_  (.D(_00205_),
    .CK(clknet_leaf_130_clk),
    .Q(\registers[6][13] ),
    .QN(_06005_));
 DFF_X1 \registers[6][14]$_SDFFCE_PN0P_  (.D(_00206_),
    .CK(clknet_leaf_128_clk),
    .Q(\registers[6][14] ),
    .QN(_06004_));
 DFF_X1 \registers[6][15]$_SDFFCE_PN0P_  (.D(_00207_),
    .CK(clknet_leaf_130_clk),
    .Q(\registers[6][15] ),
    .QN(_06003_));
 DFF_X1 \registers[6][16]$_SDFFCE_PN0P_  (.D(_00208_),
    .CK(clknet_leaf_130_clk),
    .Q(\registers[6][16] ),
    .QN(_06002_));
 DFF_X1 \registers[6][17]$_SDFFCE_PN0P_  (.D(_00209_),
    .CK(clknet_leaf_136_clk),
    .Q(\registers[6][17] ),
    .QN(_06001_));
 DFF_X1 \registers[6][18]$_SDFFCE_PN0P_  (.D(_00210_),
    .CK(clknet_leaf_136_clk),
    .Q(\registers[6][18] ),
    .QN(_06000_));
 DFF_X1 \registers[6][19]$_SDFFCE_PN0P_  (.D(_00211_),
    .CK(clknet_leaf_138_clk),
    .Q(\registers[6][19] ),
    .QN(_05999_));
 DFF_X1 \registers[6][1]$_SDFFCE_PN0P_  (.D(_00212_),
    .CK(clknet_leaf_138_clk),
    .Q(\registers[6][1] ),
    .QN(_05998_));
 DFF_X1 \registers[6][20]$_SDFFCE_PN0P_  (.D(_00213_),
    .CK(clknet_leaf_139_clk),
    .Q(\registers[6][20] ),
    .QN(_05997_));
 DFF_X1 \registers[6][21]$_SDFFCE_PN0P_  (.D(_00214_),
    .CK(clknet_leaf_139_clk),
    .Q(\registers[6][21] ),
    .QN(_05996_));
 DFF_X1 \registers[6][22]$_SDFFCE_PN0P_  (.D(_00215_),
    .CK(clknet_leaf_97_clk),
    .Q(\registers[6][22] ),
    .QN(_05995_));
 DFF_X1 \registers[6][23]$_SDFFCE_PN0P_  (.D(_00216_),
    .CK(clknet_leaf_55_clk),
    .Q(\registers[6][23] ),
    .QN(_05994_));
 DFF_X1 \registers[6][24]$_SDFFCE_PN0P_  (.D(_00217_),
    .CK(clknet_leaf_55_clk),
    .Q(\registers[6][24] ),
    .QN(_05993_));
 DFF_X1 \registers[6][25]$_SDFFCE_PN0P_  (.D(_00218_),
    .CK(clknet_leaf_56_clk),
    .Q(\registers[6][25] ),
    .QN(_05992_));
 DFF_X1 \registers[6][26]$_SDFFCE_PN0P_  (.D(_00219_),
    .CK(clknet_leaf_57_clk),
    .Q(\registers[6][26] ),
    .QN(_05991_));
 DFF_X1 \registers[6][27]$_SDFFCE_PN0P_  (.D(_00220_),
    .CK(clknet_leaf_57_clk),
    .Q(\registers[6][27] ),
    .QN(_05990_));
 DFF_X1 \registers[6][28]$_SDFFCE_PN0P_  (.D(_00221_),
    .CK(clknet_leaf_65_clk),
    .Q(\registers[6][28] ),
    .QN(_05989_));
 DFF_X1 \registers[6][29]$_SDFFCE_PN0P_  (.D(_00222_),
    .CK(clknet_leaf_63_clk),
    .Q(\registers[6][29] ),
    .QN(_05988_));
 DFF_X1 \registers[6][2]$_SDFFCE_PN0P_  (.D(_00223_),
    .CK(clknet_leaf_63_clk),
    .Q(\registers[6][2] ),
    .QN(_05987_));
 DFF_X1 \registers[6][30]$_SDFFCE_PN0P_  (.D(_00224_),
    .CK(clknet_leaf_65_clk),
    .Q(\registers[6][30] ),
    .QN(_05986_));
 DFF_X1 \registers[6][31]$_SDFFCE_PN0P_  (.D(_00225_),
    .CK(clknet_leaf_65_clk),
    .Q(\registers[6][31] ),
    .QN(_05985_));
 DFF_X1 \registers[6][3]$_SDFFCE_PN0P_  (.D(_00226_),
    .CK(clknet_leaf_62_clk),
    .Q(\registers[6][3] ),
    .QN(_05984_));
 DFF_X1 \registers[6][4]$_SDFFCE_PN0P_  (.D(_00227_),
    .CK(clknet_leaf_62_clk),
    .Q(\registers[6][4] ),
    .QN(_05983_));
 DFF_X1 \registers[6][5]$_SDFFCE_PN0P_  (.D(_00228_),
    .CK(clknet_leaf_62_clk),
    .Q(\registers[6][5] ),
    .QN(_05982_));
 DFF_X1 \registers[6][6]$_SDFFCE_PN0P_  (.D(_00229_),
    .CK(clknet_leaf_58_clk),
    .Q(\registers[6][6] ),
    .QN(_05981_));
 DFF_X1 \registers[6][7]$_SDFFCE_PN0P_  (.D(_00230_),
    .CK(clknet_leaf_58_clk),
    .Q(\registers[6][7] ),
    .QN(_05980_));
 DFF_X1 \registers[6][8]$_SDFFCE_PN0P_  (.D(_00231_),
    .CK(clknet_leaf_137_clk),
    .Q(\registers[6][8] ),
    .QN(_05979_));
 DFF_X1 \registers[6][9]$_SDFFCE_PN0P_  (.D(_00232_),
    .CK(clknet_leaf_138_clk),
    .Q(\registers[6][9] ),
    .QN(_05978_));
 DFF_X1 \registers[7][0]$_SDFFCE_PN0P_  (.D(_00233_),
    .CK(clknet_leaf_131_clk),
    .Q(\registers[7][0] ),
    .QN(_05977_));
 DFF_X1 \registers[7][10]$_SDFFCE_PN0P_  (.D(_00234_),
    .CK(clknet_leaf_127_clk),
    .Q(\registers[7][10] ),
    .QN(_05976_));
 DFF_X1 \registers[7][11]$_SDFFCE_PN0P_  (.D(_00235_),
    .CK(clknet_leaf_127_clk),
    .Q(\registers[7][11] ),
    .QN(_05975_));
 DFF_X1 \registers[7][12]$_SDFFCE_PN0P_  (.D(_00236_),
    .CK(clknet_leaf_127_clk),
    .Q(\registers[7][12] ),
    .QN(_05974_));
 DFF_X1 \registers[7][13]$_SDFFCE_PN0P_  (.D(_00237_),
    .CK(clknet_leaf_131_clk),
    .Q(\registers[7][13] ),
    .QN(_05973_));
 DFF_X1 \registers[7][14]$_SDFFCE_PN0P_  (.D(_00238_),
    .CK(clknet_leaf_130_clk),
    .Q(\registers[7][14] ),
    .QN(_05972_));
 DFF_X1 \registers[7][15]$_SDFFCE_PN0P_  (.D(_00239_),
    .CK(clknet_leaf_129_clk),
    .Q(\registers[7][15] ),
    .QN(_05971_));
 DFF_X1 \registers[7][16]$_SDFFCE_PN0P_  (.D(_00240_),
    .CK(clknet_leaf_130_clk),
    .Q(\registers[7][16] ),
    .QN(_05970_));
 DFF_X1 \registers[7][17]$_SDFFCE_PN0P_  (.D(_00241_),
    .CK(clknet_leaf_136_clk),
    .Q(\registers[7][17] ),
    .QN(_05969_));
 DFF_X1 \registers[7][18]$_SDFFCE_PN0P_  (.D(_00242_),
    .CK(clknet_leaf_136_clk),
    .Q(\registers[7][18] ),
    .QN(_05968_));
 DFF_X1 \registers[7][19]$_SDFFCE_PN0P_  (.D(_00243_),
    .CK(clknet_leaf_139_clk),
    .Q(\registers[7][19] ),
    .QN(_05967_));
 DFF_X1 \registers[7][1]$_SDFFCE_PN0P_  (.D(_00244_),
    .CK(clknet_leaf_138_clk),
    .Q(\registers[7][1] ),
    .QN(_05966_));
 DFF_X1 \registers[7][20]$_SDFFCE_PN0P_  (.D(_00245_),
    .CK(clknet_leaf_139_clk),
    .Q(\registers[7][20] ),
    .QN(_05965_));
 DFF_X1 \registers[7][21]$_SDFFCE_PN0P_  (.D(_00246_),
    .CK(clknet_leaf_97_clk),
    .Q(\registers[7][21] ),
    .QN(_05964_));
 DFF_X1 \registers[7][22]$_SDFFCE_PN0P_  (.D(_00247_),
    .CK(clknet_leaf_96_clk),
    .Q(\registers[7][22] ),
    .QN(_05963_));
 DFF_X1 \registers[7][23]$_SDFFCE_PN0P_  (.D(_00248_),
    .CK(clknet_leaf_55_clk),
    .Q(\registers[7][23] ),
    .QN(_05962_));
 DFF_X1 \registers[7][24]$_SDFFCE_PN0P_  (.D(_00249_),
    .CK(clknet_leaf_56_clk),
    .Q(\registers[7][24] ),
    .QN(_05961_));
 DFF_X1 \registers[7][25]$_SDFFCE_PN0P_  (.D(_00250_),
    .CK(clknet_leaf_57_clk),
    .Q(\registers[7][25] ),
    .QN(_05960_));
 DFF_X1 \registers[7][26]$_SDFFCE_PN0P_  (.D(_00251_),
    .CK(clknet_leaf_57_clk),
    .Q(\registers[7][26] ),
    .QN(_05959_));
 DFF_X1 \registers[7][27]$_SDFFCE_PN0P_  (.D(_00252_),
    .CK(clknet_leaf_57_clk),
    .Q(\registers[7][27] ),
    .QN(_05958_));
 DFF_X1 \registers[7][28]$_SDFFCE_PN0P_  (.D(_00253_),
    .CK(clknet_leaf_64_clk),
    .Q(\registers[7][28] ),
    .QN(_05957_));
 DFF_X1 \registers[7][29]$_SDFFCE_PN0P_  (.D(_00254_),
    .CK(clknet_leaf_63_clk),
    .Q(\registers[7][29] ),
    .QN(_05956_));
 DFF_X1 \registers[7][2]$_SDFFCE_PN0P_  (.D(_00255_),
    .CK(clknet_leaf_63_clk),
    .Q(\registers[7][2] ),
    .QN(_05955_));
 DFF_X1 \registers[7][30]$_SDFFCE_PN0P_  (.D(_00256_),
    .CK(clknet_leaf_64_clk),
    .Q(\registers[7][30] ),
    .QN(_05954_));
 DFF_X1 \registers[7][31]$_SDFFCE_PN0P_  (.D(_00257_),
    .CK(clknet_leaf_64_clk),
    .Q(\registers[7][31] ),
    .QN(_05953_));
 DFF_X1 \registers[7][3]$_SDFFCE_PN0P_  (.D(_00258_),
    .CK(clknet_leaf_63_clk),
    .Q(\registers[7][3] ),
    .QN(_05952_));
 DFF_X1 \registers[7][4]$_SDFFCE_PN0P_  (.D(_00259_),
    .CK(clknet_leaf_62_clk),
    .Q(\registers[7][4] ),
    .QN(_05951_));
 DFF_X1 \registers[7][5]$_SDFFCE_PN0P_  (.D(_00260_),
    .CK(clknet_leaf_62_clk),
    .Q(\registers[7][5] ),
    .QN(_05950_));
 DFF_X1 \registers[7][6]$_SDFFCE_PN0P_  (.D(_00261_),
    .CK(clknet_leaf_58_clk),
    .Q(\registers[7][6] ),
    .QN(_05949_));
 DFF_X1 \registers[7][7]$_SDFFCE_PN0P_  (.D(_00262_),
    .CK(clknet_leaf_58_clk),
    .Q(\registers[7][7] ),
    .QN(_05948_));
 DFF_X1 \registers[7][8]$_SDFFCE_PN0P_  (.D(_00263_),
    .CK(clknet_leaf_137_clk),
    .Q(\registers[7][8] ),
    .QN(_05947_));
 DFF_X1 \registers[7][9]$_SDFFCE_PN0P_  (.D(_00264_),
    .CK(clknet_leaf_137_clk),
    .Q(\registers[7][9] ),
    .QN(_05946_));
 DFF_X1 \registers[8][0]$_SDFFCE_PN0P_  (.D(_00265_),
    .CK(clknet_leaf_2_clk),
    .Q(\registers[8][0] ),
    .QN(_05945_));
 DFF_X1 \registers[8][10]$_SDFFCE_PN0P_  (.D(_00266_),
    .CK(clknet_leaf_155_clk),
    .Q(\registers[8][10] ),
    .QN(_05944_));
 DFF_X1 \registers[8][11]$_SDFFCE_PN0P_  (.D(_00267_),
    .CK(clknet_leaf_155_clk),
    .Q(\registers[8][11] ),
    .QN(_05943_));
 DFF_X1 \registers[8][12]$_SDFFCE_PN0P_  (.D(_00268_),
    .CK(clknet_leaf_155_clk),
    .Q(\registers[8][12] ),
    .QN(_05942_));
 DFF_X1 \registers[8][13]$_SDFFCE_PN0P_  (.D(_00269_),
    .CK(clknet_leaf_159_clk),
    .Q(\registers[8][13] ),
    .QN(_05941_));
 DFF_X1 \registers[8][14]$_SDFFCE_PN0P_  (.D(_00270_),
    .CK(clknet_leaf_0_clk),
    .Q(\registers[8][14] ),
    .QN(_05940_));
 DFF_X1 \registers[8][15]$_SDFFCE_PN0P_  (.D(_00271_),
    .CK(clknet_leaf_159_clk),
    .Q(\registers[8][15] ),
    .QN(_05939_));
 DFF_X1 \registers[8][16]$_SDFFCE_PN0P_  (.D(_00272_),
    .CK(clknet_leaf_159_clk),
    .Q(\registers[8][16] ),
    .QN(_05938_));
 DFF_X1 \registers[8][17]$_SDFFCE_PN0P_  (.D(_00273_),
    .CK(clknet_leaf_4_clk),
    .Q(\registers[8][17] ),
    .QN(_05937_));
 DFF_X1 \registers[8][18]$_SDFFCE_PN0P_  (.D(_00274_),
    .CK(clknet_leaf_5_clk),
    .Q(\registers[8][18] ),
    .QN(_05936_));
 DFF_X1 \registers[8][19]$_SDFFCE_PN0P_  (.D(_00275_),
    .CK(clknet_leaf_6_clk),
    .Q(\registers[8][19] ),
    .QN(_05935_));
 DFF_X1 \registers[8][1]$_SDFFCE_PN0P_  (.D(_00276_),
    .CK(clknet_leaf_6_clk),
    .Q(\registers[8][1] ),
    .QN(_05934_));
 DFF_X1 \registers[8][20]$_SDFFCE_PN0P_  (.D(_00277_),
    .CK(clknet_leaf_6_clk),
    .Q(\registers[8][20] ),
    .QN(_05933_));
 DFF_X1 \registers[8][21]$_SDFFCE_PN0P_  (.D(_00278_),
    .CK(clknet_leaf_7_clk),
    .Q(\registers[8][21] ),
    .QN(_05932_));
 DFF_X1 \registers[8][22]$_SDFFCE_PN0P_  (.D(_00279_),
    .CK(clknet_leaf_26_clk),
    .Q(\registers[8][22] ),
    .QN(_05931_));
 DFF_X1 \registers[8][23]$_SDFFCE_PN0P_  (.D(_00280_),
    .CK(clknet_leaf_25_clk),
    .Q(\registers[8][23] ),
    .QN(_05930_));
 DFF_X1 \registers[8][24]$_SDFFCE_PN0P_  (.D(_00281_),
    .CK(clknet_leaf_27_clk),
    .Q(\registers[8][24] ),
    .QN(_05929_));
 DFF_X1 \registers[8][25]$_SDFFCE_PN0P_  (.D(_00282_),
    .CK(clknet_leaf_27_clk),
    .Q(\registers[8][25] ),
    .QN(_05928_));
 DFF_X1 \registers[8][26]$_SDFFCE_PN0P_  (.D(_00283_),
    .CK(clknet_leaf_28_clk),
    .Q(\registers[8][26] ),
    .QN(_05927_));
 DFF_X1 \registers[8][27]$_SDFFCE_PN0P_  (.D(_00284_),
    .CK(clknet_leaf_28_clk),
    .Q(\registers[8][27] ),
    .QN(_05926_));
 DFF_X1 \registers[8][28]$_SDFFCE_PN0P_  (.D(_00285_),
    .CK(clknet_leaf_34_clk),
    .Q(\registers[8][28] ),
    .QN(_05925_));
 DFF_X1 \registers[8][29]$_SDFFCE_PN0P_  (.D(_00286_),
    .CK(clknet_leaf_34_clk),
    .Q(\registers[8][29] ),
    .QN(_05924_));
 DFF_X1 \registers[8][2]$_SDFFCE_PN0P_  (.D(_00287_),
    .CK(clknet_leaf_36_clk),
    .Q(\registers[8][2] ),
    .QN(_05923_));
 DFF_X1 \registers[8][30]$_SDFFCE_PN0P_  (.D(_00288_),
    .CK(clknet_leaf_37_clk),
    .Q(\registers[8][30] ),
    .QN(_05922_));
 DFF_X1 \registers[8][31]$_SDFFCE_PN0P_  (.D(_00289_),
    .CK(clknet_leaf_36_clk),
    .Q(\registers[8][31] ),
    .QN(_05921_));
 DFF_X1 \registers[8][3]$_SDFFCE_PN0P_  (.D(_00290_),
    .CK(clknet_leaf_38_clk),
    .Q(\registers[8][3] ),
    .QN(_05920_));
 DFF_X1 \registers[8][4]$_SDFFCE_PN0P_  (.D(_00291_),
    .CK(clknet_leaf_33_clk),
    .Q(\registers[8][4] ),
    .QN(_05919_));
 DFF_X1 \registers[8][5]$_SDFFCE_PN0P_  (.D(_00292_),
    .CK(clknet_leaf_33_clk),
    .Q(\registers[8][5] ),
    .QN(_05918_));
 DFF_X1 \registers[8][6]$_SDFFCE_PN0P_  (.D(_00293_),
    .CK(clknet_leaf_30_clk),
    .Q(\registers[8][6] ),
    .QN(_05917_));
 DFF_X1 \registers[8][7]$_SDFFCE_PN0P_  (.D(_00294_),
    .CK(clknet_leaf_30_clk),
    .Q(\registers[8][7] ),
    .QN(_05916_));
 DFF_X1 \registers[8][8]$_SDFFCE_PN0P_  (.D(_00295_),
    .CK(clknet_leaf_3_clk),
    .Q(\registers[8][8] ),
    .QN(_05915_));
 DFF_X1 \registers[8][9]$_SDFFCE_PN0P_  (.D(_00296_),
    .CK(clknet_leaf_5_clk),
    .Q(\registers[8][9] ),
    .QN(_05914_));
 DFF_X1 \registers[9][0]$_SDFFCE_PN0P_  (.D(_00297_),
    .CK(clknet_leaf_154_clk),
    .Q(\registers[9][0] ),
    .QN(_05913_));
 DFF_X1 \registers[9][10]$_SDFFCE_PN0P_  (.D(_00298_),
    .CK(clknet_leaf_154_clk),
    .Q(\registers[9][10] ),
    .QN(_05912_));
 DFF_X1 \registers[9][11]$_SDFFCE_PN0P_  (.D(_00299_),
    .CK(clknet_leaf_157_clk),
    .Q(\registers[9][11] ),
    .QN(_05911_));
 DFF_X1 \registers[9][12]$_SDFFCE_PN0P_  (.D(_00300_),
    .CK(clknet_leaf_154_clk),
    .Q(\registers[9][12] ),
    .QN(_05910_));
 DFF_X1 \registers[9][13]$_SDFFCE_PN0P_  (.D(_00301_),
    .CK(clknet_leaf_0_clk),
    .Q(\registers[9][13] ),
    .QN(_05909_));
 DFF_X1 \registers[9][14]$_SDFFCE_PN0P_  (.D(_00302_),
    .CK(clknet_leaf_158_clk),
    .Q(\registers[9][14] ),
    .QN(_05908_));
 DFF_X1 \registers[9][15]$_SDFFCE_PN0P_  (.D(_00303_),
    .CK(clknet_leaf_158_clk),
    .Q(\registers[9][15] ),
    .QN(_05907_));
 DFF_X1 \registers[9][16]$_SDFFCE_PN0P_  (.D(_00304_),
    .CK(clknet_leaf_0_clk),
    .Q(\registers[9][16] ),
    .QN(_05906_));
 DFF_X1 \registers[9][17]$_SDFFCE_PN0P_  (.D(_00305_),
    .CK(clknet_leaf_4_clk),
    .Q(\registers[9][17] ),
    .QN(_05905_));
 DFF_X1 \registers[9][18]$_SDFFCE_PN0P_  (.D(_00306_),
    .CK(clknet_leaf_4_clk),
    .Q(\registers[9][18] ),
    .QN(_05904_));
 DFF_X1 \registers[9][19]$_SDFFCE_PN0P_  (.D(_00307_),
    .CK(clknet_leaf_5_clk),
    .Q(\registers[9][19] ),
    .QN(_05903_));
 DFF_X1 \registers[9][1]$_SDFFCE_PN0P_  (.D(_00308_),
    .CK(clknet_leaf_5_clk),
    .Q(\registers[9][1] ),
    .QN(_05902_));
 DFF_X1 \registers[9][20]$_SDFFCE_PN0P_  (.D(_00309_),
    .CK(clknet_leaf_7_clk),
    .Q(\registers[9][20] ),
    .QN(_05901_));
 DFF_X1 \registers[9][21]$_SDFFCE_PN0P_  (.D(_00310_),
    .CK(clknet_leaf_7_clk),
    .Q(\registers[9][21] ),
    .QN(_05900_));
 DFF_X1 \registers[9][22]$_SDFFCE_PN0P_  (.D(_00311_),
    .CK(clknet_leaf_26_clk),
    .Q(\registers[9][22] ),
    .QN(_05899_));
 DFF_X1 \registers[9][23]$_SDFFCE_PN0P_  (.D(_00312_),
    .CK(clknet_leaf_26_clk),
    .Q(\registers[9][23] ),
    .QN(_05898_));
 DFF_X1 \registers[9][24]$_SDFFCE_PN0P_  (.D(_00313_),
    .CK(clknet_leaf_27_clk),
    .Q(\registers[9][24] ),
    .QN(_05897_));
 DFF_X1 \registers[9][25]$_SDFFCE_PN0P_  (.D(_00314_),
    .CK(clknet_leaf_27_clk),
    .Q(\registers[9][25] ),
    .QN(_05896_));
 DFF_X1 \registers[9][26]$_SDFFCE_PN0P_  (.D(_00315_),
    .CK(clknet_leaf_29_clk),
    .Q(\registers[9][26] ),
    .QN(_05895_));
 DFF_X1 \registers[9][27]$_SDFFCE_PN0P_  (.D(_00316_),
    .CK(clknet_leaf_29_clk),
    .Q(\registers[9][27] ),
    .QN(_05894_));
 DFF_X1 \registers[9][28]$_SDFFCE_PN0P_  (.D(_00317_),
    .CK(clknet_leaf_34_clk),
    .Q(\registers[9][28] ),
    .QN(_05893_));
 DFF_X1 \registers[9][29]$_SDFFCE_PN0P_  (.D(_00318_),
    .CK(clknet_leaf_35_clk),
    .Q(\registers[9][29] ),
    .QN(_05892_));
 DFF_X1 \registers[9][2]$_SDFFCE_PN0P_  (.D(_00319_),
    .CK(clknet_leaf_36_clk),
    .Q(\registers[9][2] ),
    .QN(_05891_));
 DFF_X1 \registers[9][30]$_SDFFCE_PN0P_  (.D(_00320_),
    .CK(clknet_leaf_37_clk),
    .Q(\registers[9][30] ),
    .QN(_05890_));
 DFF_X1 \registers[9][31]$_SDFFCE_PN0P_  (.D(_00321_),
    .CK(clknet_leaf_36_clk),
    .Q(\registers[9][31] ),
    .QN(_05889_));
 DFF_X1 \registers[9][3]$_SDFFCE_PN0P_  (.D(_00322_),
    .CK(clknet_leaf_37_clk),
    .Q(\registers[9][3] ),
    .QN(_05888_));
 DFF_X1 \registers[9][4]$_SDFFCE_PN0P_  (.D(_00323_),
    .CK(clknet_leaf_36_clk),
    .Q(\registers[9][4] ),
    .QN(_05887_));
 DFF_X1 \registers[9][5]$_SDFFCE_PN0P_  (.D(_00324_),
    .CK(clknet_leaf_35_clk),
    .Q(\registers[9][5] ),
    .QN(_05886_));
 DFF_X1 \registers[9][6]$_SDFFCE_PN0P_  (.D(_00325_),
    .CK(clknet_leaf_29_clk),
    .Q(\registers[9][6] ),
    .QN(_05885_));
 DFF_X1 \registers[9][7]$_SDFFCE_PN0P_  (.D(_00326_),
    .CK(clknet_leaf_29_clk),
    .Q(\registers[9][7] ),
    .QN(_05884_));
 DFF_X1 \registers[9][8]$_SDFFCE_PN0P_  (.D(_00327_),
    .CK(clknet_leaf_10_clk),
    .Q(\registers[9][8] ),
    .QN(_05883_));
 DFF_X1 \registers[9][9]$_SDFFCE_PN0P_  (.D(_00328_),
    .CK(clknet_leaf_5_clk),
    .Q(\registers[9][9] ),
    .QN(_05882_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_230 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_231 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_232 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_239 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_240 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_241 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_242 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_243 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_244 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_245 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_246 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_247 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_248 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_249 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_250 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_251 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_252 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_253 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_254 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_255 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_256 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_257 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_258 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_259 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_260 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_261 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_262 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_263 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_264 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_267 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_268 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_269 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_270 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_271 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_272 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_273 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_274 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_275 ();
 BUF_X1 input1 (.A(read_en1),
    .Z(net1));
 BUF_X1 input2 (.A(read_en2),
    .Z(net2));
 BUF_X2 input3 (.A(write_addr[3]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(write_en),
    .Z(net4));
 BUF_X1 output5 (.A(net5),
    .Z(read_data1[0]));
 BUF_X1 output6 (.A(net6),
    .Z(read_data1[10]));
 BUF_X1 output7 (.A(net7),
    .Z(read_data1[11]));
 BUF_X1 output8 (.A(net8),
    .Z(read_data1[12]));
 BUF_X1 output9 (.A(net9),
    .Z(read_data1[13]));
 BUF_X1 output10 (.A(net10),
    .Z(read_data1[14]));
 BUF_X1 output11 (.A(net11),
    .Z(read_data1[15]));
 BUF_X1 output12 (.A(net12),
    .Z(read_data1[16]));
 BUF_X1 output13 (.A(net13),
    .Z(read_data1[17]));
 BUF_X1 output14 (.A(net14),
    .Z(read_data1[18]));
 BUF_X1 output15 (.A(net15),
    .Z(read_data1[19]));
 BUF_X1 output16 (.A(net16),
    .Z(read_data1[1]));
 BUF_X1 output17 (.A(net17),
    .Z(read_data1[20]));
 BUF_X1 output18 (.A(net18),
    .Z(read_data1[21]));
 BUF_X1 output19 (.A(net19),
    .Z(read_data1[22]));
 BUF_X1 output20 (.A(net20),
    .Z(read_data1[23]));
 BUF_X1 output21 (.A(net21),
    .Z(read_data1[24]));
 BUF_X1 output22 (.A(net22),
    .Z(read_data1[25]));
 BUF_X1 output23 (.A(net23),
    .Z(read_data1[26]));
 BUF_X1 output24 (.A(net24),
    .Z(read_data1[27]));
 BUF_X1 output25 (.A(net25),
    .Z(read_data1[28]));
 BUF_X1 output26 (.A(net26),
    .Z(read_data1[29]));
 BUF_X1 output27 (.A(net27),
    .Z(read_data1[2]));
 BUF_X1 output28 (.A(net28),
    .Z(read_data1[30]));
 BUF_X1 output29 (.A(net29),
    .Z(read_data1[31]));
 BUF_X1 output30 (.A(net30),
    .Z(read_data1[3]));
 BUF_X1 output31 (.A(net31),
    .Z(read_data1[4]));
 BUF_X1 output32 (.A(net32),
    .Z(read_data1[5]));
 BUF_X1 output33 (.A(net33),
    .Z(read_data1[6]));
 BUF_X1 output34 (.A(net34),
    .Z(read_data1[7]));
 BUF_X1 output35 (.A(net35),
    .Z(read_data1[8]));
 BUF_X1 output36 (.A(net36),
    .Z(read_data1[9]));
 BUF_X1 output37 (.A(net37),
    .Z(read_data2[0]));
 BUF_X1 output38 (.A(net38),
    .Z(read_data2[10]));
 BUF_X1 output39 (.A(net39),
    .Z(read_data2[11]));
 BUF_X1 output40 (.A(net40),
    .Z(read_data2[12]));
 BUF_X1 output41 (.A(net41),
    .Z(read_data2[13]));
 BUF_X1 output42 (.A(net42),
    .Z(read_data2[14]));
 BUF_X1 output43 (.A(net43),
    .Z(read_data2[15]));
 BUF_X1 output44 (.A(net44),
    .Z(read_data2[16]));
 BUF_X1 output45 (.A(net45),
    .Z(read_data2[17]));
 BUF_X1 output46 (.A(net46),
    .Z(read_data2[18]));
 BUF_X1 output47 (.A(net47),
    .Z(read_data2[19]));
 BUF_X1 output48 (.A(net48),
    .Z(read_data2[1]));
 BUF_X1 output49 (.A(net49),
    .Z(read_data2[20]));
 BUF_X1 output50 (.A(net50),
    .Z(read_data2[21]));
 BUF_X1 output51 (.A(net51),
    .Z(read_data2[22]));
 BUF_X1 output52 (.A(net52),
    .Z(read_data2[23]));
 BUF_X1 output53 (.A(net53),
    .Z(read_data2[24]));
 BUF_X1 output54 (.A(net54),
    .Z(read_data2[25]));
 BUF_X1 output55 (.A(net55),
    .Z(read_data2[26]));
 BUF_X1 output56 (.A(net56),
    .Z(read_data2[27]));
 BUF_X1 output57 (.A(net57),
    .Z(read_data2[28]));
 BUF_X1 output58 (.A(net58),
    .Z(read_data2[29]));
 BUF_X1 output59 (.A(net59),
    .Z(read_data2[2]));
 BUF_X1 output60 (.A(net60),
    .Z(read_data2[30]));
 BUF_X1 output61 (.A(net61),
    .Z(read_data2[31]));
 BUF_X1 output62 (.A(net62),
    .Z(read_data2[3]));
 BUF_X1 output63 (.A(net63),
    .Z(read_data2[4]));
 BUF_X1 output64 (.A(net64),
    .Z(read_data2[5]));
 BUF_X1 output65 (.A(net65),
    .Z(read_data2[6]));
 BUF_X1 output66 (.A(net66),
    .Z(read_data2[7]));
 BUF_X1 output67 (.A(net67),
    .Z(read_data2[8]));
 BUF_X1 output68 (.A(net68),
    .Z(read_data2[9]));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_0_clk));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_43_clk));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_45_clk));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_47_clk));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_49_clk));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_51_clk));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_53_clk));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_55_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_58_clk));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_60_clk));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_62_clk));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_64_clk));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_66_clk));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_68_clk));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_70_clk));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_72_clk));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_74_clk));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_76_clk));
 CLKBUF_X3 clkbuf_leaf_77_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_77_clk));
 CLKBUF_X3 clkbuf_leaf_78_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_78_clk));
 CLKBUF_X3 clkbuf_leaf_79_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_79_clk));
 CLKBUF_X3 clkbuf_leaf_80_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_80_clk));
 CLKBUF_X3 clkbuf_leaf_81_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_81_clk));
 CLKBUF_X3 clkbuf_leaf_82_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_82_clk));
 CLKBUF_X3 clkbuf_leaf_83_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_83_clk));
 CLKBUF_X3 clkbuf_leaf_84_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_84_clk));
 CLKBUF_X3 clkbuf_leaf_85_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_85_clk));
 CLKBUF_X3 clkbuf_leaf_86_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_86_clk));
 CLKBUF_X3 clkbuf_leaf_87_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_87_clk));
 CLKBUF_X3 clkbuf_leaf_88_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_88_clk));
 CLKBUF_X3 clkbuf_leaf_89_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_89_clk));
 CLKBUF_X3 clkbuf_leaf_90_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_90_clk));
 CLKBUF_X3 clkbuf_leaf_91_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_91_clk));
 CLKBUF_X3 clkbuf_leaf_92_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_92_clk));
 CLKBUF_X3 clkbuf_leaf_93_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_93_clk));
 CLKBUF_X3 clkbuf_leaf_94_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_94_clk));
 CLKBUF_X3 clkbuf_leaf_95_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_95_clk));
 CLKBUF_X3 clkbuf_leaf_96_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_96_clk));
 CLKBUF_X3 clkbuf_leaf_97_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_97_clk));
 CLKBUF_X3 clkbuf_leaf_98_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_98_clk));
 CLKBUF_X3 clkbuf_leaf_99_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_99_clk));
 CLKBUF_X3 clkbuf_leaf_100_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_100_clk));
 CLKBUF_X3 clkbuf_leaf_101_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_101_clk));
 CLKBUF_X3 clkbuf_leaf_102_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_102_clk));
 CLKBUF_X3 clkbuf_leaf_103_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_103_clk));
 CLKBUF_X3 clkbuf_leaf_104_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_104_clk));
 CLKBUF_X3 clkbuf_leaf_105_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_105_clk));
 CLKBUF_X3 clkbuf_leaf_106_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_106_clk));
 CLKBUF_X3 clkbuf_leaf_107_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_107_clk));
 CLKBUF_X3 clkbuf_leaf_108_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_108_clk));
 CLKBUF_X3 clkbuf_leaf_109_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_109_clk));
 CLKBUF_X3 clkbuf_leaf_110_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_110_clk));
 CLKBUF_X3 clkbuf_leaf_111_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_111_clk));
 CLKBUF_X3 clkbuf_leaf_112_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_112_clk));
 CLKBUF_X3 clkbuf_leaf_113_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_113_clk));
 CLKBUF_X3 clkbuf_leaf_114_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_114_clk));
 CLKBUF_X3 clkbuf_leaf_115_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_115_clk));
 CLKBUF_X3 clkbuf_leaf_116_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_116_clk));
 CLKBUF_X3 clkbuf_leaf_117_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_117_clk));
 CLKBUF_X3 clkbuf_leaf_118_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_118_clk));
 CLKBUF_X3 clkbuf_leaf_119_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_119_clk));
 CLKBUF_X3 clkbuf_leaf_120_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_120_clk));
 CLKBUF_X3 clkbuf_leaf_121_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_121_clk));
 CLKBUF_X3 clkbuf_leaf_122_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_122_clk));
 CLKBUF_X3 clkbuf_leaf_123_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_123_clk));
 CLKBUF_X3 clkbuf_leaf_124_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_124_clk));
 CLKBUF_X3 clkbuf_leaf_125_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_125_clk));
 CLKBUF_X3 clkbuf_leaf_126_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_126_clk));
 CLKBUF_X3 clkbuf_leaf_127_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_127_clk));
 CLKBUF_X3 clkbuf_leaf_128_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_128_clk));
 CLKBUF_X3 clkbuf_leaf_129_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_129_clk));
 CLKBUF_X3 clkbuf_leaf_130_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_130_clk));
 CLKBUF_X3 clkbuf_leaf_131_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_131_clk));
 CLKBUF_X3 clkbuf_leaf_132_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_132_clk));
 CLKBUF_X3 clkbuf_leaf_133_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_133_clk));
 CLKBUF_X3 clkbuf_leaf_134_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_134_clk));
 CLKBUF_X3 clkbuf_leaf_135_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_135_clk));
 CLKBUF_X3 clkbuf_leaf_136_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_136_clk));
 CLKBUF_X3 clkbuf_leaf_137_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_137_clk));
 CLKBUF_X3 clkbuf_leaf_138_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_138_clk));
 CLKBUF_X3 clkbuf_leaf_139_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_139_clk));
 CLKBUF_X3 clkbuf_leaf_140_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_140_clk));
 CLKBUF_X3 clkbuf_leaf_141_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_141_clk));
 CLKBUF_X3 clkbuf_leaf_142_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_142_clk));
 CLKBUF_X3 clkbuf_leaf_143_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_143_clk));
 CLKBUF_X3 clkbuf_leaf_144_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_144_clk));
 CLKBUF_X3 clkbuf_leaf_145_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_145_clk));
 CLKBUF_X3 clkbuf_leaf_146_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_146_clk));
 CLKBUF_X3 clkbuf_leaf_147_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_147_clk));
 CLKBUF_X3 clkbuf_leaf_148_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_148_clk));
 CLKBUF_X3 clkbuf_leaf_149_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_149_clk));
 CLKBUF_X3 clkbuf_leaf_150_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_150_clk));
 CLKBUF_X3 clkbuf_leaf_151_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_151_clk));
 CLKBUF_X3 clkbuf_leaf_152_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_152_clk));
 CLKBUF_X3 clkbuf_leaf_153_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_153_clk));
 CLKBUF_X3 clkbuf_leaf_154_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_154_clk));
 CLKBUF_X3 clkbuf_leaf_155_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_155_clk));
 CLKBUF_X3 clkbuf_leaf_156_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_156_clk));
 CLKBUF_X3 clkbuf_leaf_157_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_157_clk));
 CLKBUF_X3 clkbuf_leaf_158_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_158_clk));
 CLKBUF_X3 clkbuf_leaf_159_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_159_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X2 clkload0 (.A(clknet_4_0_0_clk));
 INV_X2 clkload1 (.A(clknet_4_3_0_clk));
 INV_X2 clkload2 (.A(clknet_4_5_0_clk));
 INV_X2 clkload3 (.A(clknet_4_6_0_clk));
 CLKBUF_X3 clkload4 (.A(clknet_4_7_0_clk));
 CLKBUF_X3 clkload5 (.A(clknet_4_9_0_clk));
 CLKBUF_X3 clkload6 (.A(clknet_4_12_0_clk));
 CLKBUF_X3 clkload7 (.A(clknet_4_13_0_clk));
 CLKBUF_X3 clkload8 (.A(clknet_4_15_0_clk));
 INV_X1 clkload9 (.A(clknet_leaf_0_clk));
 INV_X1 clkload10 (.A(clknet_leaf_1_clk));
 CLKBUF_X1 clkload11 (.A(clknet_leaf_2_clk));
 INV_X1 clkload12 (.A(clknet_leaf_155_clk));
 INV_X1 clkload13 (.A(clknet_leaf_157_clk));
 INV_X1 clkload14 (.A(clknet_leaf_158_clk));
 INV_X2 clkload15 (.A(clknet_leaf_159_clk));
 CLKBUF_X1 clkload16 (.A(clknet_leaf_3_clk));
 CLKBUF_X1 clkload17 (.A(clknet_leaf_5_clk));
 INV_X1 clkload18 (.A(clknet_leaf_7_clk));
 CLKBUF_X1 clkload19 (.A(clknet_leaf_9_clk));
 INV_X1 clkload20 (.A(clknet_leaf_10_clk));
 CLKBUF_X1 clkload21 (.A(clknet_leaf_11_clk));
 INV_X1 clkload22 (.A(clknet_leaf_12_clk));
 CLKBUF_X1 clkload23 (.A(clknet_leaf_14_clk));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_144_clk));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_145_clk));
 CLKBUF_X1 clkload26 (.A(clknet_leaf_146_clk));
 INV_X2 clkload27 (.A(clknet_leaf_147_clk));
 CLKBUF_X1 clkload28 (.A(clknet_leaf_148_clk));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_150_clk));
 CLKBUF_X1 clkload30 (.A(clknet_leaf_151_clk));
 CLKBUF_X1 clkload31 (.A(clknet_leaf_152_clk));
 INV_X1 clkload32 (.A(clknet_leaf_153_clk));
 INV_X1 clkload33 (.A(clknet_leaf_154_clk));
 CLKBUF_X1 clkload34 (.A(clknet_leaf_15_clk));
 CLKBUF_X1 clkload35 (.A(clknet_leaf_16_clk));
 CLKBUF_X1 clkload36 (.A(clknet_leaf_17_clk));
 CLKBUF_X1 clkload37 (.A(clknet_leaf_19_clk));
 CLKBUF_X1 clkload38 (.A(clknet_leaf_22_clk));
 CLKBUF_X1 clkload39 (.A(clknet_leaf_23_clk));
 INV_X1 clkload40 (.A(clknet_leaf_24_clk));
 INV_X1 clkload41 (.A(clknet_leaf_25_clk));
 CLKBUF_X1 clkload42 (.A(clknet_leaf_26_clk));
 INV_X1 clkload43 (.A(clknet_leaf_28_clk));
 INV_X1 clkload44 (.A(clknet_leaf_30_clk));
 INV_X1 clkload45 (.A(clknet_leaf_31_clk));
 CLKBUF_X1 clkload46 (.A(clknet_leaf_34_clk));
 CLKBUF_X1 clkload47 (.A(clknet_leaf_36_clk));
 CLKBUF_X1 clkload48 (.A(clknet_leaf_37_clk));
 CLKBUF_X1 clkload49 (.A(clknet_leaf_18_clk));
 CLKBUF_X1 clkload50 (.A(clknet_leaf_21_clk));
 CLKBUF_X1 clkload51 (.A(clknet_leaf_51_clk));
 CLKBUF_X1 clkload52 (.A(clknet_leaf_52_clk));
 CLKBUF_X1 clkload53 (.A(clknet_leaf_53_clk));
 INV_X1 clkload54 (.A(clknet_leaf_54_clk));
 CLKBUF_X1 clkload55 (.A(clknet_leaf_55_clk));
 CLKBUF_X1 clkload56 (.A(clknet_leaf_41_clk));
 INV_X1 clkload57 (.A(clknet_leaf_42_clk));
 INV_X1 clkload58 (.A(clknet_leaf_43_clk));
 CLKBUF_X1 clkload59 (.A(clknet_leaf_45_clk));
 CLKBUF_X1 clkload60 (.A(clknet_leaf_46_clk));
 CLKBUF_X1 clkload61 (.A(clknet_leaf_47_clk));
 INV_X1 clkload62 (.A(clknet_leaf_48_clk));
 CLKBUF_X1 clkload63 (.A(clknet_leaf_49_clk));
 INV_X1 clkload64 (.A(clknet_leaf_50_clk));
 INV_X1 clkload65 (.A(clknet_leaf_123_clk));
 INV_X1 clkload66 (.A(clknet_leaf_124_clk));
 CLKBUF_X1 clkload67 (.A(clknet_leaf_125_clk));
 INV_X1 clkload68 (.A(clknet_leaf_126_clk));
 CLKBUF_X1 clkload69 (.A(clknet_leaf_127_clk));
 CLKBUF_X1 clkload70 (.A(clknet_leaf_128_clk));
 CLKBUF_X1 clkload71 (.A(clknet_leaf_130_clk));
 CLKBUF_X1 clkload72 (.A(clknet_leaf_131_clk));
 INV_X1 clkload73 (.A(clknet_leaf_132_clk));
 CLKBUF_X1 clkload74 (.A(clknet_leaf_133_clk));
 CLKBUF_X1 clkload75 (.A(clknet_leaf_99_clk));
 CLKBUF_X1 clkload76 (.A(clknet_leaf_100_clk));
 CLKBUF_X1 clkload77 (.A(clknet_leaf_134_clk));
 CLKBUF_X1 clkload78 (.A(clknet_leaf_136_clk));
 CLKBUF_X1 clkload79 (.A(clknet_leaf_137_clk));
 CLKBUF_X1 clkload80 (.A(clknet_leaf_139_clk));
 CLKBUF_X1 clkload81 (.A(clknet_leaf_112_clk));
 CLKBUF_X1 clkload82 (.A(clknet_leaf_114_clk));
 CLKBUF_X1 clkload83 (.A(clknet_leaf_115_clk));
 CLKBUF_X1 clkload84 (.A(clknet_leaf_116_clk));
 INV_X1 clkload85 (.A(clknet_leaf_117_clk));
 CLKBUF_X1 clkload86 (.A(clknet_leaf_119_clk));
 CLKBUF_X1 clkload87 (.A(clknet_leaf_120_clk));
 INV_X1 clkload88 (.A(clknet_leaf_121_clk));
 CLKBUF_X1 clkload89 (.A(clknet_leaf_122_clk));
 CLKBUF_X1 clkload90 (.A(clknet_leaf_101_clk));
 CLKBUF_X1 clkload91 (.A(clknet_leaf_103_clk));
 INV_X1 clkload92 (.A(clknet_leaf_104_clk));
 CLKBUF_X1 clkload93 (.A(clknet_leaf_105_clk));
 INV_X1 clkload94 (.A(clknet_leaf_106_clk));
 INV_X1 clkload95 (.A(clknet_leaf_108_clk));
 CLKBUF_X1 clkload96 (.A(clknet_leaf_109_clk));
 CLKBUF_X1 clkload97 (.A(clknet_leaf_110_clk));
 CLKBUF_X1 clkload98 (.A(clknet_leaf_111_clk));
 CLKBUF_X1 clkload99 (.A(clknet_leaf_56_clk));
 CLKBUF_X1 clkload100 (.A(clknet_leaf_58_clk));
 CLKBUF_X1 clkload101 (.A(clknet_leaf_59_clk));
 CLKBUF_X1 clkload102 (.A(clknet_leaf_60_clk));
 CLKBUF_X1 clkload103 (.A(clknet_leaf_92_clk));
 INV_X1 clkload104 (.A(clknet_leaf_93_clk));
 CLKBUF_X1 clkload105 (.A(clknet_leaf_94_clk));
 CLKBUF_X1 clkload106 (.A(clknet_leaf_95_clk));
 CLKBUF_X1 clkload107 (.A(clknet_leaf_96_clk));
 INV_X1 clkload108 (.A(clknet_leaf_61_clk));
 CLKBUF_X1 clkload109 (.A(clknet_leaf_62_clk));
 CLKBUF_X1 clkload110 (.A(clknet_leaf_64_clk));
 CLKBUF_X1 clkload111 (.A(clknet_leaf_65_clk));
 CLKBUF_X1 clkload112 (.A(clknet_leaf_66_clk));
 CLKBUF_X1 clkload113 (.A(clknet_leaf_67_clk));
 CLKBUF_X1 clkload114 (.A(clknet_leaf_69_clk));
 INV_X1 clkload115 (.A(clknet_leaf_70_clk));
 CLKBUF_X1 clkload116 (.A(clknet_leaf_81_clk));
 CLKBUF_X1 clkload117 (.A(clknet_leaf_82_clk));
 CLKBUF_X1 clkload118 (.A(clknet_leaf_87_clk));
 CLKBUF_X1 clkload119 (.A(clknet_leaf_89_clk));
 CLKBUF_X1 clkload120 (.A(clknet_leaf_90_clk));
 CLKBUF_X1 clkload121 (.A(clknet_leaf_91_clk));
 INV_X1 clkload122 (.A(clknet_leaf_71_clk));
 CLKBUF_X1 clkload123 (.A(clknet_leaf_72_clk));
 CLKBUF_X1 clkload124 (.A(clknet_leaf_73_clk));
 INV_X1 clkload125 (.A(clknet_leaf_74_clk));
 CLKBUF_X1 clkload126 (.A(clknet_leaf_75_clk));
 CLKBUF_X1 clkload127 (.A(clknet_leaf_76_clk));
 CLKBUF_X1 clkload128 (.A(clknet_leaf_79_clk));
 CLKBUF_X1 clkload129 (.A(clknet_leaf_80_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X8 FILLER_0_225 ();
 FILLCELL_X1 FILLER_0_233 ();
 FILLCELL_X16 FILLER_0_239 ();
 FILLCELL_X8 FILLER_0_255 ();
 FILLCELL_X4 FILLER_0_263 ();
 FILLCELL_X1 FILLER_0_267 ();
 FILLCELL_X4 FILLER_0_275 ();
 FILLCELL_X1 FILLER_0_279 ();
 FILLCELL_X2 FILLER_0_288 ();
 FILLCELL_X1 FILLER_0_290 ();
 FILLCELL_X8 FILLER_0_300 ();
 FILLCELL_X1 FILLER_0_315 ();
 FILLCELL_X4 FILLER_0_328 ();
 FILLCELL_X4 FILLER_0_354 ();
 FILLCELL_X2 FILLER_0_358 ();
 FILLCELL_X4 FILLER_0_364 ();
 FILLCELL_X2 FILLER_0_368 ();
 FILLCELL_X1 FILLER_0_373 ();
 FILLCELL_X8 FILLER_0_391 ();
 FILLCELL_X16 FILLER_0_412 ();
 FILLCELL_X8 FILLER_0_428 ();
 FILLCELL_X2 FILLER_0_436 ();
 FILLCELL_X2 FILLER_0_455 ();
 FILLCELL_X4 FILLER_0_474 ();
 FILLCELL_X2 FILLER_0_478 ();
 FILLCELL_X1 FILLER_0_480 ();
 FILLCELL_X32 FILLER_0_498 ();
 FILLCELL_X32 FILLER_0_530 ();
 FILLCELL_X32 FILLER_0_562 ();
 FILLCELL_X32 FILLER_0_594 ();
 FILLCELL_X4 FILLER_0_626 ();
 FILLCELL_X1 FILLER_0_630 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X16 FILLER_0_792 ();
 FILLCELL_X4 FILLER_0_808 ();
 FILLCELL_X2 FILLER_0_812 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X4 FILLER_1_225 ();
 FILLCELL_X1 FILLER_1_229 ();
 FILLCELL_X16 FILLER_1_237 ();
 FILLCELL_X1 FILLER_1_253 ();
 FILLCELL_X1 FILLER_1_278 ();
 FILLCELL_X4 FILLER_1_282 ();
 FILLCELL_X1 FILLER_1_286 ();
 FILLCELL_X4 FILLER_1_307 ();
 FILLCELL_X1 FILLER_1_311 ();
 FILLCELL_X8 FILLER_1_329 ();
 FILLCELL_X4 FILLER_1_337 ();
 FILLCELL_X2 FILLER_1_341 ();
 FILLCELL_X8 FILLER_1_348 ();
 FILLCELL_X2 FILLER_1_356 ();
 FILLCELL_X2 FILLER_1_375 ();
 FILLCELL_X16 FILLER_1_384 ();
 FILLCELL_X4 FILLER_1_400 ();
 FILLCELL_X1 FILLER_1_404 ();
 FILLCELL_X16 FILLER_1_422 ();
 FILLCELL_X8 FILLER_1_438 ();
 FILLCELL_X1 FILLER_1_446 ();
 FILLCELL_X4 FILLER_1_454 ();
 FILLCELL_X1 FILLER_1_458 ();
 FILLCELL_X4 FILLER_1_463 ();
 FILLCELL_X2 FILLER_1_467 ();
 FILLCELL_X2 FILLER_1_472 ();
 FILLCELL_X1 FILLER_1_474 ();
 FILLCELL_X4 FILLER_1_480 ();
 FILLCELL_X2 FILLER_1_484 ();
 FILLCELL_X1 FILLER_1_486 ();
 FILLCELL_X4 FILLER_1_491 ();
 FILLCELL_X2 FILLER_1_495 ();
 FILLCELL_X1 FILLER_1_497 ();
 FILLCELL_X32 FILLER_1_549 ();
 FILLCELL_X32 FILLER_1_581 ();
 FILLCELL_X32 FILLER_1_613 ();
 FILLCELL_X32 FILLER_1_645 ();
 FILLCELL_X32 FILLER_1_677 ();
 FILLCELL_X32 FILLER_1_709 ();
 FILLCELL_X32 FILLER_1_741 ();
 FILLCELL_X32 FILLER_1_773 ();
 FILLCELL_X8 FILLER_1_805 ();
 FILLCELL_X1 FILLER_1_813 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X4 FILLER_2_225 ();
 FILLCELL_X2 FILLER_2_229 ();
 FILLCELL_X1 FILLER_2_231 ();
 FILLCELL_X4 FILLER_2_237 ();
 FILLCELL_X2 FILLER_2_241 ();
 FILLCELL_X1 FILLER_2_243 ();
 FILLCELL_X16 FILLER_2_251 ();
 FILLCELL_X16 FILLER_2_274 ();
 FILLCELL_X2 FILLER_2_290 ();
 FILLCELL_X32 FILLER_2_299 ();
 FILLCELL_X1 FILLER_2_331 ();
 FILLCELL_X1 FILLER_2_351 ();
 FILLCELL_X2 FILLER_2_367 ();
 FILLCELL_X1 FILLER_2_372 ();
 FILLCELL_X4 FILLER_2_390 ();
 FILLCELL_X2 FILLER_2_394 ();
 FILLCELL_X1 FILLER_2_406 ();
 FILLCELL_X32 FILLER_2_414 ();
 FILLCELL_X2 FILLER_2_446 ();
 FILLCELL_X2 FILLER_2_451 ();
 FILLCELL_X1 FILLER_2_453 ();
 FILLCELL_X1 FILLER_2_460 ();
 FILLCELL_X8 FILLER_2_488 ();
 FILLCELL_X1 FILLER_2_496 ();
 FILLCELL_X1 FILLER_2_528 ();
 FILLCELL_X1 FILLER_2_539 ();
 FILLCELL_X8 FILLER_2_543 ();
 FILLCELL_X8 FILLER_2_568 ();
 FILLCELL_X32 FILLER_2_593 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X16 FILLER_2_792 ();
 FILLCELL_X4 FILLER_2_808 ();
 FILLCELL_X2 FILLER_2_812 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X8 FILLER_3_225 ();
 FILLCELL_X4 FILLER_3_233 ();
 FILLCELL_X2 FILLER_3_237 ();
 FILLCELL_X1 FILLER_3_259 ();
 FILLCELL_X1 FILLER_3_284 ();
 FILLCELL_X2 FILLER_3_292 ();
 FILLCELL_X1 FILLER_3_294 ();
 FILLCELL_X2 FILLER_3_302 ();
 FILLCELL_X2 FILLER_3_321 ();
 FILLCELL_X1 FILLER_3_323 ();
 FILLCELL_X1 FILLER_3_341 ();
 FILLCELL_X4 FILLER_3_345 ();
 FILLCELL_X1 FILLER_3_349 ();
 FILLCELL_X2 FILLER_3_372 ();
 FILLCELL_X2 FILLER_3_378 ();
 FILLCELL_X4 FILLER_3_383 ();
 FILLCELL_X2 FILLER_3_387 ();
 FILLCELL_X1 FILLER_3_389 ();
 FILLCELL_X8 FILLER_3_414 ();
 FILLCELL_X4 FILLER_3_422 ();
 FILLCELL_X1 FILLER_3_426 ();
 FILLCELL_X16 FILLER_3_444 ();
 FILLCELL_X8 FILLER_3_460 ();
 FILLCELL_X8 FILLER_3_488 ();
 FILLCELL_X4 FILLER_3_496 ();
 FILLCELL_X1 FILLER_3_500 ();
 FILLCELL_X8 FILLER_3_504 ();
 FILLCELL_X4 FILLER_3_512 ();
 FILLCELL_X2 FILLER_3_516 ();
 FILLCELL_X1 FILLER_3_518 ();
 FILLCELL_X16 FILLER_3_532 ();
 FILLCELL_X2 FILLER_3_548 ();
 FILLCELL_X1 FILLER_3_550 ();
 FILLCELL_X4 FILLER_3_575 ();
 FILLCELL_X2 FILLER_3_579 ();
 FILLCELL_X4 FILLER_3_589 ();
 FILLCELL_X2 FILLER_3_593 ();
 FILLCELL_X32 FILLER_3_616 ();
 FILLCELL_X16 FILLER_3_652 ();
 FILLCELL_X8 FILLER_3_668 ();
 FILLCELL_X2 FILLER_3_676 ();
 FILLCELL_X1 FILLER_3_682 ();
 FILLCELL_X1 FILLER_3_687 ();
 FILLCELL_X16 FILLER_3_692 ();
 FILLCELL_X1 FILLER_3_708 ();
 FILLCELL_X8 FILLER_3_726 ();
 FILLCELL_X2 FILLER_3_734 ();
 FILLCELL_X1 FILLER_3_736 ();
 FILLCELL_X32 FILLER_3_744 ();
 FILLCELL_X32 FILLER_3_776 ();
 FILLCELL_X4 FILLER_3_808 ();
 FILLCELL_X2 FILLER_3_812 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X16 FILLER_4_225 ();
 FILLCELL_X4 FILLER_4_241 ();
 FILLCELL_X4 FILLER_4_248 ();
 FILLCELL_X1 FILLER_4_252 ();
 FILLCELL_X8 FILLER_4_258 ();
 FILLCELL_X4 FILLER_4_266 ();
 FILLCELL_X2 FILLER_4_302 ();
 FILLCELL_X1 FILLER_4_304 ();
 FILLCELL_X2 FILLER_4_312 ();
 FILLCELL_X8 FILLER_4_324 ();
 FILLCELL_X8 FILLER_4_342 ();
 FILLCELL_X4 FILLER_4_355 ();
 FILLCELL_X2 FILLER_4_359 ();
 FILLCELL_X8 FILLER_4_368 ();
 FILLCELL_X2 FILLER_4_376 ();
 FILLCELL_X8 FILLER_4_383 ();
 FILLCELL_X2 FILLER_4_391 ();
 FILLCELL_X1 FILLER_4_393 ();
 FILLCELL_X8 FILLER_4_397 ();
 FILLCELL_X4 FILLER_4_425 ();
 FILLCELL_X1 FILLER_4_436 ();
 FILLCELL_X8 FILLER_4_444 ();
 FILLCELL_X1 FILLER_4_452 ();
 FILLCELL_X2 FILLER_4_457 ();
 FILLCELL_X2 FILLER_4_462 ();
 FILLCELL_X1 FILLER_4_474 ();
 FILLCELL_X8 FILLER_4_495 ();
 FILLCELL_X4 FILLER_4_503 ();
 FILLCELL_X2 FILLER_4_507 ();
 FILLCELL_X32 FILLER_4_516 ();
 FILLCELL_X8 FILLER_4_548 ();
 FILLCELL_X1 FILLER_4_556 ();
 FILLCELL_X16 FILLER_4_574 ();
 FILLCELL_X8 FILLER_4_619 ();
 FILLCELL_X4 FILLER_4_627 ();
 FILLCELL_X4 FILLER_4_632 ();
 FILLCELL_X2 FILLER_4_636 ();
 FILLCELL_X1 FILLER_4_638 ();
 FILLCELL_X16 FILLER_4_694 ();
 FILLCELL_X4 FILLER_4_710 ();
 FILLCELL_X1 FILLER_4_714 ();
 FILLCELL_X1 FILLER_4_725 ();
 FILLCELL_X1 FILLER_4_732 ();
 FILLCELL_X32 FILLER_4_750 ();
 FILLCELL_X32 FILLER_4_782 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X8 FILLER_5_161 ();
 FILLCELL_X4 FILLER_5_169 ();
 FILLCELL_X2 FILLER_5_173 ();
 FILLCELL_X1 FILLER_5_175 ();
 FILLCELL_X4 FILLER_5_193 ();
 FILLCELL_X16 FILLER_5_214 ();
 FILLCELL_X8 FILLER_5_230 ();
 FILLCELL_X4 FILLER_5_238 ();
 FILLCELL_X1 FILLER_5_242 ();
 FILLCELL_X8 FILLER_5_247 ();
 FILLCELL_X1 FILLER_5_255 ();
 FILLCELL_X1 FILLER_5_259 ();
 FILLCELL_X1 FILLER_5_265 ();
 FILLCELL_X8 FILLER_5_301 ();
 FILLCELL_X4 FILLER_5_329 ();
 FILLCELL_X1 FILLER_5_333 ();
 FILLCELL_X16 FILLER_5_341 ();
 FILLCELL_X4 FILLER_5_357 ();
 FILLCELL_X4 FILLER_5_378 ();
 FILLCELL_X2 FILLER_5_389 ();
 FILLCELL_X1 FILLER_5_391 ();
 FILLCELL_X2 FILLER_5_399 ();
 FILLCELL_X8 FILLER_5_408 ();
 FILLCELL_X4 FILLER_5_416 ();
 FILLCELL_X2 FILLER_5_420 ();
 FILLCELL_X1 FILLER_5_422 ();
 FILLCELL_X2 FILLER_5_433 ();
 FILLCELL_X4 FILLER_5_469 ();
 FILLCELL_X2 FILLER_5_473 ();
 FILLCELL_X1 FILLER_5_475 ();
 FILLCELL_X8 FILLER_5_483 ();
 FILLCELL_X1 FILLER_5_491 ();
 FILLCELL_X1 FILLER_5_499 ();
 FILLCELL_X1 FILLER_5_507 ();
 FILLCELL_X2 FILLER_5_515 ();
 FILLCELL_X4 FILLER_5_531 ();
 FILLCELL_X1 FILLER_5_535 ();
 FILLCELL_X4 FILLER_5_557 ();
 FILLCELL_X1 FILLER_5_561 ();
 FILLCELL_X4 FILLER_5_579 ();
 FILLCELL_X8 FILLER_5_600 ();
 FILLCELL_X2 FILLER_5_608 ();
 FILLCELL_X1 FILLER_5_610 ();
 FILLCELL_X16 FILLER_5_628 ();
 FILLCELL_X1 FILLER_5_644 ();
 FILLCELL_X1 FILLER_5_657 ();
 FILLCELL_X4 FILLER_5_662 ();
 FILLCELL_X16 FILLER_5_670 ();
 FILLCELL_X2 FILLER_5_686 ();
 FILLCELL_X4 FILLER_5_729 ();
 FILLCELL_X2 FILLER_5_733 ();
 FILLCELL_X32 FILLER_5_755 ();
 FILLCELL_X16 FILLER_5_787 ();
 FILLCELL_X8 FILLER_5_803 ();
 FILLCELL_X2 FILLER_5_811 ();
 FILLCELL_X1 FILLER_5_813 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X16 FILLER_6_129 ();
 FILLCELL_X16 FILLER_6_148 ();
 FILLCELL_X8 FILLER_6_164 ();
 FILLCELL_X4 FILLER_6_172 ();
 FILLCELL_X2 FILLER_6_176 ();
 FILLCELL_X1 FILLER_6_178 ();
 FILLCELL_X8 FILLER_6_189 ();
 FILLCELL_X16 FILLER_6_207 ();
 FILLCELL_X1 FILLER_6_223 ();
 FILLCELL_X4 FILLER_6_229 ();
 FILLCELL_X2 FILLER_6_238 ();
 FILLCELL_X16 FILLER_6_274 ();
 FILLCELL_X4 FILLER_6_297 ();
 FILLCELL_X2 FILLER_6_315 ();
 FILLCELL_X2 FILLER_6_336 ();
 FILLCELL_X1 FILLER_6_338 ();
 FILLCELL_X2 FILLER_6_356 ();
 FILLCELL_X4 FILLER_6_375 ();
 FILLCELL_X2 FILLER_6_379 ();
 FILLCELL_X2 FILLER_6_388 ();
 FILLCELL_X4 FILLER_6_411 ();
 FILLCELL_X2 FILLER_6_415 ();
 FILLCELL_X1 FILLER_6_417 ();
 FILLCELL_X4 FILLER_6_446 ();
 FILLCELL_X2 FILLER_6_450 ();
 FILLCELL_X4 FILLER_6_455 ();
 FILLCELL_X1 FILLER_6_459 ();
 FILLCELL_X8 FILLER_6_463 ();
 FILLCELL_X2 FILLER_6_475 ();
 FILLCELL_X1 FILLER_6_477 ();
 FILLCELL_X8 FILLER_6_481 ();
 FILLCELL_X1 FILLER_6_489 ();
 FILLCELL_X4 FILLER_6_504 ();
 FILLCELL_X2 FILLER_6_508 ();
 FILLCELL_X1 FILLER_6_510 ();
 FILLCELL_X1 FILLER_6_520 ();
 FILLCELL_X4 FILLER_6_526 ();
 FILLCELL_X2 FILLER_6_530 ();
 FILLCELL_X1 FILLER_6_532 ();
 FILLCELL_X8 FILLER_6_545 ();
 FILLCELL_X4 FILLER_6_553 ();
 FILLCELL_X2 FILLER_6_557 ();
 FILLCELL_X4 FILLER_6_564 ();
 FILLCELL_X1 FILLER_6_568 ();
 FILLCELL_X8 FILLER_6_577 ();
 FILLCELL_X2 FILLER_6_585 ();
 FILLCELL_X1 FILLER_6_587 ();
 FILLCELL_X4 FILLER_6_596 ();
 FILLCELL_X2 FILLER_6_600 ();
 FILLCELL_X8 FILLER_6_617 ();
 FILLCELL_X2 FILLER_6_625 ();
 FILLCELL_X1 FILLER_6_627 ();
 FILLCELL_X4 FILLER_6_637 ();
 FILLCELL_X1 FILLER_6_662 ();
 FILLCELL_X8 FILLER_6_674 ();
 FILLCELL_X1 FILLER_6_682 ();
 FILLCELL_X2 FILLER_6_687 ();
 FILLCELL_X1 FILLER_6_689 ();
 FILLCELL_X8 FILLER_6_699 ();
 FILLCELL_X2 FILLER_6_707 ();
 FILLCELL_X8 FILLER_6_729 ();
 FILLCELL_X1 FILLER_6_737 ();
 FILLCELL_X8 FILLER_6_745 ();
 FILLCELL_X4 FILLER_6_753 ();
 FILLCELL_X2 FILLER_6_757 ();
 FILLCELL_X32 FILLER_6_761 ();
 FILLCELL_X16 FILLER_6_793 ();
 FILLCELL_X4 FILLER_6_809 ();
 FILLCELL_X1 FILLER_6_813 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X8 FILLER_7_129 ();
 FILLCELL_X4 FILLER_7_137 ();
 FILLCELL_X2 FILLER_7_141 ();
 FILLCELL_X1 FILLER_7_143 ();
 FILLCELL_X8 FILLER_7_151 ();
 FILLCELL_X4 FILLER_7_159 ();
 FILLCELL_X2 FILLER_7_163 ();
 FILLCELL_X4 FILLER_7_169 ();
 FILLCELL_X1 FILLER_7_173 ();
 FILLCELL_X8 FILLER_7_191 ();
 FILLCELL_X4 FILLER_7_199 ();
 FILLCELL_X2 FILLER_7_203 ();
 FILLCELL_X8 FILLER_7_229 ();
 FILLCELL_X4 FILLER_7_237 ();
 FILLCELL_X1 FILLER_7_241 ();
 FILLCELL_X4 FILLER_7_254 ();
 FILLCELL_X1 FILLER_7_258 ();
 FILLCELL_X4 FILLER_7_262 ();
 FILLCELL_X2 FILLER_7_266 ();
 FILLCELL_X2 FILLER_7_278 ();
 FILLCELL_X2 FILLER_7_283 ();
 FILLCELL_X1 FILLER_7_319 ();
 FILLCELL_X2 FILLER_7_330 ();
 FILLCELL_X1 FILLER_7_332 ();
 FILLCELL_X2 FILLER_7_340 ();
 FILLCELL_X2 FILLER_7_345 ();
 FILLCELL_X1 FILLER_7_347 ();
 FILLCELL_X4 FILLER_7_353 ();
 FILLCELL_X1 FILLER_7_357 ();
 FILLCELL_X1 FILLER_7_375 ();
 FILLCELL_X8 FILLER_7_414 ();
 FILLCELL_X2 FILLER_7_422 ();
 FILLCELL_X32 FILLER_7_427 ();
 FILLCELL_X4 FILLER_7_459 ();
 FILLCELL_X2 FILLER_7_466 ();
 FILLCELL_X1 FILLER_7_468 ();
 FILLCELL_X4 FILLER_7_486 ();
 FILLCELL_X1 FILLER_7_490 ();
 FILLCELL_X2 FILLER_7_512 ();
 FILLCELL_X1 FILLER_7_514 ();
 FILLCELL_X2 FILLER_7_524 ();
 FILLCELL_X1 FILLER_7_526 ();
 FILLCELL_X16 FILLER_7_549 ();
 FILLCELL_X4 FILLER_7_565 ();
 FILLCELL_X16 FILLER_7_583 ();
 FILLCELL_X1 FILLER_7_599 ();
 FILLCELL_X2 FILLER_7_607 ();
 FILLCELL_X16 FILLER_7_626 ();
 FILLCELL_X2 FILLER_7_642 ();
 FILLCELL_X1 FILLER_7_644 ();
 FILLCELL_X1 FILLER_7_653 ();
 FILLCELL_X4 FILLER_7_676 ();
 FILLCELL_X8 FILLER_7_705 ();
 FILLCELL_X1 FILLER_7_713 ();
 FILLCELL_X4 FILLER_7_721 ();
 FILLCELL_X8 FILLER_7_732 ();
 FILLCELL_X4 FILLER_7_740 ();
 FILLCELL_X2 FILLER_7_744 ();
 FILLCELL_X1 FILLER_7_746 ();
 FILLCELL_X1 FILLER_7_751 ();
 FILLCELL_X32 FILLER_7_774 ();
 FILLCELL_X8 FILLER_7_806 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X16 FILLER_8_97 ();
 FILLCELL_X8 FILLER_8_113 ();
 FILLCELL_X4 FILLER_8_121 ();
 FILLCELL_X2 FILLER_8_125 ();
 FILLCELL_X4 FILLER_8_152 ();
 FILLCELL_X4 FILLER_8_181 ();
 FILLCELL_X2 FILLER_8_185 ();
 FILLCELL_X1 FILLER_8_187 ();
 FILLCELL_X1 FILLER_8_192 ();
 FILLCELL_X8 FILLER_8_198 ();
 FILLCELL_X2 FILLER_8_206 ();
 FILLCELL_X4 FILLER_8_211 ();
 FILLCELL_X1 FILLER_8_215 ();
 FILLCELL_X2 FILLER_8_240 ();
 FILLCELL_X4 FILLER_8_259 ();
 FILLCELL_X1 FILLER_8_263 ();
 FILLCELL_X8 FILLER_8_281 ();
 FILLCELL_X1 FILLER_8_289 ();
 FILLCELL_X4 FILLER_8_293 ();
 FILLCELL_X2 FILLER_8_297 ();
 FILLCELL_X1 FILLER_8_299 ();
 FILLCELL_X2 FILLER_8_338 ();
 FILLCELL_X1 FILLER_8_340 ();
 FILLCELL_X16 FILLER_8_345 ();
 FILLCELL_X1 FILLER_8_361 ();
 FILLCELL_X16 FILLER_8_372 ();
 FILLCELL_X4 FILLER_8_388 ();
 FILLCELL_X2 FILLER_8_392 ();
 FILLCELL_X16 FILLER_8_408 ();
 FILLCELL_X4 FILLER_8_424 ();
 FILLCELL_X2 FILLER_8_428 ();
 FILLCELL_X8 FILLER_8_437 ();
 FILLCELL_X4 FILLER_8_445 ();
 FILLCELL_X2 FILLER_8_466 ();
 FILLCELL_X4 FILLER_8_485 ();
 FILLCELL_X1 FILLER_8_489 ();
 FILLCELL_X1 FILLER_8_505 ();
 FILLCELL_X4 FILLER_8_526 ();
 FILLCELL_X2 FILLER_8_530 ();
 FILLCELL_X1 FILLER_8_547 ();
 FILLCELL_X1 FILLER_8_554 ();
 FILLCELL_X4 FILLER_8_582 ();
 FILLCELL_X1 FILLER_8_586 ();
 FILLCELL_X8 FILLER_8_623 ();
 FILLCELL_X16 FILLER_8_653 ();
 FILLCELL_X8 FILLER_8_676 ();
 FILLCELL_X4 FILLER_8_684 ();
 FILLCELL_X2 FILLER_8_688 ();
 FILLCELL_X4 FILLER_8_707 ();
 FILLCELL_X1 FILLER_8_725 ();
 FILLCELL_X8 FILLER_8_733 ();
 FILLCELL_X32 FILLER_8_775 ();
 FILLCELL_X4 FILLER_8_807 ();
 FILLCELL_X2 FILLER_8_811 ();
 FILLCELL_X1 FILLER_8_813 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X16 FILLER_9_97 ();
 FILLCELL_X8 FILLER_9_113 ();
 FILLCELL_X1 FILLER_9_121 ();
 FILLCELL_X8 FILLER_9_139 ();
 FILLCELL_X2 FILLER_9_147 ();
 FILLCELL_X16 FILLER_9_166 ();
 FILLCELL_X1 FILLER_9_198 ();
 FILLCELL_X8 FILLER_9_216 ();
 FILLCELL_X2 FILLER_9_224 ();
 FILLCELL_X4 FILLER_9_240 ();
 FILLCELL_X1 FILLER_9_244 ();
 FILLCELL_X1 FILLER_9_248 ();
 FILLCELL_X8 FILLER_9_252 ();
 FILLCELL_X4 FILLER_9_260 ();
 FILLCELL_X2 FILLER_9_264 ();
 FILLCELL_X4 FILLER_9_276 ();
 FILLCELL_X4 FILLER_9_301 ();
 FILLCELL_X1 FILLER_9_305 ();
 FILLCELL_X16 FILLER_9_313 ();
 FILLCELL_X8 FILLER_9_329 ();
 FILLCELL_X2 FILLER_9_337 ();
 FILLCELL_X1 FILLER_9_359 ();
 FILLCELL_X1 FILLER_9_377 ();
 FILLCELL_X1 FILLER_9_385 ();
 FILLCELL_X1 FILLER_9_393 ();
 FILLCELL_X16 FILLER_9_408 ();
 FILLCELL_X1 FILLER_9_424 ();
 FILLCELL_X1 FILLER_9_466 ();
 FILLCELL_X2 FILLER_9_470 ();
 FILLCELL_X8 FILLER_9_479 ();
 FILLCELL_X1 FILLER_9_487 ();
 FILLCELL_X4 FILLER_9_523 ();
 FILLCELL_X8 FILLER_9_531 ();
 FILLCELL_X2 FILLER_9_546 ();
 FILLCELL_X1 FILLER_9_548 ();
 FILLCELL_X4 FILLER_9_551 ();
 FILLCELL_X1 FILLER_9_555 ();
 FILLCELL_X8 FILLER_9_565 ();
 FILLCELL_X4 FILLER_9_573 ();
 FILLCELL_X2 FILLER_9_581 ();
 FILLCELL_X2 FILLER_9_585 ();
 FILLCELL_X8 FILLER_9_589 ();
 FILLCELL_X2 FILLER_9_597 ();
 FILLCELL_X2 FILLER_9_601 ();
 FILLCELL_X1 FILLER_9_603 ();
 FILLCELL_X16 FILLER_9_610 ();
 FILLCELL_X8 FILLER_9_626 ();
 FILLCELL_X2 FILLER_9_634 ();
 FILLCELL_X1 FILLER_9_636 ();
 FILLCELL_X4 FILLER_9_665 ();
 FILLCELL_X2 FILLER_9_669 ();
 FILLCELL_X1 FILLER_9_682 ();
 FILLCELL_X8 FILLER_9_687 ();
 FILLCELL_X16 FILLER_9_702 ();
 FILLCELL_X4 FILLER_9_718 ();
 FILLCELL_X2 FILLER_9_722 ();
 FILLCELL_X1 FILLER_9_724 ();
 FILLCELL_X16 FILLER_9_732 ();
 FILLCELL_X1 FILLER_9_748 ();
 FILLCELL_X4 FILLER_9_752 ();
 FILLCELL_X1 FILLER_9_756 ();
 FILLCELL_X1 FILLER_9_767 ();
 FILLCELL_X2 FILLER_9_771 ();
 FILLCELL_X16 FILLER_9_790 ();
 FILLCELL_X8 FILLER_9_806 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X16 FILLER_10_129 ();
 FILLCELL_X8 FILLER_10_145 ();
 FILLCELL_X4 FILLER_10_153 ();
 FILLCELL_X1 FILLER_10_157 ();
 FILLCELL_X4 FILLER_10_166 ();
 FILLCELL_X2 FILLER_10_170 ();
 FILLCELL_X1 FILLER_10_179 ();
 FILLCELL_X1 FILLER_10_187 ();
 FILLCELL_X8 FILLER_10_195 ();
 FILLCELL_X2 FILLER_10_207 ();
 FILLCELL_X4 FILLER_10_223 ();
 FILLCELL_X1 FILLER_10_227 ();
 FILLCELL_X16 FILLER_10_242 ();
 FILLCELL_X4 FILLER_10_258 ();
 FILLCELL_X8 FILLER_10_286 ();
 FILLCELL_X4 FILLER_10_301 ();
 FILLCELL_X2 FILLER_10_305 ();
 FILLCELL_X1 FILLER_10_307 ();
 FILLCELL_X8 FILLER_10_311 ();
 FILLCELL_X16 FILLER_10_326 ();
 FILLCELL_X1 FILLER_10_342 ();
 FILLCELL_X32 FILLER_10_350 ();
 FILLCELL_X1 FILLER_10_386 ();
 FILLCELL_X1 FILLER_10_390 ();
 FILLCELL_X32 FILLER_10_398 ();
 FILLCELL_X4 FILLER_10_430 ();
 FILLCELL_X1 FILLER_10_434 ();
 FILLCELL_X8 FILLER_10_438 ();
 FILLCELL_X4 FILLER_10_446 ();
 FILLCELL_X4 FILLER_10_460 ();
 FILLCELL_X1 FILLER_10_464 ();
 FILLCELL_X2 FILLER_10_475 ();
 FILLCELL_X32 FILLER_10_480 ();
 FILLCELL_X2 FILLER_10_521 ();
 FILLCELL_X4 FILLER_10_527 ();
 FILLCELL_X8 FILLER_10_539 ();
 FILLCELL_X2 FILLER_10_547 ();
 FILLCELL_X2 FILLER_10_568 ();
 FILLCELL_X1 FILLER_10_587 ();
 FILLCELL_X2 FILLER_10_607 ();
 FILLCELL_X4 FILLER_10_613 ();
 FILLCELL_X1 FILLER_10_617 ();
 FILLCELL_X8 FILLER_10_620 ();
 FILLCELL_X1 FILLER_10_628 ();
 FILLCELL_X16 FILLER_10_632 ();
 FILLCELL_X8 FILLER_10_648 ();
 FILLCELL_X4 FILLER_10_656 ();
 FILLCELL_X2 FILLER_10_660 ();
 FILLCELL_X4 FILLER_10_669 ();
 FILLCELL_X4 FILLER_10_690 ();
 FILLCELL_X4 FILLER_10_715 ();
 FILLCELL_X1 FILLER_10_719 ();
 FILLCELL_X8 FILLER_10_734 ();
 FILLCELL_X1 FILLER_10_742 ();
 FILLCELL_X2 FILLER_10_750 ();
 FILLCELL_X16 FILLER_10_769 ();
 FILLCELL_X1 FILLER_10_785 ();
 FILLCELL_X2 FILLER_10_792 ();
 FILLCELL_X8 FILLER_10_801 ();
 FILLCELL_X4 FILLER_10_809 ();
 FILLCELL_X1 FILLER_10_813 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X8 FILLER_11_97 ();
 FILLCELL_X4 FILLER_11_105 ();
 FILLCELL_X2 FILLER_11_109 ();
 FILLCELL_X1 FILLER_11_111 ();
 FILLCELL_X4 FILLER_11_184 ();
 FILLCELL_X4 FILLER_11_213 ();
 FILLCELL_X1 FILLER_11_217 ();
 FILLCELL_X2 FILLER_11_225 ();
 FILLCELL_X1 FILLER_11_227 ();
 FILLCELL_X2 FILLER_11_235 ();
 FILLCELL_X1 FILLER_11_246 ();
 FILLCELL_X2 FILLER_11_254 ();
 FILLCELL_X1 FILLER_11_256 ();
 FILLCELL_X16 FILLER_11_260 ();
 FILLCELL_X4 FILLER_11_276 ();
 FILLCELL_X2 FILLER_11_280 ();
 FILLCELL_X1 FILLER_11_285 ();
 FILLCELL_X2 FILLER_11_303 ();
 FILLCELL_X2 FILLER_11_309 ();
 FILLCELL_X2 FILLER_11_328 ();
 FILLCELL_X4 FILLER_11_333 ();
 FILLCELL_X16 FILLER_11_354 ();
 FILLCELL_X8 FILLER_11_370 ();
 FILLCELL_X2 FILLER_11_378 ();
 FILLCELL_X2 FILLER_11_383 ();
 FILLCELL_X2 FILLER_11_388 ();
 FILLCELL_X1 FILLER_11_390 ();
 FILLCELL_X16 FILLER_11_425 ();
 FILLCELL_X4 FILLER_11_441 ();
 FILLCELL_X1 FILLER_11_445 ();
 FILLCELL_X8 FILLER_11_449 ();
 FILLCELL_X1 FILLER_11_457 ();
 FILLCELL_X1 FILLER_11_467 ();
 FILLCELL_X2 FILLER_11_485 ();
 FILLCELL_X1 FILLER_11_487 ();
 FILLCELL_X16 FILLER_11_492 ();
 FILLCELL_X8 FILLER_11_508 ();
 FILLCELL_X4 FILLER_11_524 ();
 FILLCELL_X2 FILLER_11_528 ();
 FILLCELL_X1 FILLER_11_530 ();
 FILLCELL_X8 FILLER_11_548 ();
 FILLCELL_X1 FILLER_11_556 ();
 FILLCELL_X2 FILLER_11_561 ();
 FILLCELL_X2 FILLER_11_567 ();
 FILLCELL_X1 FILLER_11_569 ();
 FILLCELL_X1 FILLER_11_577 ();
 FILLCELL_X2 FILLER_11_582 ();
 FILLCELL_X1 FILLER_11_595 ();
 FILLCELL_X8 FILLER_11_607 ();
 FILLCELL_X2 FILLER_11_639 ();
 FILLCELL_X2 FILLER_11_662 ();
 FILLCELL_X4 FILLER_11_668 ();
 FILLCELL_X2 FILLER_11_672 ();
 FILLCELL_X2 FILLER_11_677 ();
 FILLCELL_X8 FILLER_11_683 ();
 FILLCELL_X4 FILLER_11_691 ();
 FILLCELL_X2 FILLER_11_695 ();
 FILLCELL_X8 FILLER_11_710 ();
 FILLCELL_X2 FILLER_11_725 ();
 FILLCELL_X4 FILLER_11_734 ();
 FILLCELL_X1 FILLER_11_738 ();
 FILLCELL_X16 FILLER_11_759 ();
 FILLCELL_X8 FILLER_11_775 ();
 FILLCELL_X2 FILLER_11_783 ();
 FILLCELL_X4 FILLER_11_789 ();
 FILLCELL_X4 FILLER_11_810 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X16 FILLER_12_65 ();
 FILLCELL_X8 FILLER_12_81 ();
 FILLCELL_X2 FILLER_12_89 ();
 FILLCELL_X8 FILLER_12_94 ();
 FILLCELL_X2 FILLER_12_102 ();
 FILLCELL_X4 FILLER_12_118 ();
 FILLCELL_X8 FILLER_12_136 ();
 FILLCELL_X4 FILLER_12_144 ();
 FILLCELL_X16 FILLER_12_155 ();
 FILLCELL_X4 FILLER_12_171 ();
 FILLCELL_X2 FILLER_12_175 ();
 FILLCELL_X8 FILLER_12_181 ();
 FILLCELL_X4 FILLER_12_189 ();
 FILLCELL_X1 FILLER_12_234 ();
 FILLCELL_X2 FILLER_12_261 ();
 FILLCELL_X1 FILLER_12_263 ();
 FILLCELL_X8 FILLER_12_288 ();
 FILLCELL_X4 FILLER_12_296 ();
 FILLCELL_X16 FILLER_12_303 ();
 FILLCELL_X8 FILLER_12_326 ();
 FILLCELL_X2 FILLER_12_334 ();
 FILLCELL_X1 FILLER_12_336 ();
 FILLCELL_X4 FILLER_12_341 ();
 FILLCELL_X4 FILLER_12_348 ();
 FILLCELL_X8 FILLER_12_367 ();
 FILLCELL_X2 FILLER_12_379 ();
 FILLCELL_X1 FILLER_12_381 ();
 FILLCELL_X2 FILLER_12_399 ();
 FILLCELL_X2 FILLER_12_408 ();
 FILLCELL_X2 FILLER_12_414 ();
 FILLCELL_X2 FILLER_12_419 ();
 FILLCELL_X1 FILLER_12_421 ();
 FILLCELL_X4 FILLER_12_439 ();
 FILLCELL_X1 FILLER_12_443 ();
 FILLCELL_X8 FILLER_12_448 ();
 FILLCELL_X8 FILLER_12_476 ();
 FILLCELL_X4 FILLER_12_504 ();
 FILLCELL_X2 FILLER_12_508 ();
 FILLCELL_X1 FILLER_12_510 ();
 FILLCELL_X4 FILLER_12_528 ();
 FILLCELL_X2 FILLER_12_532 ();
 FILLCELL_X1 FILLER_12_534 ();
 FILLCELL_X16 FILLER_12_542 ();
 FILLCELL_X4 FILLER_12_558 ();
 FILLCELL_X2 FILLER_12_583 ();
 FILLCELL_X4 FILLER_12_587 ();
 FILLCELL_X1 FILLER_12_591 ();
 FILLCELL_X4 FILLER_12_605 ();
 FILLCELL_X1 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X2 FILLER_12_632 ();
 FILLCELL_X1 FILLER_12_634 ();
 FILLCELL_X2 FILLER_12_637 ();
 FILLCELL_X4 FILLER_12_670 ();
 FILLCELL_X2 FILLER_12_674 ();
 FILLCELL_X1 FILLER_12_676 ();
 FILLCELL_X1 FILLER_12_701 ();
 FILLCELL_X1 FILLER_12_705 ();
 FILLCELL_X1 FILLER_12_711 ();
 FILLCELL_X1 FILLER_12_717 ();
 FILLCELL_X1 FILLER_12_721 ();
 FILLCELL_X8 FILLER_12_735 ();
 FILLCELL_X4 FILLER_12_743 ();
 FILLCELL_X1 FILLER_12_747 ();
 FILLCELL_X8 FILLER_12_751 ();
 FILLCELL_X4 FILLER_12_759 ();
 FILLCELL_X1 FILLER_12_763 ();
 FILLCELL_X4 FILLER_12_809 ();
 FILLCELL_X1 FILLER_12_813 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X16 FILLER_13_65 ();
 FILLCELL_X4 FILLER_13_81 ();
 FILLCELL_X1 FILLER_13_85 ();
 FILLCELL_X4 FILLER_13_90 ();
 FILLCELL_X2 FILLER_13_94 ();
 FILLCELL_X2 FILLER_13_113 ();
 FILLCELL_X1 FILLER_13_132 ();
 FILLCELL_X4 FILLER_13_154 ();
 FILLCELL_X1 FILLER_13_158 ();
 FILLCELL_X4 FILLER_13_164 ();
 FILLCELL_X2 FILLER_13_168 ();
 FILLCELL_X8 FILLER_13_187 ();
 FILLCELL_X4 FILLER_13_195 ();
 FILLCELL_X1 FILLER_13_199 ();
 FILLCELL_X4 FILLER_13_204 ();
 FILLCELL_X1 FILLER_13_208 ();
 FILLCELL_X16 FILLER_13_212 ();
 FILLCELL_X8 FILLER_13_235 ();
 FILLCELL_X4 FILLER_13_243 ();
 FILLCELL_X2 FILLER_13_247 ();
 FILLCELL_X1 FILLER_13_249 ();
 FILLCELL_X4 FILLER_13_254 ();
 FILLCELL_X1 FILLER_13_258 ();
 FILLCELL_X2 FILLER_13_262 ();
 FILLCELL_X1 FILLER_13_271 ();
 FILLCELL_X2 FILLER_13_279 ();
 FILLCELL_X8 FILLER_13_288 ();
 FILLCELL_X2 FILLER_13_296 ();
 FILLCELL_X2 FILLER_13_312 ();
 FILLCELL_X2 FILLER_13_331 ();
 FILLCELL_X4 FILLER_13_353 ();
 FILLCELL_X1 FILLER_13_357 ();
 FILLCELL_X4 FILLER_13_365 ();
 FILLCELL_X1 FILLER_13_417 ();
 FILLCELL_X2 FILLER_13_431 ();
 FILLCELL_X8 FILLER_13_450 ();
 FILLCELL_X2 FILLER_13_458 ();
 FILLCELL_X16 FILLER_13_463 ();
 FILLCELL_X4 FILLER_13_479 ();
 FILLCELL_X2 FILLER_13_493 ();
 FILLCELL_X1 FILLER_13_495 ();
 FILLCELL_X16 FILLER_13_510 ();
 FILLCELL_X8 FILLER_13_526 ();
 FILLCELL_X2 FILLER_13_534 ();
 FILLCELL_X1 FILLER_13_536 ();
 FILLCELL_X16 FILLER_13_548 ();
 FILLCELL_X1 FILLER_13_564 ();
 FILLCELL_X2 FILLER_13_569 ();
 FILLCELL_X4 FILLER_13_579 ();
 FILLCELL_X8 FILLER_13_585 ();
 FILLCELL_X1 FILLER_13_593 ();
 FILLCELL_X2 FILLER_13_610 ();
 FILLCELL_X1 FILLER_13_612 ();
 FILLCELL_X16 FILLER_13_621 ();
 FILLCELL_X4 FILLER_13_637 ();
 FILLCELL_X2 FILLER_13_641 ();
 FILLCELL_X1 FILLER_13_643 ();
 FILLCELL_X4 FILLER_13_651 ();
 FILLCELL_X8 FILLER_13_685 ();
 FILLCELL_X4 FILLER_13_700 ();
 FILLCELL_X4 FILLER_13_713 ();
 FILLCELL_X8 FILLER_13_734 ();
 FILLCELL_X1 FILLER_13_742 ();
 FILLCELL_X4 FILLER_13_745 ();
 FILLCELL_X2 FILLER_13_749 ();
 FILLCELL_X8 FILLER_13_755 ();
 FILLCELL_X2 FILLER_13_763 ();
 FILLCELL_X1 FILLER_13_765 ();
 FILLCELL_X8 FILLER_13_780 ();
 FILLCELL_X16 FILLER_13_798 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X4 FILLER_14_65 ();
 FILLCELL_X2 FILLER_14_69 ();
 FILLCELL_X8 FILLER_14_94 ();
 FILLCELL_X4 FILLER_14_102 ();
 FILLCELL_X16 FILLER_14_109 ();
 FILLCELL_X16 FILLER_14_128 ();
 FILLCELL_X1 FILLER_14_144 ();
 FILLCELL_X2 FILLER_14_184 ();
 FILLCELL_X4 FILLER_14_193 ();
 FILLCELL_X2 FILLER_14_206 ();
 FILLCELL_X8 FILLER_14_229 ();
 FILLCELL_X8 FILLER_14_261 ();
 FILLCELL_X2 FILLER_14_269 ();
 FILLCELL_X8 FILLER_14_278 ();
 FILLCELL_X1 FILLER_14_286 ();
 FILLCELL_X8 FILLER_14_307 ();
 FILLCELL_X1 FILLER_14_315 ();
 FILLCELL_X1 FILLER_14_323 ();
 FILLCELL_X8 FILLER_14_327 ();
 FILLCELL_X4 FILLER_14_335 ();
 FILLCELL_X2 FILLER_14_339 ();
 FILLCELL_X1 FILLER_14_341 ();
 FILLCELL_X2 FILLER_14_345 ();
 FILLCELL_X1 FILLER_14_347 ();
 FILLCELL_X8 FILLER_14_362 ();
 FILLCELL_X4 FILLER_14_370 ();
 FILLCELL_X2 FILLER_14_374 ();
 FILLCELL_X4 FILLER_14_379 ();
 FILLCELL_X2 FILLER_14_383 ();
 FILLCELL_X1 FILLER_14_385 ();
 FILLCELL_X16 FILLER_14_407 ();
 FILLCELL_X8 FILLER_14_423 ();
 FILLCELL_X2 FILLER_14_431 ();
 FILLCELL_X4 FILLER_14_440 ();
 FILLCELL_X1 FILLER_14_444 ();
 FILLCELL_X2 FILLER_14_452 ();
 FILLCELL_X1 FILLER_14_454 ();
 FILLCELL_X1 FILLER_14_458 ();
 FILLCELL_X1 FILLER_14_463 ();
 FILLCELL_X1 FILLER_14_467 ();
 FILLCELL_X1 FILLER_14_485 ();
 FILLCELL_X1 FILLER_14_493 ();
 FILLCELL_X2 FILLER_14_506 ();
 FILLCELL_X2 FILLER_14_513 ();
 FILLCELL_X1 FILLER_14_515 ();
 FILLCELL_X8 FILLER_14_532 ();
 FILLCELL_X1 FILLER_14_540 ();
 FILLCELL_X8 FILLER_14_571 ();
 FILLCELL_X4 FILLER_14_579 ();
 FILLCELL_X2 FILLER_14_583 ();
 FILLCELL_X1 FILLER_14_585 ();
 FILLCELL_X4 FILLER_14_600 ();
 FILLCELL_X4 FILLER_14_623 ();
 FILLCELL_X1 FILLER_14_627 ();
 FILLCELL_X8 FILLER_14_632 ();
 FILLCELL_X4 FILLER_14_640 ();
 FILLCELL_X2 FILLER_14_661 ();
 FILLCELL_X8 FILLER_14_668 ();
 FILLCELL_X4 FILLER_14_676 ();
 FILLCELL_X2 FILLER_14_680 ();
 FILLCELL_X1 FILLER_14_682 ();
 FILLCELL_X8 FILLER_14_690 ();
 FILLCELL_X1 FILLER_14_698 ();
 FILLCELL_X4 FILLER_14_706 ();
 FILLCELL_X1 FILLER_14_710 ();
 FILLCELL_X4 FILLER_14_714 ();
 FILLCELL_X1 FILLER_14_718 ();
 FILLCELL_X4 FILLER_14_722 ();
 FILLCELL_X1 FILLER_14_726 ();
 FILLCELL_X8 FILLER_14_733 ();
 FILLCELL_X2 FILLER_14_741 ();
 FILLCELL_X4 FILLER_14_786 ();
 FILLCELL_X2 FILLER_14_790 ();
 FILLCELL_X4 FILLER_14_809 ();
 FILLCELL_X1 FILLER_14_813 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X16 FILLER_15_33 ();
 FILLCELL_X4 FILLER_15_49 ();
 FILLCELL_X4 FILLER_15_74 ();
 FILLCELL_X2 FILLER_15_78 ();
 FILLCELL_X4 FILLER_15_101 ();
 FILLCELL_X2 FILLER_15_105 ();
 FILLCELL_X1 FILLER_15_107 ();
 FILLCELL_X16 FILLER_15_115 ();
 FILLCELL_X8 FILLER_15_131 ();
 FILLCELL_X8 FILLER_15_155 ();
 FILLCELL_X1 FILLER_15_163 ();
 FILLCELL_X4 FILLER_15_172 ();
 FILLCELL_X1 FILLER_15_176 ();
 FILLCELL_X4 FILLER_15_180 ();
 FILLCELL_X1 FILLER_15_184 ();
 FILLCELL_X2 FILLER_15_206 ();
 FILLCELL_X2 FILLER_15_211 ();
 FILLCELL_X8 FILLER_15_216 ();
 FILLCELL_X2 FILLER_15_224 ();
 FILLCELL_X8 FILLER_15_240 ();
 FILLCELL_X2 FILLER_15_248 ();
 FILLCELL_X16 FILLER_15_253 ();
 FILLCELL_X2 FILLER_15_269 ();
 FILLCELL_X1 FILLER_15_271 ();
 FILLCELL_X4 FILLER_15_286 ();
 FILLCELL_X2 FILLER_15_290 ();
 FILLCELL_X1 FILLER_15_292 ();
 FILLCELL_X1 FILLER_15_300 ();
 FILLCELL_X4 FILLER_15_308 ();
 FILLCELL_X1 FILLER_15_319 ();
 FILLCELL_X1 FILLER_15_327 ();
 FILLCELL_X8 FILLER_15_342 ();
 FILLCELL_X4 FILLER_15_350 ();
 FILLCELL_X16 FILLER_15_361 ();
 FILLCELL_X8 FILLER_15_377 ();
 FILLCELL_X4 FILLER_15_385 ();
 FILLCELL_X2 FILLER_15_389 ();
 FILLCELL_X8 FILLER_15_419 ();
 FILLCELL_X2 FILLER_15_427 ();
 FILLCELL_X2 FILLER_15_463 ();
 FILLCELL_X2 FILLER_15_469 ();
 FILLCELL_X16 FILLER_15_474 ();
 FILLCELL_X4 FILLER_15_490 ();
 FILLCELL_X4 FILLER_15_506 ();
 FILLCELL_X1 FILLER_15_510 ();
 FILLCELL_X2 FILLER_15_540 ();
 FILLCELL_X1 FILLER_15_559 ();
 FILLCELL_X2 FILLER_15_565 ();
 FILLCELL_X2 FILLER_15_586 ();
 FILLCELL_X4 FILLER_15_594 ();
 FILLCELL_X1 FILLER_15_598 ();
 FILLCELL_X4 FILLER_15_604 ();
 FILLCELL_X1 FILLER_15_608 ();
 FILLCELL_X16 FILLER_15_611 ();
 FILLCELL_X8 FILLER_15_631 ();
 FILLCELL_X1 FILLER_15_639 ();
 FILLCELL_X2 FILLER_15_647 ();
 FILLCELL_X1 FILLER_15_649 ();
 FILLCELL_X1 FILLER_15_665 ();
 FILLCELL_X4 FILLER_15_673 ();
 FILLCELL_X2 FILLER_15_677 ();
 FILLCELL_X4 FILLER_15_696 ();
 FILLCELL_X1 FILLER_15_700 ();
 FILLCELL_X4 FILLER_15_704 ();
 FILLCELL_X1 FILLER_15_711 ();
 FILLCELL_X1 FILLER_15_721 ();
 FILLCELL_X4 FILLER_15_728 ();
 FILLCELL_X2 FILLER_15_732 ();
 FILLCELL_X1 FILLER_15_734 ();
 FILLCELL_X2 FILLER_15_746 ();
 FILLCELL_X4 FILLER_15_755 ();
 FILLCELL_X4 FILLER_15_766 ();
 FILLCELL_X2 FILLER_15_770 ();
 FILLCELL_X1 FILLER_15_772 ();
 FILLCELL_X8 FILLER_15_783 ();
 FILLCELL_X1 FILLER_15_791 ();
 FILLCELL_X1 FILLER_15_795 ();
 FILLCELL_X1 FILLER_15_813 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X16 FILLER_16_33 ();
 FILLCELL_X8 FILLER_16_49 ();
 FILLCELL_X4 FILLER_16_57 ();
 FILLCELL_X2 FILLER_16_85 ();
 FILLCELL_X1 FILLER_16_87 ();
 FILLCELL_X4 FILLER_16_95 ();
 FILLCELL_X2 FILLER_16_99 ();
 FILLCELL_X2 FILLER_16_118 ();
 FILLCELL_X1 FILLER_16_120 ();
 FILLCELL_X16 FILLER_16_131 ();
 FILLCELL_X4 FILLER_16_156 ();
 FILLCELL_X8 FILLER_16_168 ();
 FILLCELL_X4 FILLER_16_180 ();
 FILLCELL_X2 FILLER_16_184 ();
 FILLCELL_X1 FILLER_16_186 ();
 FILLCELL_X2 FILLER_16_190 ();
 FILLCELL_X1 FILLER_16_192 ();
 FILLCELL_X4 FILLER_16_200 ();
 FILLCELL_X2 FILLER_16_204 ();
 FILLCELL_X1 FILLER_16_206 ();
 FILLCELL_X4 FILLER_16_214 ();
 FILLCELL_X16 FILLER_16_232 ();
 FILLCELL_X1 FILLER_16_248 ();
 FILLCELL_X2 FILLER_16_253 ();
 FILLCELL_X1 FILLER_16_255 ();
 FILLCELL_X4 FILLER_16_259 ();
 FILLCELL_X2 FILLER_16_263 ();
 FILLCELL_X1 FILLER_16_265 ();
 FILLCELL_X4 FILLER_16_273 ();
 FILLCELL_X1 FILLER_16_277 ();
 FILLCELL_X4 FILLER_16_283 ();
 FILLCELL_X1 FILLER_16_287 ();
 FILLCELL_X2 FILLER_16_295 ();
 FILLCELL_X8 FILLER_16_311 ();
 FILLCELL_X4 FILLER_16_319 ();
 FILLCELL_X2 FILLER_16_323 ();
 FILLCELL_X1 FILLER_16_325 ();
 FILLCELL_X1 FILLER_16_329 ();
 FILLCELL_X8 FILLER_16_337 ();
 FILLCELL_X4 FILLER_16_345 ();
 FILLCELL_X1 FILLER_16_349 ();
 FILLCELL_X4 FILLER_16_357 ();
 FILLCELL_X2 FILLER_16_361 ();
 FILLCELL_X1 FILLER_16_363 ();
 FILLCELL_X8 FILLER_16_381 ();
 FILLCELL_X2 FILLER_16_389 ();
 FILLCELL_X32 FILLER_16_398 ();
 FILLCELL_X2 FILLER_16_430 ();
 FILLCELL_X1 FILLER_16_432 ();
 FILLCELL_X8 FILLER_16_436 ();
 FILLCELL_X4 FILLER_16_444 ();
 FILLCELL_X1 FILLER_16_448 ();
 FILLCELL_X4 FILLER_16_452 ();
 FILLCELL_X2 FILLER_16_456 ();
 FILLCELL_X16 FILLER_16_478 ();
 FILLCELL_X1 FILLER_16_494 ();
 FILLCELL_X4 FILLER_16_509 ();
 FILLCELL_X2 FILLER_16_513 ();
 FILLCELL_X1 FILLER_16_515 ();
 FILLCELL_X8 FILLER_16_530 ();
 FILLCELL_X2 FILLER_16_538 ();
 FILLCELL_X1 FILLER_16_557 ();
 FILLCELL_X1 FILLER_16_571 ();
 FILLCELL_X4 FILLER_16_610 ();
 FILLCELL_X8 FILLER_16_635 ();
 FILLCELL_X2 FILLER_16_643 ();
 FILLCELL_X1 FILLER_16_645 ();
 FILLCELL_X4 FILLER_16_662 ();
 FILLCELL_X2 FILLER_16_683 ();
 FILLCELL_X4 FILLER_16_688 ();
 FILLCELL_X4 FILLER_16_699 ();
 FILLCELL_X1 FILLER_16_703 ();
 FILLCELL_X1 FILLER_16_713 ();
 FILLCELL_X8 FILLER_16_740 ();
 FILLCELL_X16 FILLER_16_755 ();
 FILLCELL_X2 FILLER_16_771 ();
 FILLCELL_X1 FILLER_16_773 ();
 FILLCELL_X1 FILLER_16_780 ();
 FILLCELL_X4 FILLER_16_784 ();
 FILLCELL_X1 FILLER_16_788 ();
 FILLCELL_X8 FILLER_16_803 ();
 FILLCELL_X2 FILLER_16_811 ();
 FILLCELL_X1 FILLER_16_813 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X8 FILLER_17_69 ();
 FILLCELL_X2 FILLER_17_91 ();
 FILLCELL_X1 FILLER_17_93 ();
 FILLCELL_X2 FILLER_17_111 ();
 FILLCELL_X1 FILLER_17_154 ();
 FILLCELL_X4 FILLER_17_196 ();
 FILLCELL_X2 FILLER_17_200 ();
 FILLCELL_X1 FILLER_17_202 ();
 FILLCELL_X1 FILLER_17_220 ();
 FILLCELL_X2 FILLER_17_228 ();
 FILLCELL_X2 FILLER_17_237 ();
 FILLCELL_X2 FILLER_17_256 ();
 FILLCELL_X1 FILLER_17_258 ();
 FILLCELL_X4 FILLER_17_276 ();
 FILLCELL_X1 FILLER_17_280 ();
 FILLCELL_X2 FILLER_17_286 ();
 FILLCELL_X4 FILLER_17_295 ();
 FILLCELL_X1 FILLER_17_299 ();
 FILLCELL_X8 FILLER_17_338 ();
 FILLCELL_X2 FILLER_17_360 ();
 FILLCELL_X1 FILLER_17_362 ();
 FILLCELL_X1 FILLER_17_373 ();
 FILLCELL_X1 FILLER_17_377 ();
 FILLCELL_X2 FILLER_17_392 ();
 FILLCELL_X1 FILLER_17_394 ();
 FILLCELL_X1 FILLER_17_409 ();
 FILLCELL_X4 FILLER_17_427 ();
 FILLCELL_X4 FILLER_17_448 ();
 FILLCELL_X8 FILLER_17_459 ();
 FILLCELL_X1 FILLER_17_467 ();
 FILLCELL_X16 FILLER_17_475 ();
 FILLCELL_X32 FILLER_17_495 ();
 FILLCELL_X8 FILLER_17_529 ();
 FILLCELL_X4 FILLER_17_537 ();
 FILLCELL_X2 FILLER_17_541 ();
 FILLCELL_X8 FILLER_17_564 ();
 FILLCELL_X1 FILLER_17_572 ();
 FILLCELL_X1 FILLER_17_577 ();
 FILLCELL_X4 FILLER_17_587 ();
 FILLCELL_X2 FILLER_17_591 ();
 FILLCELL_X4 FILLER_17_598 ();
 FILLCELL_X2 FILLER_17_602 ();
 FILLCELL_X4 FILLER_17_617 ();
 FILLCELL_X2 FILLER_17_621 ();
 FILLCELL_X2 FILLER_17_639 ();
 FILLCELL_X8 FILLER_17_658 ();
 FILLCELL_X16 FILLER_17_674 ();
 FILLCELL_X2 FILLER_17_690 ();
 FILLCELL_X2 FILLER_17_703 ();
 FILLCELL_X1 FILLER_17_705 ();
 FILLCELL_X4 FILLER_17_718 ();
 FILLCELL_X8 FILLER_17_726 ();
 FILLCELL_X2 FILLER_17_741 ();
 FILLCELL_X1 FILLER_17_743 ();
 FILLCELL_X8 FILLER_17_751 ();
 FILLCELL_X1 FILLER_17_759 ();
 FILLCELL_X8 FILLER_17_784 ();
 FILLCELL_X8 FILLER_17_802 ();
 FILLCELL_X4 FILLER_17_810 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X8 FILLER_18_33 ();
 FILLCELL_X4 FILLER_18_41 ();
 FILLCELL_X2 FILLER_18_45 ();
 FILLCELL_X1 FILLER_18_47 ();
 FILLCELL_X8 FILLER_18_69 ();
 FILLCELL_X4 FILLER_18_77 ();
 FILLCELL_X2 FILLER_18_81 ();
 FILLCELL_X8 FILLER_18_86 ();
 FILLCELL_X4 FILLER_18_94 ();
 FILLCELL_X2 FILLER_18_98 ();
 FILLCELL_X1 FILLER_18_100 ();
 FILLCELL_X1 FILLER_18_109 ();
 FILLCELL_X8 FILLER_18_124 ();
 FILLCELL_X2 FILLER_18_132 ();
 FILLCELL_X1 FILLER_18_134 ();
 FILLCELL_X4 FILLER_18_142 ();
 FILLCELL_X1 FILLER_18_146 ();
 FILLCELL_X32 FILLER_18_154 ();
 FILLCELL_X4 FILLER_18_186 ();
 FILLCELL_X2 FILLER_18_190 ();
 FILLCELL_X1 FILLER_18_192 ();
 FILLCELL_X16 FILLER_18_210 ();
 FILLCELL_X4 FILLER_18_226 ();
 FILLCELL_X2 FILLER_18_230 ();
 FILLCELL_X1 FILLER_18_232 ();
 FILLCELL_X8 FILLER_18_240 ();
 FILLCELL_X1 FILLER_18_248 ();
 FILLCELL_X16 FILLER_18_252 ();
 FILLCELL_X1 FILLER_18_268 ();
 FILLCELL_X8 FILLER_18_272 ();
 FILLCELL_X1 FILLER_18_280 ();
 FILLCELL_X8 FILLER_18_288 ();
 FILLCELL_X4 FILLER_18_296 ();
 FILLCELL_X8 FILLER_18_308 ();
 FILLCELL_X2 FILLER_18_316 ();
 FILLCELL_X1 FILLER_18_318 ();
 FILLCELL_X8 FILLER_18_333 ();
 FILLCELL_X2 FILLER_18_341 ();
 FILLCELL_X4 FILLER_18_371 ();
 FILLCELL_X2 FILLER_18_375 ();
 FILLCELL_X2 FILLER_18_398 ();
 FILLCELL_X2 FILLER_18_407 ();
 FILLCELL_X1 FILLER_18_416 ();
 FILLCELL_X2 FILLER_18_424 ();
 FILLCELL_X1 FILLER_18_429 ();
 FILLCELL_X2 FILLER_18_440 ();
 FILLCELL_X8 FILLER_18_474 ();
 FILLCELL_X4 FILLER_18_482 ();
 FILLCELL_X4 FILLER_18_508 ();
 FILLCELL_X8 FILLER_18_530 ();
 FILLCELL_X4 FILLER_18_538 ();
 FILLCELL_X1 FILLER_18_553 ();
 FILLCELL_X4 FILLER_18_558 ();
 FILLCELL_X2 FILLER_18_562 ();
 FILLCELL_X1 FILLER_18_564 ();
 FILLCELL_X8 FILLER_18_576 ();
 FILLCELL_X4 FILLER_18_584 ();
 FILLCELL_X2 FILLER_18_588 ();
 FILLCELL_X1 FILLER_18_590 ();
 FILLCELL_X4 FILLER_18_614 ();
 FILLCELL_X2 FILLER_18_618 ();
 FILLCELL_X8 FILLER_18_622 ();
 FILLCELL_X1 FILLER_18_630 ();
 FILLCELL_X4 FILLER_18_636 ();
 FILLCELL_X8 FILLER_18_652 ();
 FILLCELL_X4 FILLER_18_660 ();
 FILLCELL_X2 FILLER_18_664 ();
 FILLCELL_X1 FILLER_18_666 ();
 FILLCELL_X16 FILLER_18_675 ();
 FILLCELL_X1 FILLER_18_691 ();
 FILLCELL_X1 FILLER_18_702 ();
 FILLCELL_X8 FILLER_18_707 ();
 FILLCELL_X4 FILLER_18_715 ();
 FILLCELL_X1 FILLER_18_719 ();
 FILLCELL_X4 FILLER_18_725 ();
 FILLCELL_X2 FILLER_18_729 ();
 FILLCELL_X16 FILLER_18_747 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X16 FILLER_19_33 ();
 FILLCELL_X8 FILLER_19_49 ();
 FILLCELL_X1 FILLER_19_61 ();
 FILLCELL_X1 FILLER_19_66 ();
 FILLCELL_X8 FILLER_19_91 ();
 FILLCELL_X2 FILLER_19_99 ();
 FILLCELL_X1 FILLER_19_101 ();
 FILLCELL_X2 FILLER_19_117 ();
 FILLCELL_X1 FILLER_19_119 ();
 FILLCELL_X4 FILLER_19_122 ();
 FILLCELL_X2 FILLER_19_126 ();
 FILLCELL_X8 FILLER_19_136 ();
 FILLCELL_X1 FILLER_19_144 ();
 FILLCELL_X32 FILLER_19_152 ();
 FILLCELL_X2 FILLER_19_184 ();
 FILLCELL_X1 FILLER_19_186 ();
 FILLCELL_X1 FILLER_19_203 ();
 FILLCELL_X2 FILLER_19_211 ();
 FILLCELL_X8 FILLER_19_216 ();
 FILLCELL_X1 FILLER_19_231 ();
 FILLCELL_X2 FILLER_19_239 ();
 FILLCELL_X16 FILLER_19_244 ();
 FILLCELL_X8 FILLER_19_260 ();
 FILLCELL_X1 FILLER_19_268 ();
 FILLCELL_X1 FILLER_19_276 ();
 FILLCELL_X2 FILLER_19_280 ();
 FILLCELL_X2 FILLER_19_299 ();
 FILLCELL_X2 FILLER_19_310 ();
 FILLCELL_X1 FILLER_19_312 ();
 FILLCELL_X2 FILLER_19_322 ();
 FILLCELL_X1 FILLER_19_324 ();
 FILLCELL_X2 FILLER_19_332 ();
 FILLCELL_X8 FILLER_19_355 ();
 FILLCELL_X1 FILLER_19_385 ();
 FILLCELL_X8 FILLER_19_394 ();
 FILLCELL_X32 FILLER_19_409 ();
 FILLCELL_X4 FILLER_19_441 ();
 FILLCELL_X4 FILLER_19_448 ();
 FILLCELL_X2 FILLER_19_452 ();
 FILLCELL_X4 FILLER_19_457 ();
 FILLCELL_X2 FILLER_19_488 ();
 FILLCELL_X1 FILLER_19_493 ();
 FILLCELL_X2 FILLER_19_497 ();
 FILLCELL_X1 FILLER_19_499 ();
 FILLCELL_X2 FILLER_19_507 ();
 FILLCELL_X1 FILLER_19_512 ();
 FILLCELL_X2 FILLER_19_528 ();
 FILLCELL_X8 FILLER_19_545 ();
 FILLCELL_X4 FILLER_19_553 ();
 FILLCELL_X1 FILLER_19_557 ();
 FILLCELL_X16 FILLER_19_570 ();
 FILLCELL_X8 FILLER_19_586 ();
 FILLCELL_X8 FILLER_19_600 ();
 FILLCELL_X1 FILLER_19_608 ();
 FILLCELL_X8 FILLER_19_626 ();
 FILLCELL_X2 FILLER_19_638 ();
 FILLCELL_X8 FILLER_19_660 ();
 FILLCELL_X2 FILLER_19_676 ();
 FILLCELL_X1 FILLER_19_678 ();
 FILLCELL_X2 FILLER_19_700 ();
 FILLCELL_X1 FILLER_19_702 ();
 FILLCELL_X4 FILLER_19_710 ();
 FILLCELL_X2 FILLER_19_714 ();
 FILLCELL_X16 FILLER_19_733 ();
 FILLCELL_X1 FILLER_19_749 ();
 FILLCELL_X16 FILLER_19_757 ();
 FILLCELL_X4 FILLER_19_773 ();
 FILLCELL_X2 FILLER_19_777 ();
 FILLCELL_X1 FILLER_19_779 ();
 FILLCELL_X2 FILLER_19_783 ();
 FILLCELL_X1 FILLER_19_785 ();
 FILLCELL_X4 FILLER_19_808 ();
 FILLCELL_X2 FILLER_19_812 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X8 FILLER_20_33 ();
 FILLCELL_X4 FILLER_20_41 ();
 FILLCELL_X2 FILLER_20_45 ();
 FILLCELL_X1 FILLER_20_73 ();
 FILLCELL_X2 FILLER_20_81 ();
 FILLCELL_X2 FILLER_20_90 ();
 FILLCELL_X1 FILLER_20_116 ();
 FILLCELL_X4 FILLER_20_139 ();
 FILLCELL_X2 FILLER_20_143 ();
 FILLCELL_X8 FILLER_20_168 ();
 FILLCELL_X2 FILLER_20_201 ();
 FILLCELL_X2 FILLER_20_220 ();
 FILLCELL_X1 FILLER_20_231 ();
 FILLCELL_X2 FILLER_20_244 ();
 FILLCELL_X2 FILLER_20_253 ();
 FILLCELL_X1 FILLER_20_255 ();
 FILLCELL_X2 FILLER_20_259 ();
 FILLCELL_X16 FILLER_20_278 ();
 FILLCELL_X4 FILLER_20_294 ();
 FILLCELL_X2 FILLER_20_298 ();
 FILLCELL_X1 FILLER_20_317 ();
 FILLCELL_X4 FILLER_20_338 ();
 FILLCELL_X2 FILLER_20_342 ();
 FILLCELL_X8 FILLER_20_351 ();
 FILLCELL_X2 FILLER_20_359 ();
 FILLCELL_X1 FILLER_20_361 ();
 FILLCELL_X2 FILLER_20_373 ();
 FILLCELL_X2 FILLER_20_378 ();
 FILLCELL_X4 FILLER_20_384 ();
 FILLCELL_X16 FILLER_20_416 ();
 FILLCELL_X2 FILLER_20_432 ();
 FILLCELL_X1 FILLER_20_438 ();
 FILLCELL_X8 FILLER_20_442 ();
 FILLCELL_X2 FILLER_20_450 ();
 FILLCELL_X32 FILLER_20_456 ();
 FILLCELL_X4 FILLER_20_488 ();
 FILLCELL_X2 FILLER_20_492 ();
 FILLCELL_X4 FILLER_20_496 ();
 FILLCELL_X1 FILLER_20_500 ();
 FILLCELL_X16 FILLER_20_511 ();
 FILLCELL_X4 FILLER_20_533 ();
 FILLCELL_X1 FILLER_20_537 ();
 FILLCELL_X2 FILLER_20_547 ();
 FILLCELL_X2 FILLER_20_554 ();
 FILLCELL_X1 FILLER_20_556 ();
 FILLCELL_X4 FILLER_20_559 ();
 FILLCELL_X2 FILLER_20_563 ();
 FILLCELL_X2 FILLER_20_586 ();
 FILLCELL_X1 FILLER_20_588 ();
 FILLCELL_X16 FILLER_20_600 ();
 FILLCELL_X8 FILLER_20_620 ();
 FILLCELL_X8 FILLER_20_632 ();
 FILLCELL_X4 FILLER_20_640 ();
 FILLCELL_X1 FILLER_20_644 ();
 FILLCELL_X4 FILLER_20_648 ();
 FILLCELL_X2 FILLER_20_652 ();
 FILLCELL_X1 FILLER_20_654 ();
 FILLCELL_X8 FILLER_20_659 ();
 FILLCELL_X4 FILLER_20_684 ();
 FILLCELL_X4 FILLER_20_710 ();
 FILLCELL_X2 FILLER_20_714 ();
 FILLCELL_X4 FILLER_20_730 ();
 FILLCELL_X1 FILLER_20_734 ();
 FILLCELL_X4 FILLER_20_737 ();
 FILLCELL_X2 FILLER_20_741 ();
 FILLCELL_X1 FILLER_20_743 ();
 FILLCELL_X8 FILLER_20_761 ();
 FILLCELL_X2 FILLER_20_776 ();
 FILLCELL_X1 FILLER_20_778 ();
 FILLCELL_X4 FILLER_20_783 ();
 FILLCELL_X2 FILLER_20_787 ();
 FILLCELL_X8 FILLER_20_802 ();
 FILLCELL_X4 FILLER_20_810 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X16 FILLER_21_33 ();
 FILLCELL_X8 FILLER_21_49 ();
 FILLCELL_X8 FILLER_21_60 ();
 FILLCELL_X4 FILLER_21_68 ();
 FILLCELL_X2 FILLER_21_72 ();
 FILLCELL_X8 FILLER_21_88 ();
 FILLCELL_X2 FILLER_21_96 ();
 FILLCELL_X1 FILLER_21_98 ();
 FILLCELL_X8 FILLER_21_120 ();
 FILLCELL_X2 FILLER_21_128 ();
 FILLCELL_X8 FILLER_21_165 ();
 FILLCELL_X2 FILLER_21_173 ();
 FILLCELL_X8 FILLER_21_179 ();
 FILLCELL_X4 FILLER_21_211 ();
 FILLCELL_X1 FILLER_21_215 ();
 FILLCELL_X4 FILLER_21_219 ();
 FILLCELL_X4 FILLER_21_237 ();
 FILLCELL_X2 FILLER_21_241 ();
 FILLCELL_X4 FILLER_21_260 ();
 FILLCELL_X8 FILLER_21_285 ();
 FILLCELL_X1 FILLER_21_293 ();
 FILLCELL_X8 FILLER_21_302 ();
 FILLCELL_X2 FILLER_21_310 ();
 FILLCELL_X1 FILLER_21_312 ();
 FILLCELL_X16 FILLER_21_316 ();
 FILLCELL_X4 FILLER_21_332 ();
 FILLCELL_X1 FILLER_21_336 ();
 FILLCELL_X2 FILLER_21_354 ();
 FILLCELL_X4 FILLER_21_373 ();
 FILLCELL_X1 FILLER_21_377 ();
 FILLCELL_X16 FILLER_21_395 ();
 FILLCELL_X4 FILLER_21_411 ();
 FILLCELL_X1 FILLER_21_415 ();
 FILLCELL_X4 FILLER_21_426 ();
 FILLCELL_X2 FILLER_21_447 ();
 FILLCELL_X1 FILLER_21_449 ();
 FILLCELL_X2 FILLER_21_470 ();
 FILLCELL_X2 FILLER_21_476 ();
 FILLCELL_X4 FILLER_21_481 ();
 FILLCELL_X1 FILLER_21_485 ();
 FILLCELL_X1 FILLER_21_505 ();
 FILLCELL_X8 FILLER_21_513 ();
 FILLCELL_X2 FILLER_21_521 ();
 FILLCELL_X1 FILLER_21_523 ();
 FILLCELL_X1 FILLER_21_537 ();
 FILLCELL_X2 FILLER_21_572 ();
 FILLCELL_X4 FILLER_21_578 ();
 FILLCELL_X2 FILLER_21_582 ();
 FILLCELL_X1 FILLER_21_597 ();
 FILLCELL_X4 FILLER_21_663 ();
 FILLCELL_X1 FILLER_21_680 ();
 FILLCELL_X8 FILLER_21_686 ();
 FILLCELL_X4 FILLER_21_700 ();
 FILLCELL_X2 FILLER_21_708 ();
 FILLCELL_X16 FILLER_21_730 ();
 FILLCELL_X4 FILLER_21_746 ();
 FILLCELL_X2 FILLER_21_750 ();
 FILLCELL_X4 FILLER_21_755 ();
 FILLCELL_X2 FILLER_21_759 ();
 FILLCELL_X1 FILLER_21_765 ();
 FILLCELL_X2 FILLER_21_793 ();
 FILLCELL_X1 FILLER_21_795 ();
 FILLCELL_X1 FILLER_21_813 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X16 FILLER_22_33 ();
 FILLCELL_X8 FILLER_22_49 ();
 FILLCELL_X1 FILLER_22_57 ();
 FILLCELL_X1 FILLER_22_62 ();
 FILLCELL_X4 FILLER_22_67 ();
 FILLCELL_X1 FILLER_22_71 ();
 FILLCELL_X4 FILLER_22_83 ();
 FILLCELL_X16 FILLER_22_90 ();
 FILLCELL_X4 FILLER_22_106 ();
 FILLCELL_X1 FILLER_22_131 ();
 FILLCELL_X4 FILLER_22_135 ();
 FILLCELL_X1 FILLER_22_139 ();
 FILLCELL_X1 FILLER_22_152 ();
 FILLCELL_X8 FILLER_22_160 ();
 FILLCELL_X2 FILLER_22_168 ();
 FILLCELL_X1 FILLER_22_170 ();
 FILLCELL_X8 FILLER_22_188 ();
 FILLCELL_X8 FILLER_22_203 ();
 FILLCELL_X2 FILLER_22_211 ();
 FILLCELL_X1 FILLER_22_213 ();
 FILLCELL_X8 FILLER_22_238 ();
 FILLCELL_X2 FILLER_22_246 ();
 FILLCELL_X1 FILLER_22_248 ();
 FILLCELL_X16 FILLER_22_253 ();
 FILLCELL_X2 FILLER_22_290 ();
 FILLCELL_X4 FILLER_22_309 ();
 FILLCELL_X16 FILLER_22_320 ();
 FILLCELL_X8 FILLER_22_336 ();
 FILLCELL_X4 FILLER_22_344 ();
 FILLCELL_X2 FILLER_22_348 ();
 FILLCELL_X2 FILLER_22_353 ();
 FILLCELL_X1 FILLER_22_355 ();
 FILLCELL_X16 FILLER_22_366 ();
 FILLCELL_X4 FILLER_22_382 ();
 FILLCELL_X1 FILLER_22_386 ();
 FILLCELL_X16 FILLER_22_391 ();
 FILLCELL_X8 FILLER_22_407 ();
 FILLCELL_X2 FILLER_22_432 ();
 FILLCELL_X1 FILLER_22_434 ();
 FILLCELL_X4 FILLER_22_438 ();
 FILLCELL_X2 FILLER_22_442 ();
 FILLCELL_X1 FILLER_22_444 ();
 FILLCELL_X2 FILLER_22_448 ();
 FILLCELL_X8 FILLER_22_460 ();
 FILLCELL_X2 FILLER_22_492 ();
 FILLCELL_X2 FILLER_22_511 ();
 FILLCELL_X1 FILLER_22_513 ();
 FILLCELL_X16 FILLER_22_519 ();
 FILLCELL_X1 FILLER_22_535 ();
 FILLCELL_X16 FILLER_22_543 ();
 FILLCELL_X4 FILLER_22_559 ();
 FILLCELL_X2 FILLER_22_563 ();
 FILLCELL_X1 FILLER_22_570 ();
 FILLCELL_X1 FILLER_22_592 ();
 FILLCELL_X4 FILLER_22_598 ();
 FILLCELL_X2 FILLER_22_602 ();
 FILLCELL_X1 FILLER_22_604 ();
 FILLCELL_X8 FILLER_22_622 ();
 FILLCELL_X1 FILLER_22_630 ();
 FILLCELL_X8 FILLER_22_632 ();
 FILLCELL_X1 FILLER_22_640 ();
 FILLCELL_X16 FILLER_22_658 ();
 FILLCELL_X2 FILLER_22_674 ();
 FILLCELL_X8 FILLER_22_684 ();
 FILLCELL_X2 FILLER_22_722 ();
 FILLCELL_X8 FILLER_22_731 ();
 FILLCELL_X4 FILLER_22_739 ();
 FILLCELL_X1 FILLER_22_743 ();
 FILLCELL_X1 FILLER_22_751 ();
 FILLCELL_X32 FILLER_22_759 ();
 FILLCELL_X16 FILLER_22_794 ();
 FILLCELL_X4 FILLER_22_810 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X16 FILLER_23_33 ();
 FILLCELL_X8 FILLER_23_49 ();
 FILLCELL_X2 FILLER_23_57 ();
 FILLCELL_X1 FILLER_23_59 ();
 FILLCELL_X2 FILLER_23_91 ();
 FILLCELL_X8 FILLER_23_103 ();
 FILLCELL_X4 FILLER_23_111 ();
 FILLCELL_X2 FILLER_23_115 ();
 FILLCELL_X1 FILLER_23_117 ();
 FILLCELL_X1 FILLER_23_142 ();
 FILLCELL_X16 FILLER_23_160 ();
 FILLCELL_X16 FILLER_23_180 ();
 FILLCELL_X4 FILLER_23_196 ();
 FILLCELL_X1 FILLER_23_200 ();
 FILLCELL_X1 FILLER_23_208 ();
 FILLCELL_X2 FILLER_23_212 ();
 FILLCELL_X1 FILLER_23_214 ();
 FILLCELL_X16 FILLER_23_218 ();
 FILLCELL_X8 FILLER_23_234 ();
 FILLCELL_X1 FILLER_23_242 ();
 FILLCELL_X8 FILLER_23_260 ();
 FILLCELL_X2 FILLER_23_268 ();
 FILLCELL_X1 FILLER_23_270 ();
 FILLCELL_X1 FILLER_23_278 ();
 FILLCELL_X1 FILLER_23_296 ();
 FILLCELL_X2 FILLER_23_304 ();
 FILLCELL_X2 FILLER_23_313 ();
 FILLCELL_X4 FILLER_23_335 ();
 FILLCELL_X8 FILLER_23_347 ();
 FILLCELL_X2 FILLER_23_355 ();
 FILLCELL_X1 FILLER_23_357 ();
 FILLCELL_X4 FILLER_23_376 ();
 FILLCELL_X1 FILLER_23_380 ();
 FILLCELL_X1 FILLER_23_413 ();
 FILLCELL_X16 FILLER_23_421 ();
 FILLCELL_X8 FILLER_23_437 ();
 FILLCELL_X2 FILLER_23_445 ();
 FILLCELL_X8 FILLER_23_467 ();
 FILLCELL_X16 FILLER_23_478 ();
 FILLCELL_X4 FILLER_23_494 ();
 FILLCELL_X2 FILLER_23_498 ();
 FILLCELL_X8 FILLER_23_510 ();
 FILLCELL_X4 FILLER_23_518 ();
 FILLCELL_X2 FILLER_23_522 ();
 FILLCELL_X4 FILLER_23_541 ();
 FILLCELL_X4 FILLER_23_556 ();
 FILLCELL_X8 FILLER_23_562 ();
 FILLCELL_X4 FILLER_23_570 ();
 FILLCELL_X1 FILLER_23_574 ();
 FILLCELL_X2 FILLER_23_581 ();
 FILLCELL_X1 FILLER_23_583 ();
 FILLCELL_X4 FILLER_23_588 ();
 FILLCELL_X2 FILLER_23_592 ();
 FILLCELL_X1 FILLER_23_594 ();
 FILLCELL_X4 FILLER_23_614 ();
 FILLCELL_X2 FILLER_23_625 ();
 FILLCELL_X4 FILLER_23_630 ();
 FILLCELL_X2 FILLER_23_634 ();
 FILLCELL_X8 FILLER_23_640 ();
 FILLCELL_X1 FILLER_23_648 ();
 FILLCELL_X4 FILLER_23_653 ();
 FILLCELL_X1 FILLER_23_657 ();
 FILLCELL_X8 FILLER_23_662 ();
 FILLCELL_X2 FILLER_23_670 ();
 FILLCELL_X1 FILLER_23_672 ();
 FILLCELL_X2 FILLER_23_690 ();
 FILLCELL_X1 FILLER_23_692 ();
 FILLCELL_X8 FILLER_23_710 ();
 FILLCELL_X1 FILLER_23_718 ();
 FILLCELL_X1 FILLER_23_760 ();
 FILLCELL_X4 FILLER_23_768 ();
 FILLCELL_X2 FILLER_23_772 ();
 FILLCELL_X1 FILLER_23_774 ();
 FILLCELL_X2 FILLER_23_788 ();
 FILLCELL_X1 FILLER_23_790 ();
 FILLCELL_X2 FILLER_23_812 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X16 FILLER_24_33 ();
 FILLCELL_X4 FILLER_24_49 ();
 FILLCELL_X1 FILLER_24_53 ();
 FILLCELL_X2 FILLER_24_71 ();
 FILLCELL_X1 FILLER_24_73 ();
 FILLCELL_X8 FILLER_24_77 ();
 FILLCELL_X4 FILLER_24_85 ();
 FILLCELL_X16 FILLER_24_106 ();
 FILLCELL_X2 FILLER_24_122 ();
 FILLCELL_X1 FILLER_24_124 ();
 FILLCELL_X2 FILLER_24_132 ();
 FILLCELL_X8 FILLER_24_137 ();
 FILLCELL_X2 FILLER_24_145 ();
 FILLCELL_X1 FILLER_24_150 ();
 FILLCELL_X32 FILLER_24_154 ();
 FILLCELL_X8 FILLER_24_186 ();
 FILLCELL_X1 FILLER_24_194 ();
 FILLCELL_X2 FILLER_24_212 ();
 FILLCELL_X8 FILLER_24_238 ();
 FILLCELL_X4 FILLER_24_246 ();
 FILLCELL_X8 FILLER_24_253 ();
 FILLCELL_X2 FILLER_24_261 ();
 FILLCELL_X16 FILLER_24_280 ();
 FILLCELL_X2 FILLER_24_303 ();
 FILLCELL_X1 FILLER_24_305 ();
 FILLCELL_X4 FILLER_24_309 ();
 FILLCELL_X1 FILLER_24_313 ();
 FILLCELL_X2 FILLER_24_321 ();
 FILLCELL_X1 FILLER_24_323 ();
 FILLCELL_X8 FILLER_24_331 ();
 FILLCELL_X1 FILLER_24_339 ();
 FILLCELL_X8 FILLER_24_344 ();
 FILLCELL_X4 FILLER_24_352 ();
 FILLCELL_X2 FILLER_24_356 ();
 FILLCELL_X4 FILLER_24_380 ();
 FILLCELL_X2 FILLER_24_384 ();
 FILLCELL_X1 FILLER_24_386 ();
 FILLCELL_X2 FILLER_24_394 ();
 FILLCELL_X4 FILLER_24_399 ();
 FILLCELL_X2 FILLER_24_403 ();
 FILLCELL_X1 FILLER_24_405 ();
 FILLCELL_X8 FILLER_24_427 ();
 FILLCELL_X4 FILLER_24_442 ();
 FILLCELL_X1 FILLER_24_446 ();
 FILLCELL_X1 FILLER_24_462 ();
 FILLCELL_X16 FILLER_24_484 ();
 FILLCELL_X4 FILLER_24_500 ();
 FILLCELL_X2 FILLER_24_518 ();
 FILLCELL_X4 FILLER_24_544 ();
 FILLCELL_X1 FILLER_24_548 ();
 FILLCELL_X2 FILLER_24_568 ();
 FILLCELL_X8 FILLER_24_591 ();
 FILLCELL_X2 FILLER_24_599 ();
 FILLCELL_X1 FILLER_24_601 ();
 FILLCELL_X4 FILLER_24_626 ();
 FILLCELL_X1 FILLER_24_630 ();
 FILLCELL_X4 FILLER_24_673 ();
 FILLCELL_X1 FILLER_24_677 ();
 FILLCELL_X32 FILLER_24_687 ();
 FILLCELL_X2 FILLER_24_719 ();
 FILLCELL_X1 FILLER_24_724 ();
 FILLCELL_X4 FILLER_24_731 ();
 FILLCELL_X4 FILLER_24_742 ();
 FILLCELL_X1 FILLER_24_746 ();
 FILLCELL_X1 FILLER_24_751 ();
 FILLCELL_X2 FILLER_24_758 ();
 FILLCELL_X4 FILLER_24_767 ();
 FILLCELL_X1 FILLER_24_771 ();
 FILLCELL_X16 FILLER_24_789 ();
 FILLCELL_X8 FILLER_24_805 ();
 FILLCELL_X1 FILLER_24_813 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X8 FILLER_25_33 ();
 FILLCELL_X4 FILLER_25_41 ();
 FILLCELL_X2 FILLER_25_45 ();
 FILLCELL_X2 FILLER_25_64 ();
 FILLCELL_X1 FILLER_25_66 ();
 FILLCELL_X8 FILLER_25_71 ();
 FILLCELL_X2 FILLER_25_79 ();
 FILLCELL_X1 FILLER_25_81 ();
 FILLCELL_X1 FILLER_25_86 ();
 FILLCELL_X1 FILLER_25_94 ();
 FILLCELL_X2 FILLER_25_98 ();
 FILLCELL_X2 FILLER_25_107 ();
 FILLCELL_X2 FILLER_25_116 ();
 FILLCELL_X1 FILLER_25_118 ();
 FILLCELL_X8 FILLER_25_136 ();
 FILLCELL_X4 FILLER_25_144 ();
 FILLCELL_X2 FILLER_25_158 ();
 FILLCELL_X1 FILLER_25_160 ();
 FILLCELL_X4 FILLER_25_168 ();
 FILLCELL_X2 FILLER_25_172 ();
 FILLCELL_X2 FILLER_25_181 ();
 FILLCELL_X1 FILLER_25_183 ();
 FILLCELL_X4 FILLER_25_188 ();
 FILLCELL_X2 FILLER_25_192 ();
 FILLCELL_X4 FILLER_25_214 ();
 FILLCELL_X4 FILLER_25_246 ();
 FILLCELL_X2 FILLER_25_250 ();
 FILLCELL_X2 FILLER_25_256 ();
 FILLCELL_X16 FILLER_25_261 ();
 FILLCELL_X2 FILLER_25_277 ();
 FILLCELL_X1 FILLER_25_279 ();
 FILLCELL_X2 FILLER_25_307 ();
 FILLCELL_X16 FILLER_25_316 ();
 FILLCELL_X2 FILLER_25_332 ();
 FILLCELL_X8 FILLER_25_354 ();
 FILLCELL_X2 FILLER_25_362 ();
 FILLCELL_X1 FILLER_25_371 ();
 FILLCELL_X4 FILLER_25_375 ();
 FILLCELL_X4 FILLER_25_403 ();
 FILLCELL_X2 FILLER_25_407 ();
 FILLCELL_X1 FILLER_25_430 ();
 FILLCELL_X16 FILLER_25_465 ();
 FILLCELL_X1 FILLER_25_516 ();
 FILLCELL_X4 FILLER_25_527 ();
 FILLCELL_X1 FILLER_25_531 ();
 FILLCELL_X16 FILLER_25_536 ();
 FILLCELL_X4 FILLER_25_552 ();
 FILLCELL_X2 FILLER_25_556 ();
 FILLCELL_X1 FILLER_25_558 ();
 FILLCELL_X4 FILLER_25_563 ();
 FILLCELL_X2 FILLER_25_575 ();
 FILLCELL_X1 FILLER_25_577 ();
 FILLCELL_X4 FILLER_25_585 ();
 FILLCELL_X2 FILLER_25_597 ();
 FILLCELL_X1 FILLER_25_599 ();
 FILLCELL_X2 FILLER_25_609 ();
 FILLCELL_X16 FILLER_25_613 ();
 FILLCELL_X8 FILLER_25_629 ();
 FILLCELL_X1 FILLER_25_637 ();
 FILLCELL_X16 FILLER_25_642 ();
 FILLCELL_X8 FILLER_25_658 ();
 FILLCELL_X2 FILLER_25_670 ();
 FILLCELL_X1 FILLER_25_672 ();
 FILLCELL_X4 FILLER_25_675 ();
 FILLCELL_X1 FILLER_25_679 ();
 FILLCELL_X1 FILLER_25_682 ();
 FILLCELL_X2 FILLER_25_690 ();
 FILLCELL_X1 FILLER_25_696 ();
 FILLCELL_X2 FILLER_25_700 ();
 FILLCELL_X2 FILLER_25_707 ();
 FILLCELL_X4 FILLER_25_716 ();
 FILLCELL_X8 FILLER_25_724 ();
 FILLCELL_X2 FILLER_25_749 ();
 FILLCELL_X4 FILLER_25_761 ();
 FILLCELL_X2 FILLER_25_765 ();
 FILLCELL_X1 FILLER_25_781 ();
 FILLCELL_X2 FILLER_25_788 ();
 FILLCELL_X1 FILLER_25_790 ();
 FILLCELL_X2 FILLER_25_795 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X16 FILLER_26_33 ();
 FILLCELL_X8 FILLER_26_49 ();
 FILLCELL_X2 FILLER_26_69 ();
 FILLCELL_X1 FILLER_26_71 ();
 FILLCELL_X1 FILLER_26_89 ();
 FILLCELL_X16 FILLER_26_97 ();
 FILLCELL_X8 FILLER_26_113 ();
 FILLCELL_X4 FILLER_26_121 ();
 FILLCELL_X1 FILLER_26_125 ();
 FILLCELL_X1 FILLER_26_130 ();
 FILLCELL_X4 FILLER_26_142 ();
 FILLCELL_X8 FILLER_26_170 ();
 FILLCELL_X1 FILLER_26_178 ();
 FILLCELL_X1 FILLER_26_207 ();
 FILLCELL_X16 FILLER_26_211 ();
 FILLCELL_X4 FILLER_26_241 ();
 FILLCELL_X8 FILLER_26_265 ();
 FILLCELL_X2 FILLER_26_273 ();
 FILLCELL_X1 FILLER_26_275 ();
 FILLCELL_X8 FILLER_26_284 ();
 FILLCELL_X4 FILLER_26_292 ();
 FILLCELL_X2 FILLER_26_296 ();
 FILLCELL_X8 FILLER_26_318 ();
 FILLCELL_X2 FILLER_26_326 ();
 FILLCELL_X1 FILLER_26_335 ();
 FILLCELL_X8 FILLER_26_339 ();
 FILLCELL_X4 FILLER_26_347 ();
 FILLCELL_X4 FILLER_26_356 ();
 FILLCELL_X2 FILLER_26_360 ();
 FILLCELL_X2 FILLER_26_379 ();
 FILLCELL_X8 FILLER_26_388 ();
 FILLCELL_X2 FILLER_26_396 ();
 FILLCELL_X8 FILLER_26_426 ();
 FILLCELL_X2 FILLER_26_434 ();
 FILLCELL_X8 FILLER_26_439 ();
 FILLCELL_X4 FILLER_26_447 ();
 FILLCELL_X4 FILLER_26_454 ();
 FILLCELL_X8 FILLER_26_478 ();
 FILLCELL_X1 FILLER_26_486 ();
 FILLCELL_X8 FILLER_26_508 ();
 FILLCELL_X2 FILLER_26_516 ();
 FILLCELL_X1 FILLER_26_518 ();
 FILLCELL_X4 FILLER_26_528 ();
 FILLCELL_X16 FILLER_26_536 ();
 FILLCELL_X4 FILLER_26_552 ();
 FILLCELL_X1 FILLER_26_567 ();
 FILLCELL_X1 FILLER_26_572 ();
 FILLCELL_X1 FILLER_26_577 ();
 FILLCELL_X1 FILLER_26_585 ();
 FILLCELL_X8 FILLER_26_618 ();
 FILLCELL_X4 FILLER_26_626 ();
 FILLCELL_X1 FILLER_26_630 ();
 FILLCELL_X2 FILLER_26_632 ();
 FILLCELL_X1 FILLER_26_634 ();
 FILLCELL_X4 FILLER_26_639 ();
 FILLCELL_X1 FILLER_26_646 ();
 FILLCELL_X1 FILLER_26_651 ();
 FILLCELL_X2 FILLER_26_663 ();
 FILLCELL_X16 FILLER_26_730 ();
 FILLCELL_X8 FILLER_26_746 ();
 FILLCELL_X4 FILLER_26_754 ();
 FILLCELL_X1 FILLER_26_758 ();
 FILLCELL_X32 FILLER_26_780 ();
 FILLCELL_X2 FILLER_26_812 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X16 FILLER_27_33 ();
 FILLCELL_X16 FILLER_27_66 ();
 FILLCELL_X2 FILLER_27_82 ();
 FILLCELL_X1 FILLER_27_84 ();
 FILLCELL_X1 FILLER_27_88 ();
 FILLCELL_X2 FILLER_27_103 ();
 FILLCELL_X2 FILLER_27_112 ();
 FILLCELL_X1 FILLER_27_114 ();
 FILLCELL_X16 FILLER_27_139 ();
 FILLCELL_X1 FILLER_27_162 ();
 FILLCELL_X1 FILLER_27_171 ();
 FILLCELL_X8 FILLER_27_180 ();
 FILLCELL_X4 FILLER_27_188 ();
 FILLCELL_X2 FILLER_27_192 ();
 FILLCELL_X1 FILLER_27_194 ();
 FILLCELL_X4 FILLER_27_203 ();
 FILLCELL_X8 FILLER_27_211 ();
 FILLCELL_X2 FILLER_27_219 ();
 FILLCELL_X32 FILLER_27_245 ();
 FILLCELL_X4 FILLER_27_277 ();
 FILLCELL_X1 FILLER_27_281 ();
 FILLCELL_X2 FILLER_27_285 ();
 FILLCELL_X1 FILLER_27_287 ();
 FILLCELL_X8 FILLER_27_291 ();
 FILLCELL_X4 FILLER_27_299 ();
 FILLCELL_X4 FILLER_27_307 ();
 FILLCELL_X2 FILLER_27_311 ();
 FILLCELL_X1 FILLER_27_313 ();
 FILLCELL_X1 FILLER_27_321 ();
 FILLCELL_X4 FILLER_27_339 ();
 FILLCELL_X2 FILLER_27_343 ();
 FILLCELL_X1 FILLER_27_345 ();
 FILLCELL_X1 FILLER_27_353 ();
 FILLCELL_X2 FILLER_27_359 ();
 FILLCELL_X4 FILLER_27_368 ();
 FILLCELL_X1 FILLER_27_372 ();
 FILLCELL_X16 FILLER_27_377 ();
 FILLCELL_X2 FILLER_27_393 ();
 FILLCELL_X1 FILLER_27_395 ();
 FILLCELL_X32 FILLER_27_406 ();
 FILLCELL_X8 FILLER_27_438 ();
 FILLCELL_X4 FILLER_27_446 ();
 FILLCELL_X1 FILLER_27_450 ();
 FILLCELL_X4 FILLER_27_454 ();
 FILLCELL_X32 FILLER_27_462 ();
 FILLCELL_X4 FILLER_27_494 ();
 FILLCELL_X2 FILLER_27_498 ();
 FILLCELL_X1 FILLER_27_503 ();
 FILLCELL_X1 FILLER_27_528 ();
 FILLCELL_X2 FILLER_27_563 ();
 FILLCELL_X16 FILLER_27_582 ();
 FILLCELL_X8 FILLER_27_598 ();
 FILLCELL_X2 FILLER_27_606 ();
 FILLCELL_X1 FILLER_27_627 ();
 FILLCELL_X8 FILLER_27_669 ();
 FILLCELL_X1 FILLER_27_677 ();
 FILLCELL_X2 FILLER_27_683 ();
 FILLCELL_X1 FILLER_27_685 ();
 FILLCELL_X16 FILLER_27_694 ();
 FILLCELL_X8 FILLER_27_710 ();
 FILLCELL_X2 FILLER_27_718 ();
 FILLCELL_X4 FILLER_27_723 ();
 FILLCELL_X1 FILLER_27_727 ();
 FILLCELL_X2 FILLER_27_757 ();
 FILLCELL_X1 FILLER_27_759 ();
 FILLCELL_X1 FILLER_27_765 ();
 FILLCELL_X16 FILLER_27_783 ();
 FILLCELL_X8 FILLER_27_799 ();
 FILLCELL_X4 FILLER_27_807 ();
 FILLCELL_X2 FILLER_27_811 ();
 FILLCELL_X1 FILLER_27_813 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X16 FILLER_28_65 ();
 FILLCELL_X4 FILLER_28_81 ();
 FILLCELL_X2 FILLER_28_85 ();
 FILLCELL_X16 FILLER_28_94 ();
 FILLCELL_X1 FILLER_28_110 ();
 FILLCELL_X8 FILLER_28_125 ();
 FILLCELL_X2 FILLER_28_133 ();
 FILLCELL_X1 FILLER_28_135 ();
 FILLCELL_X2 FILLER_28_152 ();
 FILLCELL_X8 FILLER_28_161 ();
 FILLCELL_X2 FILLER_28_186 ();
 FILLCELL_X1 FILLER_28_205 ();
 FILLCELL_X1 FILLER_28_223 ();
 FILLCELL_X1 FILLER_28_238 ();
 FILLCELL_X8 FILLER_28_246 ();
 FILLCELL_X4 FILLER_28_254 ();
 FILLCELL_X2 FILLER_28_265 ();
 FILLCELL_X16 FILLER_28_302 ();
 FILLCELL_X2 FILLER_28_330 ();
 FILLCELL_X1 FILLER_28_332 ();
 FILLCELL_X1 FILLER_28_355 ();
 FILLCELL_X1 FILLER_28_373 ();
 FILLCELL_X2 FILLER_28_377 ();
 FILLCELL_X8 FILLER_28_382 ();
 FILLCELL_X4 FILLER_28_390 ();
 FILLCELL_X16 FILLER_28_411 ();
 FILLCELL_X4 FILLER_28_427 ();
 FILLCELL_X2 FILLER_28_431 ();
 FILLCELL_X1 FILLER_28_433 ();
 FILLCELL_X4 FILLER_28_448 ();
 FILLCELL_X2 FILLER_28_452 ();
 FILLCELL_X1 FILLER_28_458 ();
 FILLCELL_X4 FILLER_28_462 ();
 FILLCELL_X2 FILLER_28_466 ();
 FILLCELL_X1 FILLER_28_468 ();
 FILLCELL_X8 FILLER_28_476 ();
 FILLCELL_X1 FILLER_28_484 ();
 FILLCELL_X8 FILLER_28_489 ();
 FILLCELL_X4 FILLER_28_497 ();
 FILLCELL_X2 FILLER_28_501 ();
 FILLCELL_X4 FILLER_28_533 ();
 FILLCELL_X2 FILLER_28_537 ();
 FILLCELL_X4 FILLER_28_546 ();
 FILLCELL_X2 FILLER_28_550 ();
 FILLCELL_X8 FILLER_28_563 ();
 FILLCELL_X2 FILLER_28_571 ();
 FILLCELL_X1 FILLER_28_573 ();
 FILLCELL_X8 FILLER_28_578 ();
 FILLCELL_X2 FILLER_28_586 ();
 FILLCELL_X1 FILLER_28_588 ();
 FILLCELL_X4 FILLER_28_598 ();
 FILLCELL_X1 FILLER_28_602 ();
 FILLCELL_X8 FILLER_28_617 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X4 FILLER_28_632 ();
 FILLCELL_X1 FILLER_28_636 ();
 FILLCELL_X8 FILLER_28_640 ();
 FILLCELL_X4 FILLER_28_648 ();
 FILLCELL_X4 FILLER_28_660 ();
 FILLCELL_X16 FILLER_28_669 ();
 FILLCELL_X8 FILLER_28_685 ();
 FILLCELL_X2 FILLER_28_700 ();
 FILLCELL_X4 FILLER_28_709 ();
 FILLCELL_X8 FILLER_28_716 ();
 FILLCELL_X2 FILLER_28_724 ();
 FILLCELL_X1 FILLER_28_726 ();
 FILLCELL_X2 FILLER_28_744 ();
 FILLCELL_X1 FILLER_28_753 ();
 FILLCELL_X8 FILLER_28_761 ();
 FILLCELL_X2 FILLER_28_769 ();
 FILLCELL_X1 FILLER_28_774 ();
 FILLCELL_X1 FILLER_28_778 ();
 FILLCELL_X1 FILLER_28_783 ();
 FILLCELL_X1 FILLER_28_787 ();
 FILLCELL_X8 FILLER_28_802 ();
 FILLCELL_X4 FILLER_28_810 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X8 FILLER_29_33 ();
 FILLCELL_X4 FILLER_29_48 ();
 FILLCELL_X4 FILLER_29_69 ();
 FILLCELL_X1 FILLER_29_73 ();
 FILLCELL_X2 FILLER_29_81 ();
 FILLCELL_X1 FILLER_29_83 ();
 FILLCELL_X8 FILLER_29_91 ();
 FILLCELL_X4 FILLER_29_99 ();
 FILLCELL_X1 FILLER_29_103 ();
 FILLCELL_X1 FILLER_29_108 ();
 FILLCELL_X8 FILLER_29_113 ();
 FILLCELL_X1 FILLER_29_125 ();
 FILLCELL_X2 FILLER_29_129 ();
 FILLCELL_X2 FILLER_29_138 ();
 FILLCELL_X2 FILLER_29_157 ();
 FILLCELL_X1 FILLER_29_159 ();
 FILLCELL_X32 FILLER_29_167 ();
 FILLCELL_X16 FILLER_29_199 ();
 FILLCELL_X8 FILLER_29_215 ();
 FILLCELL_X4 FILLER_29_223 ();
 FILLCELL_X1 FILLER_29_227 ();
 FILLCELL_X4 FILLER_29_242 ();
 FILLCELL_X2 FILLER_29_246 ();
 FILLCELL_X1 FILLER_29_248 ();
 FILLCELL_X4 FILLER_29_254 ();
 FILLCELL_X2 FILLER_29_258 ();
 FILLCELL_X4 FILLER_29_285 ();
 FILLCELL_X1 FILLER_29_289 ();
 FILLCELL_X1 FILLER_29_298 ();
 FILLCELL_X1 FILLER_29_316 ();
 FILLCELL_X1 FILLER_29_334 ();
 FILLCELL_X4 FILLER_29_342 ();
 FILLCELL_X2 FILLER_29_346 ();
 FILLCELL_X1 FILLER_29_348 ();
 FILLCELL_X4 FILLER_29_357 ();
 FILLCELL_X1 FILLER_29_361 ();
 FILLCELL_X4 FILLER_29_365 ();
 FILLCELL_X2 FILLER_29_369 ();
 FILLCELL_X1 FILLER_29_371 ();
 FILLCELL_X8 FILLER_29_396 ();
 FILLCELL_X4 FILLER_29_404 ();
 FILLCELL_X2 FILLER_29_408 ();
 FILLCELL_X2 FILLER_29_434 ();
 FILLCELL_X4 FILLER_29_470 ();
 FILLCELL_X2 FILLER_29_474 ();
 FILLCELL_X2 FILLER_29_500 ();
 FILLCELL_X4 FILLER_29_509 ();
 FILLCELL_X1 FILLER_29_513 ();
 FILLCELL_X16 FILLER_29_531 ();
 FILLCELL_X1 FILLER_29_547 ();
 FILLCELL_X2 FILLER_29_567 ();
 FILLCELL_X2 FILLER_29_586 ();
 FILLCELL_X1 FILLER_29_588 ();
 FILLCELL_X2 FILLER_29_606 ();
 FILLCELL_X1 FILLER_29_608 ();
 FILLCELL_X32 FILLER_29_614 ();
 FILLCELL_X4 FILLER_29_646 ();
 FILLCELL_X2 FILLER_29_655 ();
 FILLCELL_X1 FILLER_29_657 ();
 FILLCELL_X4 FILLER_29_679 ();
 FILLCELL_X4 FILLER_29_720 ();
 FILLCELL_X1 FILLER_29_727 ();
 FILLCELL_X2 FILLER_29_748 ();
 FILLCELL_X1 FILLER_29_750 ();
 FILLCELL_X2 FILLER_29_762 ();
 FILLCELL_X4 FILLER_29_781 ();
 FILLCELL_X2 FILLER_29_785 ();
 FILLCELL_X1 FILLER_29_792 ();
 FILLCELL_X1 FILLER_29_796 ();
 FILLCELL_X16 FILLER_30_1 ();
 FILLCELL_X8 FILLER_30_17 ();
 FILLCELL_X4 FILLER_30_25 ();
 FILLCELL_X1 FILLER_30_29 ();
 FILLCELL_X8 FILLER_30_47 ();
 FILLCELL_X2 FILLER_30_71 ();
 FILLCELL_X1 FILLER_30_73 ();
 FILLCELL_X2 FILLER_30_95 ();
 FILLCELL_X1 FILLER_30_97 ();
 FILLCELL_X1 FILLER_30_115 ();
 FILLCELL_X1 FILLER_30_145 ();
 FILLCELL_X2 FILLER_30_156 ();
 FILLCELL_X8 FILLER_30_172 ();
 FILLCELL_X1 FILLER_30_180 ();
 FILLCELL_X4 FILLER_30_186 ();
 FILLCELL_X2 FILLER_30_190 ();
 FILLCELL_X1 FILLER_30_192 ();
 FILLCELL_X8 FILLER_30_197 ();
 FILLCELL_X4 FILLER_30_229 ();
 FILLCELL_X2 FILLER_30_233 ();
 FILLCELL_X1 FILLER_30_235 ();
 FILLCELL_X1 FILLER_30_248 ();
 FILLCELL_X1 FILLER_30_270 ();
 FILLCELL_X2 FILLER_30_274 ();
 FILLCELL_X1 FILLER_30_276 ();
 FILLCELL_X4 FILLER_30_289 ();
 FILLCELL_X2 FILLER_30_300 ();
 FILLCELL_X4 FILLER_30_306 ();
 FILLCELL_X2 FILLER_30_310 ();
 FILLCELL_X2 FILLER_30_315 ();
 FILLCELL_X1 FILLER_30_317 ();
 FILLCELL_X2 FILLER_30_321 ();
 FILLCELL_X1 FILLER_30_323 ();
 FILLCELL_X4 FILLER_30_329 ();
 FILLCELL_X1 FILLER_30_333 ();
 FILLCELL_X2 FILLER_30_348 ();
 FILLCELL_X1 FILLER_30_350 ();
 FILLCELL_X8 FILLER_30_358 ();
 FILLCELL_X4 FILLER_30_366 ();
 FILLCELL_X2 FILLER_30_370 ();
 FILLCELL_X1 FILLER_30_372 ();
 FILLCELL_X1 FILLER_30_377 ();
 FILLCELL_X1 FILLER_30_385 ();
 FILLCELL_X16 FILLER_30_400 ();
 FILLCELL_X2 FILLER_30_416 ();
 FILLCELL_X1 FILLER_30_418 ();
 FILLCELL_X1 FILLER_30_426 ();
 FILLCELL_X8 FILLER_30_430 ();
 FILLCELL_X4 FILLER_30_438 ();
 FILLCELL_X1 FILLER_30_442 ();
 FILLCELL_X4 FILLER_30_446 ();
 FILLCELL_X2 FILLER_30_450 ();
 FILLCELL_X8 FILLER_30_455 ();
 FILLCELL_X4 FILLER_30_463 ();
 FILLCELL_X2 FILLER_30_467 ();
 FILLCELL_X8 FILLER_30_476 ();
 FILLCELL_X4 FILLER_30_484 ();
 FILLCELL_X1 FILLER_30_488 ();
 FILLCELL_X2 FILLER_30_492 ();
 FILLCELL_X16 FILLER_30_499 ();
 FILLCELL_X8 FILLER_30_515 ();
 FILLCELL_X1 FILLER_30_527 ();
 FILLCELL_X4 FILLER_30_539 ();
 FILLCELL_X2 FILLER_30_543 ();
 FILLCELL_X4 FILLER_30_549 ();
 FILLCELL_X2 FILLER_30_553 ();
 FILLCELL_X1 FILLER_30_555 ();
 FILLCELL_X8 FILLER_30_561 ();
 FILLCELL_X4 FILLER_30_569 ();
 FILLCELL_X2 FILLER_30_573 ();
 FILLCELL_X1 FILLER_30_575 ();
 FILLCELL_X4 FILLER_30_585 ();
 FILLCELL_X4 FILLER_30_597 ();
 FILLCELL_X2 FILLER_30_624 ();
 FILLCELL_X1 FILLER_30_626 ();
 FILLCELL_X1 FILLER_30_632 ();
 FILLCELL_X1 FILLER_30_644 ();
 FILLCELL_X4 FILLER_30_652 ();
 FILLCELL_X4 FILLER_30_660 ();
 FILLCELL_X8 FILLER_30_668 ();
 FILLCELL_X2 FILLER_30_676 ();
 FILLCELL_X4 FILLER_30_683 ();
 FILLCELL_X1 FILLER_30_687 ();
 FILLCELL_X1 FILLER_30_692 ();
 FILLCELL_X2 FILLER_30_697 ();
 FILLCELL_X8 FILLER_30_706 ();
 FILLCELL_X2 FILLER_30_714 ();
 FILLCELL_X16 FILLER_30_736 ();
 FILLCELL_X8 FILLER_30_752 ();
 FILLCELL_X4 FILLER_30_760 ();
 FILLCELL_X1 FILLER_30_764 ();
 FILLCELL_X1 FILLER_30_777 ();
 FILLCELL_X2 FILLER_30_790 ();
 FILLCELL_X16 FILLER_30_797 ();
 FILLCELL_X1 FILLER_30_813 ();
 FILLCELL_X8 FILLER_31_1 ();
 FILLCELL_X1 FILLER_31_9 ();
 FILLCELL_X16 FILLER_31_17 ();
 FILLCELL_X4 FILLER_31_33 ();
 FILLCELL_X2 FILLER_31_47 ();
 FILLCELL_X1 FILLER_31_49 ();
 FILLCELL_X16 FILLER_31_86 ();
 FILLCELL_X4 FILLER_31_102 ();
 FILLCELL_X4 FILLER_31_114 ();
 FILLCELL_X8 FILLER_31_126 ();
 FILLCELL_X4 FILLER_31_134 ();
 FILLCELL_X2 FILLER_31_138 ();
 FILLCELL_X1 FILLER_31_140 ();
 FILLCELL_X2 FILLER_31_148 ();
 FILLCELL_X1 FILLER_31_150 ();
 FILLCELL_X8 FILLER_31_167 ();
 FILLCELL_X4 FILLER_31_175 ();
 FILLCELL_X2 FILLER_31_183 ();
 FILLCELL_X1 FILLER_31_185 ();
 FILLCELL_X4 FILLER_31_194 ();
 FILLCELL_X2 FILLER_31_198 ();
 FILLCELL_X1 FILLER_31_200 ();
 FILLCELL_X4 FILLER_31_225 ();
 FILLCELL_X2 FILLER_31_229 ();
 FILLCELL_X1 FILLER_31_236 ();
 FILLCELL_X2 FILLER_31_275 ();
 FILLCELL_X1 FILLER_31_297 ();
 FILLCELL_X1 FILLER_31_301 ();
 FILLCELL_X4 FILLER_31_305 ();
 FILLCELL_X8 FILLER_31_313 ();
 FILLCELL_X4 FILLER_31_324 ();
 FILLCELL_X1 FILLER_31_345 ();
 FILLCELL_X8 FILLER_31_379 ();
 FILLCELL_X4 FILLER_31_401 ();
 FILLCELL_X2 FILLER_31_405 ();
 FILLCELL_X8 FILLER_31_425 ();
 FILLCELL_X2 FILLER_31_433 ();
 FILLCELL_X1 FILLER_31_435 ();
 FILLCELL_X2 FILLER_31_440 ();
 FILLCELL_X4 FILLER_31_445 ();
 FILLCELL_X4 FILLER_31_453 ();
 FILLCELL_X1 FILLER_31_457 ();
 FILLCELL_X1 FILLER_31_461 ();
 FILLCELL_X2 FILLER_31_466 ();
 FILLCELL_X1 FILLER_31_468 ();
 FILLCELL_X4 FILLER_31_479 ();
 FILLCELL_X2 FILLER_31_483 ();
 FILLCELL_X8 FILLER_31_504 ();
 FILLCELL_X1 FILLER_31_516 ();
 FILLCELL_X4 FILLER_31_524 ();
 FILLCELL_X2 FILLER_31_535 ();
 FILLCELL_X4 FILLER_31_543 ();
 FILLCELL_X2 FILLER_31_547 ();
 FILLCELL_X2 FILLER_31_556 ();
 FILLCELL_X2 FILLER_31_563 ();
 FILLCELL_X1 FILLER_31_565 ();
 FILLCELL_X8 FILLER_31_568 ();
 FILLCELL_X2 FILLER_31_576 ();
 FILLCELL_X1 FILLER_31_578 ();
 FILLCELL_X2 FILLER_31_618 ();
 FILLCELL_X1 FILLER_31_620 ();
 FILLCELL_X8 FILLER_31_640 ();
 FILLCELL_X4 FILLER_31_661 ();
 FILLCELL_X1 FILLER_31_665 ();
 FILLCELL_X2 FILLER_31_671 ();
 FILLCELL_X1 FILLER_31_673 ();
 FILLCELL_X2 FILLER_31_679 ();
 FILLCELL_X2 FILLER_31_686 ();
 FILLCELL_X1 FILLER_31_688 ();
 FILLCELL_X16 FILLER_31_697 ();
 FILLCELL_X8 FILLER_31_713 ();
 FILLCELL_X2 FILLER_31_721 ();
 FILLCELL_X1 FILLER_31_723 ();
 FILLCELL_X1 FILLER_31_731 ();
 FILLCELL_X1 FILLER_31_743 ();
 FILLCELL_X2 FILLER_31_748 ();
 FILLCELL_X1 FILLER_31_750 ();
 FILLCELL_X4 FILLER_31_755 ();
 FILLCELL_X4 FILLER_31_766 ();
 FILLCELL_X1 FILLER_31_780 ();
 FILLCELL_X2 FILLER_31_788 ();
 FILLCELL_X1 FILLER_31_790 ();
 FILLCELL_X16 FILLER_31_796 ();
 FILLCELL_X2 FILLER_31_812 ();
 FILLCELL_X16 FILLER_32_1 ();
 FILLCELL_X8 FILLER_32_17 ();
 FILLCELL_X2 FILLER_32_25 ();
 FILLCELL_X1 FILLER_32_27 ();
 FILLCELL_X4 FILLER_32_53 ();
 FILLCELL_X2 FILLER_32_57 ();
 FILLCELL_X1 FILLER_32_59 ();
 FILLCELL_X16 FILLER_32_68 ();
 FILLCELL_X2 FILLER_32_84 ();
 FILLCELL_X8 FILLER_32_113 ();
 FILLCELL_X2 FILLER_32_121 ();
 FILLCELL_X1 FILLER_32_123 ();
 FILLCELL_X8 FILLER_32_131 ();
 FILLCELL_X2 FILLER_32_163 ();
 FILLCELL_X1 FILLER_32_165 ();
 FILLCELL_X8 FILLER_32_205 ();
 FILLCELL_X2 FILLER_32_213 ();
 FILLCELL_X1 FILLER_32_215 ();
 FILLCELL_X2 FILLER_32_232 ();
 FILLCELL_X8 FILLER_32_251 ();
 FILLCELL_X2 FILLER_32_259 ();
 FILLCELL_X1 FILLER_32_261 ();
 FILLCELL_X2 FILLER_32_267 ();
 FILLCELL_X1 FILLER_32_275 ();
 FILLCELL_X8 FILLER_32_281 ();
 FILLCELL_X2 FILLER_32_289 ();
 FILLCELL_X1 FILLER_32_291 ();
 FILLCELL_X2 FILLER_32_304 ();
 FILLCELL_X1 FILLER_32_323 ();
 FILLCELL_X2 FILLER_32_340 ();
 FILLCELL_X16 FILLER_32_360 ();
 FILLCELL_X2 FILLER_32_376 ();
 FILLCELL_X16 FILLER_32_390 ();
 FILLCELL_X4 FILLER_32_406 ();
 FILLCELL_X2 FILLER_32_427 ();
 FILLCELL_X2 FILLER_32_480 ();
 FILLCELL_X2 FILLER_32_499 ();
 FILLCELL_X2 FILLER_32_527 ();
 FILLCELL_X2 FILLER_32_537 ();
 FILLCELL_X1 FILLER_32_539 ();
 FILLCELL_X4 FILLER_32_549 ();
 FILLCELL_X2 FILLER_32_553 ();
 FILLCELL_X2 FILLER_32_574 ();
 FILLCELL_X4 FILLER_32_580 ();
 FILLCELL_X1 FILLER_32_584 ();
 FILLCELL_X4 FILLER_32_594 ();
 FILLCELL_X1 FILLER_32_614 ();
 FILLCELL_X8 FILLER_32_622 ();
 FILLCELL_X1 FILLER_32_630 ();
 FILLCELL_X2 FILLER_32_632 ();
 FILLCELL_X2 FILLER_32_655 ();
 FILLCELL_X1 FILLER_32_657 ();
 FILLCELL_X4 FILLER_32_672 ();
 FILLCELL_X16 FILLER_32_710 ();
 FILLCELL_X4 FILLER_32_726 ();
 FILLCELL_X2 FILLER_32_730 ();
 FILLCELL_X1 FILLER_32_732 ();
 FILLCELL_X4 FILLER_32_757 ();
 FILLCELL_X2 FILLER_32_761 ();
 FILLCELL_X4 FILLER_32_780 ();
 FILLCELL_X2 FILLER_32_784 ();
 FILLCELL_X1 FILLER_32_793 ();
 FILLCELL_X8 FILLER_32_804 ();
 FILLCELL_X2 FILLER_32_812 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X16 FILLER_33_33 ();
 FILLCELL_X2 FILLER_33_49 ();
 FILLCELL_X1 FILLER_33_51 ();
 FILLCELL_X4 FILLER_33_69 ();
 FILLCELL_X2 FILLER_33_73 ();
 FILLCELL_X1 FILLER_33_75 ();
 FILLCELL_X16 FILLER_33_90 ();
 FILLCELL_X8 FILLER_33_106 ();
 FILLCELL_X2 FILLER_33_114 ();
 FILLCELL_X1 FILLER_33_123 ();
 FILLCELL_X4 FILLER_33_153 ();
 FILLCELL_X1 FILLER_33_157 ();
 FILLCELL_X4 FILLER_33_165 ();
 FILLCELL_X2 FILLER_33_169 ();
 FILLCELL_X4 FILLER_33_181 ();
 FILLCELL_X1 FILLER_33_189 ();
 FILLCELL_X4 FILLER_33_193 ();
 FILLCELL_X1 FILLER_33_197 ();
 FILLCELL_X8 FILLER_33_217 ();
 FILLCELL_X4 FILLER_33_225 ();
 FILLCELL_X2 FILLER_33_229 ();
 FILLCELL_X16 FILLER_33_262 ();
 FILLCELL_X8 FILLER_33_278 ();
 FILLCELL_X4 FILLER_33_286 ();
 FILLCELL_X2 FILLER_33_290 ();
 FILLCELL_X8 FILLER_33_309 ();
 FILLCELL_X4 FILLER_33_317 ();
 FILLCELL_X1 FILLER_33_321 ();
 FILLCELL_X8 FILLER_33_332 ();
 FILLCELL_X8 FILLER_33_347 ();
 FILLCELL_X4 FILLER_33_355 ();
 FILLCELL_X2 FILLER_33_359 ();
 FILLCELL_X1 FILLER_33_365 ();
 FILLCELL_X4 FILLER_33_374 ();
 FILLCELL_X2 FILLER_33_385 ();
 FILLCELL_X2 FILLER_33_394 ();
 FILLCELL_X1 FILLER_33_396 ();
 FILLCELL_X2 FILLER_33_404 ();
 FILLCELL_X1 FILLER_33_406 ();
 FILLCELL_X4 FILLER_33_412 ();
 FILLCELL_X2 FILLER_33_427 ();
 FILLCELL_X2 FILLER_33_440 ();
 FILLCELL_X1 FILLER_33_442 ();
 FILLCELL_X1 FILLER_33_451 ();
 FILLCELL_X8 FILLER_33_455 ();
 FILLCELL_X4 FILLER_33_463 ();
 FILLCELL_X2 FILLER_33_467 ();
 FILLCELL_X2 FILLER_33_476 ();
 FILLCELL_X4 FILLER_33_483 ();
 FILLCELL_X1 FILLER_33_487 ();
 FILLCELL_X1 FILLER_33_491 ();
 FILLCELL_X1 FILLER_33_495 ();
 FILLCELL_X8 FILLER_33_503 ();
 FILLCELL_X2 FILLER_33_511 ();
 FILLCELL_X4 FILLER_33_518 ();
 FILLCELL_X2 FILLER_33_522 ();
 FILLCELL_X4 FILLER_33_561 ();
 FILLCELL_X2 FILLER_33_565 ();
 FILLCELL_X1 FILLER_33_588 ();
 FILLCELL_X2 FILLER_33_600 ();
 FILLCELL_X1 FILLER_33_608 ();
 FILLCELL_X8 FILLER_33_626 ();
 FILLCELL_X4 FILLER_33_634 ();
 FILLCELL_X2 FILLER_33_638 ();
 FILLCELL_X1 FILLER_33_640 ();
 FILLCELL_X8 FILLER_33_665 ();
 FILLCELL_X4 FILLER_33_673 ();
 FILLCELL_X1 FILLER_33_677 ();
 FILLCELL_X2 FILLER_33_682 ();
 FILLCELL_X1 FILLER_33_684 ();
 FILLCELL_X4 FILLER_33_694 ();
 FILLCELL_X4 FILLER_33_702 ();
 FILLCELL_X1 FILLER_33_706 ();
 FILLCELL_X8 FILLER_33_716 ();
 FILLCELL_X4 FILLER_33_724 ();
 FILLCELL_X1 FILLER_33_728 ();
 FILLCELL_X2 FILLER_33_734 ();
 FILLCELL_X8 FILLER_33_746 ();
 FILLCELL_X4 FILLER_33_754 ();
 FILLCELL_X4 FILLER_33_765 ();
 FILLCELL_X4 FILLER_33_792 ();
 FILLCELL_X1 FILLER_33_796 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X4 FILLER_34_33 ();
 FILLCELL_X1 FILLER_34_37 ();
 FILLCELL_X1 FILLER_34_46 ();
 FILLCELL_X8 FILLER_34_64 ();
 FILLCELL_X4 FILLER_34_72 ();
 FILLCELL_X2 FILLER_34_76 ();
 FILLCELL_X8 FILLER_34_92 ();
 FILLCELL_X4 FILLER_34_100 ();
 FILLCELL_X1 FILLER_34_104 ();
 FILLCELL_X8 FILLER_34_133 ();
 FILLCELL_X2 FILLER_34_141 ();
 FILLCELL_X4 FILLER_34_159 ();
 FILLCELL_X2 FILLER_34_163 ();
 FILLCELL_X1 FILLER_34_174 ();
 FILLCELL_X4 FILLER_34_192 ();
 FILLCELL_X1 FILLER_34_196 ();
 FILLCELL_X8 FILLER_34_217 ();
 FILLCELL_X2 FILLER_34_225 ();
 FILLCELL_X1 FILLER_34_227 ();
 FILLCELL_X2 FILLER_34_252 ();
 FILLCELL_X8 FILLER_34_275 ();
 FILLCELL_X2 FILLER_34_283 ();
 FILLCELL_X1 FILLER_34_285 ();
 FILLCELL_X4 FILLER_34_307 ();
 FILLCELL_X4 FILLER_34_328 ();
 FILLCELL_X2 FILLER_34_332 ();
 FILLCELL_X2 FILLER_34_351 ();
 FILLCELL_X1 FILLER_34_382 ();
 FILLCELL_X2 FILLER_34_397 ();
 FILLCELL_X1 FILLER_34_399 ();
 FILLCELL_X4 FILLER_34_428 ();
 FILLCELL_X2 FILLER_34_432 ();
 FILLCELL_X2 FILLER_34_444 ();
 FILLCELL_X1 FILLER_34_446 ();
 FILLCELL_X1 FILLER_34_452 ();
 FILLCELL_X2 FILLER_34_456 ();
 FILLCELL_X1 FILLER_34_458 ();
 FILLCELL_X16 FILLER_34_466 ();
 FILLCELL_X4 FILLER_34_482 ();
 FILLCELL_X2 FILLER_34_486 ();
 FILLCELL_X1 FILLER_34_493 ();
 FILLCELL_X8 FILLER_34_499 ();
 FILLCELL_X1 FILLER_34_507 ();
 FILLCELL_X2 FILLER_34_518 ();
 FILLCELL_X8 FILLER_34_525 ();
 FILLCELL_X4 FILLER_34_533 ();
 FILLCELL_X1 FILLER_34_537 ();
 FILLCELL_X1 FILLER_34_559 ();
 FILLCELL_X4 FILLER_34_594 ();
 FILLCELL_X2 FILLER_34_598 ();
 FILLCELL_X2 FILLER_34_607 ();
 FILLCELL_X1 FILLER_34_611 ();
 FILLCELL_X4 FILLER_34_617 ();
 FILLCELL_X2 FILLER_34_621 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X16 FILLER_34_632 ();
 FILLCELL_X2 FILLER_34_648 ();
 FILLCELL_X1 FILLER_34_650 ();
 FILLCELL_X8 FILLER_34_656 ();
 FILLCELL_X4 FILLER_34_664 ();
 FILLCELL_X2 FILLER_34_668 ();
 FILLCELL_X1 FILLER_34_670 ();
 FILLCELL_X4 FILLER_34_685 ();
 FILLCELL_X2 FILLER_34_689 ();
 FILLCELL_X1 FILLER_34_724 ();
 FILLCELL_X2 FILLER_34_734 ();
 FILLCELL_X1 FILLER_34_736 ();
 FILLCELL_X2 FILLER_34_744 ();
 FILLCELL_X1 FILLER_34_746 ();
 FILLCELL_X1 FILLER_34_771 ();
 FILLCELL_X32 FILLER_34_774 ();
 FILLCELL_X8 FILLER_34_806 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X4 FILLER_35_33 ();
 FILLCELL_X1 FILLER_35_37 ();
 FILLCELL_X2 FILLER_35_42 ();
 FILLCELL_X2 FILLER_35_83 ();
 FILLCELL_X2 FILLER_35_116 ();
 FILLCELL_X8 FILLER_35_123 ();
 FILLCELL_X4 FILLER_35_131 ();
 FILLCELL_X2 FILLER_35_135 ();
 FILLCELL_X2 FILLER_35_141 ();
 FILLCELL_X4 FILLER_35_147 ();
 FILLCELL_X16 FILLER_35_161 ();
 FILLCELL_X8 FILLER_35_177 ();
 FILLCELL_X2 FILLER_35_196 ();
 FILLCELL_X1 FILLER_35_198 ();
 FILLCELL_X2 FILLER_35_202 ();
 FILLCELL_X1 FILLER_35_204 ();
 FILLCELL_X4 FILLER_35_208 ();
 FILLCELL_X1 FILLER_35_212 ();
 FILLCELL_X32 FILLER_35_220 ();
 FILLCELL_X8 FILLER_35_252 ();
 FILLCELL_X1 FILLER_35_260 ();
 FILLCELL_X1 FILLER_35_264 ();
 FILLCELL_X4 FILLER_35_279 ();
 FILLCELL_X2 FILLER_35_283 ();
 FILLCELL_X2 FILLER_35_309 ();
 FILLCELL_X1 FILLER_35_311 ();
 FILLCELL_X16 FILLER_35_319 ();
 FILLCELL_X4 FILLER_35_335 ();
 FILLCELL_X2 FILLER_35_339 ();
 FILLCELL_X16 FILLER_35_349 ();
 FILLCELL_X8 FILLER_35_365 ();
 FILLCELL_X16 FILLER_35_390 ();
 FILLCELL_X8 FILLER_35_406 ();
 FILLCELL_X4 FILLER_35_414 ();
 FILLCELL_X2 FILLER_35_418 ();
 FILLCELL_X1 FILLER_35_420 ();
 FILLCELL_X2 FILLER_35_425 ();
 FILLCELL_X1 FILLER_35_431 ();
 FILLCELL_X2 FILLER_35_435 ();
 FILLCELL_X4 FILLER_35_442 ();
 FILLCELL_X2 FILLER_35_446 ();
 FILLCELL_X2 FILLER_35_453 ();
 FILLCELL_X1 FILLER_35_455 ();
 FILLCELL_X8 FILLER_35_473 ();
 FILLCELL_X4 FILLER_35_489 ();
 FILLCELL_X2 FILLER_35_493 ();
 FILLCELL_X2 FILLER_35_505 ();
 FILLCELL_X16 FILLER_35_536 ();
 FILLCELL_X8 FILLER_35_552 ();
 FILLCELL_X1 FILLER_35_560 ();
 FILLCELL_X2 FILLER_35_566 ();
 FILLCELL_X1 FILLER_35_568 ();
 FILLCELL_X2 FILLER_35_579 ();
 FILLCELL_X1 FILLER_35_581 ();
 FILLCELL_X2 FILLER_35_606 ();
 FILLCELL_X4 FILLER_35_631 ();
 FILLCELL_X2 FILLER_35_642 ();
 FILLCELL_X2 FILLER_35_653 ();
 FILLCELL_X2 FILLER_35_670 ();
 FILLCELL_X1 FILLER_35_689 ();
 FILLCELL_X2 FILLER_35_704 ();
 FILLCELL_X1 FILLER_35_706 ();
 FILLCELL_X8 FILLER_35_711 ();
 FILLCELL_X4 FILLER_35_719 ();
 FILLCELL_X1 FILLER_35_723 ();
 FILLCELL_X1 FILLER_35_731 ();
 FILLCELL_X8 FILLER_35_749 ();
 FILLCELL_X2 FILLER_35_757 ();
 FILLCELL_X1 FILLER_35_759 ();
 FILLCELL_X4 FILLER_35_764 ();
 FILLCELL_X4 FILLER_35_771 ();
 FILLCELL_X1 FILLER_35_775 ();
 FILLCELL_X2 FILLER_35_783 ();
 FILLCELL_X4 FILLER_35_792 ();
 FILLCELL_X1 FILLER_35_796 ();
 FILLCELL_X16 FILLER_36_1 ();
 FILLCELL_X8 FILLER_36_17 ();
 FILLCELL_X2 FILLER_36_25 ();
 FILLCELL_X4 FILLER_36_67 ();
 FILLCELL_X1 FILLER_36_71 ();
 FILLCELL_X4 FILLER_36_77 ();
 FILLCELL_X1 FILLER_36_81 ();
 FILLCELL_X1 FILLER_36_98 ();
 FILLCELL_X4 FILLER_36_103 ();
 FILLCELL_X2 FILLER_36_107 ();
 FILLCELL_X1 FILLER_36_109 ();
 FILLCELL_X8 FILLER_36_113 ();
 FILLCELL_X2 FILLER_36_121 ();
 FILLCELL_X1 FILLER_36_123 ();
 FILLCELL_X1 FILLER_36_148 ();
 FILLCELL_X8 FILLER_36_166 ();
 FILLCELL_X4 FILLER_36_178 ();
 FILLCELL_X8 FILLER_36_185 ();
 FILLCELL_X2 FILLER_36_193 ();
 FILLCELL_X4 FILLER_36_202 ();
 FILLCELL_X2 FILLER_36_206 ();
 FILLCELL_X1 FILLER_36_208 ();
 FILLCELL_X1 FILLER_36_212 ();
 FILLCELL_X4 FILLER_36_230 ();
 FILLCELL_X2 FILLER_36_234 ();
 FILLCELL_X8 FILLER_36_267 ();
 FILLCELL_X4 FILLER_36_275 ();
 FILLCELL_X1 FILLER_36_286 ();
 FILLCELL_X2 FILLER_36_294 ();
 FILLCELL_X1 FILLER_36_296 ();
 FILLCELL_X4 FILLER_36_316 ();
 FILLCELL_X2 FILLER_36_320 ();
 FILLCELL_X1 FILLER_36_322 ();
 FILLCELL_X2 FILLER_36_327 ();
 FILLCELL_X4 FILLER_36_333 ();
 FILLCELL_X2 FILLER_36_337 ();
 FILLCELL_X16 FILLER_36_346 ();
 FILLCELL_X4 FILLER_36_368 ();
 FILLCELL_X1 FILLER_36_379 ();
 FILLCELL_X8 FILLER_36_387 ();
 FILLCELL_X4 FILLER_36_395 ();
 FILLCELL_X1 FILLER_36_399 ();
 FILLCELL_X1 FILLER_36_441 ();
 FILLCELL_X2 FILLER_36_447 ();
 FILLCELL_X1 FILLER_36_449 ();
 FILLCELL_X8 FILLER_36_460 ();
 FILLCELL_X4 FILLER_36_468 ();
 FILLCELL_X2 FILLER_36_472 ();
 FILLCELL_X1 FILLER_36_491 ();
 FILLCELL_X1 FILLER_36_509 ();
 FILLCELL_X4 FILLER_36_514 ();
 FILLCELL_X2 FILLER_36_518 ();
 FILLCELL_X4 FILLER_36_544 ();
 FILLCELL_X2 FILLER_36_548 ();
 FILLCELL_X2 FILLER_36_557 ();
 FILLCELL_X1 FILLER_36_559 ();
 FILLCELL_X8 FILLER_36_565 ();
 FILLCELL_X4 FILLER_36_573 ();
 FILLCELL_X2 FILLER_36_577 ();
 FILLCELL_X2 FILLER_36_584 ();
 FILLCELL_X1 FILLER_36_586 ();
 FILLCELL_X16 FILLER_36_595 ();
 FILLCELL_X4 FILLER_36_611 ();
 FILLCELL_X2 FILLER_36_615 ();
 FILLCELL_X1 FILLER_36_617 ();
 FILLCELL_X1 FILLER_36_630 ();
 FILLCELL_X2 FILLER_36_632 ();
 FILLCELL_X1 FILLER_36_634 ();
 FILLCELL_X1 FILLER_36_637 ();
 FILLCELL_X4 FILLER_36_693 ();
 FILLCELL_X1 FILLER_36_714 ();
 FILLCELL_X1 FILLER_36_722 ();
 FILLCELL_X8 FILLER_36_726 ();
 FILLCELL_X4 FILLER_36_734 ();
 FILLCELL_X2 FILLER_36_738 ();
 FILLCELL_X1 FILLER_36_740 ();
 FILLCELL_X2 FILLER_36_744 ();
 FILLCELL_X1 FILLER_36_746 ();
 FILLCELL_X4 FILLER_36_764 ();
 FILLCELL_X1 FILLER_36_768 ();
 FILLCELL_X4 FILLER_36_772 ();
 FILLCELL_X1 FILLER_36_776 ();
 FILLCELL_X8 FILLER_36_785 ();
 FILLCELL_X4 FILLER_36_807 ();
 FILLCELL_X2 FILLER_36_811 ();
 FILLCELL_X1 FILLER_36_813 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X16 FILLER_37_33 ();
 FILLCELL_X4 FILLER_37_49 ();
 FILLCELL_X2 FILLER_37_53 ();
 FILLCELL_X4 FILLER_37_60 ();
 FILLCELL_X8 FILLER_37_69 ();
 FILLCELL_X1 FILLER_37_77 ();
 FILLCELL_X1 FILLER_37_82 ();
 FILLCELL_X2 FILLER_37_100 ();
 FILLCELL_X2 FILLER_37_109 ();
 FILLCELL_X2 FILLER_37_118 ();
 FILLCELL_X1 FILLER_37_120 ();
 FILLCELL_X1 FILLER_37_142 ();
 FILLCELL_X2 FILLER_37_148 ();
 FILLCELL_X1 FILLER_37_150 ();
 FILLCELL_X2 FILLER_37_165 ();
 FILLCELL_X1 FILLER_37_167 ();
 FILLCELL_X2 FILLER_37_185 ();
 FILLCELL_X1 FILLER_37_187 ();
 FILLCELL_X4 FILLER_37_205 ();
 FILLCELL_X1 FILLER_37_209 ();
 FILLCELL_X4 FILLER_37_224 ();
 FILLCELL_X16 FILLER_37_235 ();
 FILLCELL_X4 FILLER_37_251 ();
 FILLCELL_X2 FILLER_37_262 ();
 FILLCELL_X8 FILLER_37_285 ();
 FILLCELL_X1 FILLER_37_293 ();
 FILLCELL_X4 FILLER_37_312 ();
 FILLCELL_X1 FILLER_37_316 ();
 FILLCELL_X4 FILLER_37_334 ();
 FILLCELL_X1 FILLER_37_338 ();
 FILLCELL_X2 FILLER_37_346 ();
 FILLCELL_X1 FILLER_37_348 ();
 FILLCELL_X8 FILLER_37_356 ();
 FILLCELL_X1 FILLER_37_364 ();
 FILLCELL_X1 FILLER_37_369 ();
 FILLCELL_X1 FILLER_37_373 ();
 FILLCELL_X2 FILLER_37_377 ();
 FILLCELL_X2 FILLER_37_386 ();
 FILLCELL_X2 FILLER_37_395 ();
 FILLCELL_X16 FILLER_37_404 ();
 FILLCELL_X2 FILLER_37_420 ();
 FILLCELL_X1 FILLER_37_422 ();
 FILLCELL_X8 FILLER_37_432 ();
 FILLCELL_X1 FILLER_37_440 ();
 FILLCELL_X1 FILLER_37_448 ();
 FILLCELL_X8 FILLER_37_473 ();
 FILLCELL_X2 FILLER_37_481 ();
 FILLCELL_X1 FILLER_37_483 ();
 FILLCELL_X2 FILLER_37_488 ();
 FILLCELL_X1 FILLER_37_490 ();
 FILLCELL_X32 FILLER_37_494 ();
 FILLCELL_X8 FILLER_37_526 ();
 FILLCELL_X4 FILLER_37_534 ();
 FILLCELL_X2 FILLER_37_538 ();
 FILLCELL_X1 FILLER_37_540 ();
 FILLCELL_X2 FILLER_37_546 ();
 FILLCELL_X1 FILLER_37_548 ();
 FILLCELL_X2 FILLER_37_568 ();
 FILLCELL_X1 FILLER_37_570 ();
 FILLCELL_X2 FILLER_37_575 ();
 FILLCELL_X1 FILLER_37_577 ();
 FILLCELL_X4 FILLER_37_582 ();
 FILLCELL_X2 FILLER_37_586 ();
 FILLCELL_X8 FILLER_37_605 ();
 FILLCELL_X1 FILLER_37_619 ();
 FILLCELL_X4 FILLER_37_637 ();
 FILLCELL_X4 FILLER_37_661 ();
 FILLCELL_X2 FILLER_37_665 ();
 FILLCELL_X1 FILLER_37_667 ();
 FILLCELL_X4 FILLER_37_702 ();
 FILLCELL_X1 FILLER_37_706 ();
 FILLCELL_X2 FILLER_37_711 ();
 FILLCELL_X1 FILLER_37_713 ();
 FILLCELL_X2 FILLER_37_721 ();
 FILLCELL_X4 FILLER_37_726 ();
 FILLCELL_X4 FILLER_37_739 ();
 FILLCELL_X2 FILLER_37_753 ();
 FILLCELL_X1 FILLER_37_755 ();
 FILLCELL_X8 FILLER_37_760 ();
 FILLCELL_X8 FILLER_37_772 ();
 FILLCELL_X4 FILLER_37_787 ();
 FILLCELL_X16 FILLER_38_1 ();
 FILLCELL_X8 FILLER_38_17 ();
 FILLCELL_X1 FILLER_38_25 ();
 FILLCELL_X8 FILLER_38_48 ();
 FILLCELL_X2 FILLER_38_56 ();
 FILLCELL_X1 FILLER_38_58 ();
 FILLCELL_X8 FILLER_38_93 ();
 FILLCELL_X8 FILLER_38_122 ();
 FILLCELL_X4 FILLER_38_130 ();
 FILLCELL_X2 FILLER_38_134 ();
 FILLCELL_X1 FILLER_38_136 ();
 FILLCELL_X4 FILLER_38_141 ();
 FILLCELL_X2 FILLER_38_145 ();
 FILLCELL_X1 FILLER_38_147 ();
 FILLCELL_X8 FILLER_38_155 ();
 FILLCELL_X4 FILLER_38_170 ();
 FILLCELL_X8 FILLER_38_177 ();
 FILLCELL_X16 FILLER_38_192 ();
 FILLCELL_X1 FILLER_38_208 ();
 FILLCELL_X8 FILLER_38_230 ();
 FILLCELL_X4 FILLER_38_238 ();
 FILLCELL_X4 FILLER_38_283 ();
 FILLCELL_X1 FILLER_38_287 ();
 FILLCELL_X2 FILLER_38_305 ();
 FILLCELL_X16 FILLER_38_310 ();
 FILLCELL_X8 FILLER_38_326 ();
 FILLCELL_X1 FILLER_38_334 ();
 FILLCELL_X4 FILLER_38_356 ();
 FILLCELL_X2 FILLER_38_377 ();
 FILLCELL_X16 FILLER_38_393 ();
 FILLCELL_X2 FILLER_38_409 ();
 FILLCELL_X1 FILLER_38_411 ();
 FILLCELL_X1 FILLER_38_415 ();
 FILLCELL_X8 FILLER_38_426 ();
 FILLCELL_X4 FILLER_38_434 ();
 FILLCELL_X2 FILLER_38_442 ();
 FILLCELL_X4 FILLER_38_447 ();
 FILLCELL_X1 FILLER_38_470 ();
 FILLCELL_X2 FILLER_38_474 ();
 FILLCELL_X2 FILLER_38_483 ();
 FILLCELL_X2 FILLER_38_499 ();
 FILLCELL_X8 FILLER_38_515 ();
 FILLCELL_X2 FILLER_38_523 ();
 FILLCELL_X1 FILLER_38_525 ();
 FILLCELL_X4 FILLER_38_542 ();
 FILLCELL_X1 FILLER_38_546 ();
 FILLCELL_X8 FILLER_38_553 ();
 FILLCELL_X4 FILLER_38_561 ();
 FILLCELL_X2 FILLER_38_565 ();
 FILLCELL_X1 FILLER_38_567 ();
 FILLCELL_X1 FILLER_38_587 ();
 FILLCELL_X2 FILLER_38_595 ();
 FILLCELL_X1 FILLER_38_597 ();
 FILLCELL_X4 FILLER_38_605 ();
 FILLCELL_X2 FILLER_38_609 ();
 FILLCELL_X1 FILLER_38_611 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X8 FILLER_38_632 ();
 FILLCELL_X1 FILLER_38_640 ();
 FILLCELL_X4 FILLER_38_650 ();
 FILLCELL_X2 FILLER_38_654 ();
 FILLCELL_X1 FILLER_38_656 ();
 FILLCELL_X2 FILLER_38_660 ();
 FILLCELL_X1 FILLER_38_676 ();
 FILLCELL_X16 FILLER_38_682 ();
 FILLCELL_X4 FILLER_38_698 ();
 FILLCELL_X1 FILLER_38_702 ();
 FILLCELL_X8 FILLER_38_707 ();
 FILLCELL_X4 FILLER_38_715 ();
 FILLCELL_X1 FILLER_38_719 ();
 FILLCELL_X1 FILLER_38_729 ();
 FILLCELL_X1 FILLER_38_734 ();
 FILLCELL_X1 FILLER_38_738 ();
 FILLCELL_X4 FILLER_38_751 ();
 FILLCELL_X1 FILLER_38_755 ();
 FILLCELL_X4 FILLER_38_761 ();
 FILLCELL_X2 FILLER_38_765 ();
 FILLCELL_X1 FILLER_38_767 ();
 FILLCELL_X4 FILLER_38_771 ();
 FILLCELL_X8 FILLER_38_799 ();
 FILLCELL_X4 FILLER_38_807 ();
 FILLCELL_X2 FILLER_38_811 ();
 FILLCELL_X1 FILLER_38_813 ();
 FILLCELL_X16 FILLER_39_1 ();
 FILLCELL_X8 FILLER_39_17 ();
 FILLCELL_X4 FILLER_39_25 ();
 FILLCELL_X2 FILLER_39_29 ();
 FILLCELL_X16 FILLER_39_48 ();
 FILLCELL_X1 FILLER_39_64 ();
 FILLCELL_X8 FILLER_39_76 ();
 FILLCELL_X2 FILLER_39_84 ();
 FILLCELL_X1 FILLER_39_86 ();
 FILLCELL_X2 FILLER_39_91 ();
 FILLCELL_X1 FILLER_39_93 ();
 FILLCELL_X8 FILLER_39_100 ();
 FILLCELL_X2 FILLER_39_108 ();
 FILLCELL_X16 FILLER_39_117 ();
 FILLCELL_X1 FILLER_39_133 ();
 FILLCELL_X1 FILLER_39_141 ();
 FILLCELL_X2 FILLER_39_145 ();
 FILLCELL_X1 FILLER_39_147 ();
 FILLCELL_X1 FILLER_39_155 ();
 FILLCELL_X4 FILLER_39_163 ();
 FILLCELL_X2 FILLER_39_167 ();
 FILLCELL_X1 FILLER_39_169 ();
 FILLCELL_X1 FILLER_39_177 ();
 FILLCELL_X2 FILLER_39_181 ();
 FILLCELL_X1 FILLER_39_190 ();
 FILLCELL_X2 FILLER_39_198 ();
 FILLCELL_X8 FILLER_39_209 ();
 FILLCELL_X4 FILLER_39_217 ();
 FILLCELL_X16 FILLER_39_239 ();
 FILLCELL_X4 FILLER_39_255 ();
 FILLCELL_X2 FILLER_39_259 ();
 FILLCELL_X2 FILLER_39_266 ();
 FILLCELL_X4 FILLER_39_275 ();
 FILLCELL_X1 FILLER_39_303 ();
 FILLCELL_X1 FILLER_39_308 ();
 FILLCELL_X1 FILLER_39_312 ();
 FILLCELL_X8 FILLER_39_317 ();
 FILLCELL_X1 FILLER_39_325 ();
 FILLCELL_X1 FILLER_39_346 ();
 FILLCELL_X16 FILLER_39_354 ();
 FILLCELL_X4 FILLER_39_377 ();
 FILLCELL_X2 FILLER_39_381 ();
 FILLCELL_X1 FILLER_39_383 ();
 FILLCELL_X2 FILLER_39_391 ();
 FILLCELL_X4 FILLER_39_400 ();
 FILLCELL_X1 FILLER_39_404 ();
 FILLCELL_X2 FILLER_39_492 ();
 FILLCELL_X2 FILLER_39_511 ();
 FILLCELL_X1 FILLER_39_532 ();
 FILLCELL_X2 FILLER_39_535 ();
 FILLCELL_X2 FILLER_39_541 ();
 FILLCELL_X1 FILLER_39_543 ();
 FILLCELL_X4 FILLER_39_548 ();
 FILLCELL_X2 FILLER_39_552 ();
 FILLCELL_X2 FILLER_39_564 ();
 FILLCELL_X2 FILLER_39_570 ();
 FILLCELL_X1 FILLER_39_572 ();
 FILLCELL_X1 FILLER_39_580 ();
 FILLCELL_X1 FILLER_39_588 ();
 FILLCELL_X1 FILLER_39_591 ();
 FILLCELL_X1 FILLER_39_603 ();
 FILLCELL_X8 FILLER_39_606 ();
 FILLCELL_X2 FILLER_39_614 ();
 FILLCELL_X1 FILLER_39_616 ();
 FILLCELL_X1 FILLER_39_623 ();
 FILLCELL_X2 FILLER_39_629 ();
 FILLCELL_X1 FILLER_39_631 ();
 FILLCELL_X1 FILLER_39_658 ();
 FILLCELL_X2 FILLER_39_664 ();
 FILLCELL_X1 FILLER_39_666 ();
 FILLCELL_X8 FILLER_39_679 ();
 FILLCELL_X2 FILLER_39_687 ();
 FILLCELL_X8 FILLER_39_694 ();
 FILLCELL_X1 FILLER_39_702 ();
 FILLCELL_X16 FILLER_39_710 ();
 FILLCELL_X1 FILLER_39_726 ();
 FILLCELL_X1 FILLER_39_735 ();
 FILLCELL_X4 FILLER_39_743 ();
 FILLCELL_X1 FILLER_39_747 ();
 FILLCELL_X1 FILLER_39_755 ();
 FILLCELL_X16 FILLER_39_773 ();
 FILLCELL_X4 FILLER_39_789 ();
 FILLCELL_X2 FILLER_39_793 ();
 FILLCELL_X8 FILLER_39_803 ();
 FILLCELL_X8 FILLER_40_1 ();
 FILLCELL_X8 FILLER_40_13 ();
 FILLCELL_X4 FILLER_40_21 ();
 FILLCELL_X2 FILLER_40_25 ();
 FILLCELL_X1 FILLER_40_27 ();
 FILLCELL_X4 FILLER_40_39 ();
 FILLCELL_X2 FILLER_40_46 ();
 FILLCELL_X2 FILLER_40_51 ();
 FILLCELL_X1 FILLER_40_53 ();
 FILLCELL_X1 FILLER_40_71 ();
 FILLCELL_X2 FILLER_40_86 ();
 FILLCELL_X2 FILLER_40_105 ();
 FILLCELL_X1 FILLER_40_107 ();
 FILLCELL_X2 FILLER_40_112 ();
 FILLCELL_X1 FILLER_40_114 ();
 FILLCELL_X8 FILLER_40_118 ();
 FILLCELL_X4 FILLER_40_126 ();
 FILLCELL_X1 FILLER_40_130 ();
 FILLCELL_X8 FILLER_40_153 ();
 FILLCELL_X4 FILLER_40_161 ();
 FILLCELL_X2 FILLER_40_165 ();
 FILLCELL_X1 FILLER_40_167 ();
 FILLCELL_X1 FILLER_40_185 ();
 FILLCELL_X8 FILLER_40_200 ();
 FILLCELL_X4 FILLER_40_208 ();
 FILLCELL_X1 FILLER_40_212 ();
 FILLCELL_X16 FILLER_40_225 ();
 FILLCELL_X4 FILLER_40_241 ();
 FILLCELL_X2 FILLER_40_245 ();
 FILLCELL_X1 FILLER_40_247 ();
 FILLCELL_X2 FILLER_40_252 ();
 FILLCELL_X1 FILLER_40_254 ();
 FILLCELL_X8 FILLER_40_258 ();
 FILLCELL_X1 FILLER_40_266 ();
 FILLCELL_X8 FILLER_40_272 ();
 FILLCELL_X4 FILLER_40_280 ();
 FILLCELL_X1 FILLER_40_284 ();
 FILLCELL_X4 FILLER_40_292 ();
 FILLCELL_X1 FILLER_40_296 ();
 FILLCELL_X8 FILLER_40_300 ();
 FILLCELL_X16 FILLER_40_350 ();
 FILLCELL_X8 FILLER_40_386 ();
 FILLCELL_X8 FILLER_40_401 ();
 FILLCELL_X2 FILLER_40_409 ();
 FILLCELL_X1 FILLER_40_411 ();
 FILLCELL_X8 FILLER_40_429 ();
 FILLCELL_X1 FILLER_40_437 ();
 FILLCELL_X4 FILLER_40_441 ();
 FILLCELL_X1 FILLER_40_445 ();
 FILLCELL_X32 FILLER_40_455 ();
 FILLCELL_X8 FILLER_40_487 ();
 FILLCELL_X2 FILLER_40_495 ();
 FILLCELL_X8 FILLER_40_504 ();
 FILLCELL_X4 FILLER_40_512 ();
 FILLCELL_X2 FILLER_40_516 ();
 FILLCELL_X1 FILLER_40_521 ();
 FILLCELL_X4 FILLER_40_561 ();
 FILLCELL_X2 FILLER_40_565 ();
 FILLCELL_X8 FILLER_40_569 ();
 FILLCELL_X1 FILLER_40_577 ();
 FILLCELL_X2 FILLER_40_593 ();
 FILLCELL_X1 FILLER_40_609 ();
 FILLCELL_X2 FILLER_40_615 ();
 FILLCELL_X1 FILLER_40_617 ();
 FILLCELL_X8 FILLER_40_623 ();
 FILLCELL_X2 FILLER_40_632 ();
 FILLCELL_X4 FILLER_40_636 ();
 FILLCELL_X1 FILLER_40_640 ();
 FILLCELL_X8 FILLER_40_643 ();
 FILLCELL_X2 FILLER_40_651 ();
 FILLCELL_X2 FILLER_40_660 ();
 FILLCELL_X8 FILLER_40_667 ();
 FILLCELL_X8 FILLER_40_682 ();
 FILLCELL_X4 FILLER_40_690 ();
 FILLCELL_X1 FILLER_40_694 ();
 FILLCELL_X2 FILLER_40_719 ();
 FILLCELL_X1 FILLER_40_721 ();
 FILLCELL_X8 FILLER_40_727 ();
 FILLCELL_X2 FILLER_40_745 ();
 FILLCELL_X1 FILLER_40_747 ();
 FILLCELL_X4 FILLER_40_755 ();
 FILLCELL_X1 FILLER_40_759 ();
 FILLCELL_X32 FILLER_40_765 ();
 FILLCELL_X1 FILLER_40_810 ();
 FILLCELL_X16 FILLER_41_1 ();
 FILLCELL_X2 FILLER_41_17 ();
 FILLCELL_X4 FILLER_41_39 ();
 FILLCELL_X1 FILLER_41_85 ();
 FILLCELL_X4 FILLER_41_93 ();
 FILLCELL_X2 FILLER_41_97 ();
 FILLCELL_X1 FILLER_41_99 ();
 FILLCELL_X1 FILLER_41_117 ();
 FILLCELL_X32 FILLER_41_125 ();
 FILLCELL_X8 FILLER_41_164 ();
 FILLCELL_X2 FILLER_41_172 ();
 FILLCELL_X4 FILLER_41_181 ();
 FILLCELL_X2 FILLER_41_185 ();
 FILLCELL_X1 FILLER_41_187 ();
 FILLCELL_X8 FILLER_41_195 ();
 FILLCELL_X8 FILLER_41_210 ();
 FILLCELL_X1 FILLER_41_238 ();
 FILLCELL_X1 FILLER_41_256 ();
 FILLCELL_X32 FILLER_41_274 ();
 FILLCELL_X2 FILLER_41_306 ();
 FILLCELL_X4 FILLER_41_316 ();
 FILLCELL_X1 FILLER_41_320 ();
 FILLCELL_X4 FILLER_41_328 ();
 FILLCELL_X8 FILLER_41_337 ();
 FILLCELL_X4 FILLER_41_345 ();
 FILLCELL_X2 FILLER_41_349 ();
 FILLCELL_X4 FILLER_41_372 ();
 FILLCELL_X2 FILLER_41_376 ();
 FILLCELL_X16 FILLER_41_383 ();
 FILLCELL_X8 FILLER_41_399 ();
 FILLCELL_X4 FILLER_41_407 ();
 FILLCELL_X1 FILLER_41_411 ();
 FILLCELL_X32 FILLER_41_426 ();
 FILLCELL_X32 FILLER_41_458 ();
 FILLCELL_X16 FILLER_41_490 ();
 FILLCELL_X8 FILLER_41_506 ();
 FILLCELL_X1 FILLER_41_514 ();
 FILLCELL_X8 FILLER_41_520 ();
 FILLCELL_X4 FILLER_41_528 ();
 FILLCELL_X2 FILLER_41_532 ();
 FILLCELL_X2 FILLER_41_539 ();
 FILLCELL_X2 FILLER_41_587 ();
 FILLCELL_X1 FILLER_41_612 ();
 FILLCELL_X1 FILLER_41_618 ();
 FILLCELL_X4 FILLER_41_621 ();
 FILLCELL_X1 FILLER_41_625 ();
 FILLCELL_X4 FILLER_41_645 ();
 FILLCELL_X2 FILLER_41_649 ();
 FILLCELL_X8 FILLER_41_668 ();
 FILLCELL_X1 FILLER_41_676 ();
 FILLCELL_X2 FILLER_41_684 ();
 FILLCELL_X1 FILLER_41_686 ();
 FILLCELL_X2 FILLER_41_733 ();
 FILLCELL_X1 FILLER_41_735 ();
 FILLCELL_X1 FILLER_41_743 ();
 FILLCELL_X1 FILLER_41_747 ();
 FILLCELL_X2 FILLER_41_762 ();
 FILLCELL_X8 FILLER_41_768 ();
 FILLCELL_X1 FILLER_41_793 ();
 FILLCELL_X16 FILLER_42_1 ();
 FILLCELL_X4 FILLER_42_17 ();
 FILLCELL_X1 FILLER_42_21 ();
 FILLCELL_X4 FILLER_42_32 ();
 FILLCELL_X2 FILLER_42_36 ();
 FILLCELL_X8 FILLER_42_43 ();
 FILLCELL_X4 FILLER_42_51 ();
 FILLCELL_X16 FILLER_42_69 ();
 FILLCELL_X4 FILLER_42_85 ();
 FILLCELL_X1 FILLER_42_89 ();
 FILLCELL_X8 FILLER_42_95 ();
 FILLCELL_X4 FILLER_42_103 ();
 FILLCELL_X2 FILLER_42_107 ();
 FILLCELL_X1 FILLER_42_109 ();
 FILLCELL_X1 FILLER_42_113 ();
 FILLCELL_X2 FILLER_42_154 ();
 FILLCELL_X1 FILLER_42_156 ();
 FILLCELL_X2 FILLER_42_164 ();
 FILLCELL_X8 FILLER_42_175 ();
 FILLCELL_X1 FILLER_42_183 ();
 FILLCELL_X2 FILLER_42_191 ();
 FILLCELL_X4 FILLER_42_196 ();
 FILLCELL_X2 FILLER_42_200 ();
 FILLCELL_X1 FILLER_42_202 ();
 FILLCELL_X1 FILLER_42_216 ();
 FILLCELL_X2 FILLER_42_248 ();
 FILLCELL_X4 FILLER_42_253 ();
 FILLCELL_X2 FILLER_42_257 ();
 FILLCELL_X4 FILLER_42_266 ();
 FILLCELL_X1 FILLER_42_270 ();
 FILLCELL_X8 FILLER_42_288 ();
 FILLCELL_X4 FILLER_42_296 ();
 FILLCELL_X2 FILLER_42_300 ();
 FILLCELL_X1 FILLER_42_302 ();
 FILLCELL_X8 FILLER_42_320 ();
 FILLCELL_X1 FILLER_42_328 ();
 FILLCELL_X8 FILLER_42_339 ();
 FILLCELL_X2 FILLER_42_347 ();
 FILLCELL_X1 FILLER_42_358 ();
 FILLCELL_X1 FILLER_42_366 ();
 FILLCELL_X1 FILLER_42_381 ();
 FILLCELL_X4 FILLER_42_389 ();
 FILLCELL_X1 FILLER_42_393 ();
 FILLCELL_X4 FILLER_42_401 ();
 FILLCELL_X2 FILLER_42_405 ();
 FILLCELL_X4 FILLER_42_418 ();
 FILLCELL_X1 FILLER_42_422 ();
 FILLCELL_X4 FILLER_42_426 ();
 FILLCELL_X2 FILLER_42_430 ();
 FILLCELL_X1 FILLER_42_432 ();
 FILLCELL_X1 FILLER_42_437 ();
 FILLCELL_X1 FILLER_42_444 ();
 FILLCELL_X2 FILLER_42_462 ();
 FILLCELL_X2 FILLER_42_467 ();
 FILLCELL_X1 FILLER_42_469 ();
 FILLCELL_X1 FILLER_42_482 ();
 FILLCELL_X2 FILLER_42_500 ();
 FILLCELL_X1 FILLER_42_502 ();
 FILLCELL_X2 FILLER_42_506 ();
 FILLCELL_X4 FILLER_42_525 ();
 FILLCELL_X2 FILLER_42_529 ();
 FILLCELL_X1 FILLER_42_531 ();
 FILLCELL_X2 FILLER_42_539 ();
 FILLCELL_X1 FILLER_42_541 ();
 FILLCELL_X4 FILLER_42_550 ();
 FILLCELL_X2 FILLER_42_554 ();
 FILLCELL_X2 FILLER_42_563 ();
 FILLCELL_X2 FILLER_42_594 ();
 FILLCELL_X1 FILLER_42_596 ();
 FILLCELL_X4 FILLER_42_605 ();
 FILLCELL_X8 FILLER_42_632 ();
 FILLCELL_X4 FILLER_42_640 ();
 FILLCELL_X2 FILLER_42_652 ();
 FILLCELL_X1 FILLER_42_662 ();
 FILLCELL_X4 FILLER_42_671 ();
 FILLCELL_X2 FILLER_42_675 ();
 FILLCELL_X1 FILLER_42_677 ();
 FILLCELL_X8 FILLER_42_685 ();
 FILLCELL_X2 FILLER_42_693 ();
 FILLCELL_X1 FILLER_42_707 ();
 FILLCELL_X2 FILLER_42_712 ();
 FILLCELL_X2 FILLER_42_718 ();
 FILLCELL_X2 FILLER_42_729 ();
 FILLCELL_X1 FILLER_42_731 ();
 FILLCELL_X1 FILLER_42_736 ();
 FILLCELL_X4 FILLER_42_754 ();
 FILLCELL_X2 FILLER_42_805 ();
 FILLCELL_X1 FILLER_42_807 ();
 FILLCELL_X2 FILLER_42_811 ();
 FILLCELL_X1 FILLER_42_813 ();
 FILLCELL_X8 FILLER_43_1 ();
 FILLCELL_X4 FILLER_43_9 ();
 FILLCELL_X1 FILLER_43_13 ();
 FILLCELL_X16 FILLER_43_18 ();
 FILLCELL_X8 FILLER_43_34 ();
 FILLCELL_X4 FILLER_43_42 ();
 FILLCELL_X1 FILLER_43_71 ();
 FILLCELL_X4 FILLER_43_86 ();
 FILLCELL_X4 FILLER_43_107 ();
 FILLCELL_X2 FILLER_43_111 ();
 FILLCELL_X16 FILLER_43_123 ();
 FILLCELL_X4 FILLER_43_139 ();
 FILLCELL_X1 FILLER_43_150 ();
 FILLCELL_X8 FILLER_43_161 ();
 FILLCELL_X1 FILLER_43_169 ();
 FILLCELL_X4 FILLER_43_194 ();
 FILLCELL_X1 FILLER_43_198 ();
 FILLCELL_X8 FILLER_43_223 ();
 FILLCELL_X4 FILLER_43_231 ();
 FILLCELL_X1 FILLER_43_235 ();
 FILLCELL_X8 FILLER_43_239 ();
 FILLCELL_X1 FILLER_43_247 ();
 FILLCELL_X4 FILLER_43_262 ();
 FILLCELL_X1 FILLER_43_266 ();
 FILLCELL_X8 FILLER_43_295 ();
 FILLCELL_X1 FILLER_43_303 ();
 FILLCELL_X16 FILLER_43_311 ();
 FILLCELL_X1 FILLER_43_327 ();
 FILLCELL_X2 FILLER_43_345 ();
 FILLCELL_X2 FILLER_43_351 ();
 FILLCELL_X1 FILLER_43_353 ();
 FILLCELL_X2 FILLER_43_357 ();
 FILLCELL_X1 FILLER_43_373 ();
 FILLCELL_X16 FILLER_43_381 ();
 FILLCELL_X4 FILLER_43_397 ();
 FILLCELL_X1 FILLER_43_427 ();
 FILLCELL_X1 FILLER_43_454 ();
 FILLCELL_X4 FILLER_43_459 ();
 FILLCELL_X2 FILLER_43_463 ();
 FILLCELL_X1 FILLER_43_465 ();
 FILLCELL_X2 FILLER_43_471 ();
 FILLCELL_X1 FILLER_43_473 ();
 FILLCELL_X2 FILLER_43_481 ();
 FILLCELL_X2 FILLER_43_490 ();
 FILLCELL_X1 FILLER_43_495 ();
 FILLCELL_X2 FILLER_43_501 ();
 FILLCELL_X1 FILLER_43_503 ();
 FILLCELL_X1 FILLER_43_532 ();
 FILLCELL_X1 FILLER_43_535 ();
 FILLCELL_X1 FILLER_43_540 ();
 FILLCELL_X2 FILLER_43_564 ();
 FILLCELL_X1 FILLER_43_566 ();
 FILLCELL_X1 FILLER_43_571 ();
 FILLCELL_X4 FILLER_43_574 ();
 FILLCELL_X2 FILLER_43_578 ();
 FILLCELL_X16 FILLER_43_584 ();
 FILLCELL_X8 FILLER_43_600 ();
 FILLCELL_X16 FILLER_43_616 ();
 FILLCELL_X4 FILLER_43_632 ();
 FILLCELL_X2 FILLER_43_636 ();
 FILLCELL_X2 FILLER_43_655 ();
 FILLCELL_X8 FILLER_43_677 ();
 FILLCELL_X4 FILLER_43_685 ();
 FILLCELL_X4 FILLER_43_693 ();
 FILLCELL_X1 FILLER_43_697 ();
 FILLCELL_X1 FILLER_43_702 ();
 FILLCELL_X1 FILLER_43_711 ();
 FILLCELL_X2 FILLER_43_733 ();
 FILLCELL_X8 FILLER_43_742 ();
 FILLCELL_X1 FILLER_43_750 ();
 FILLCELL_X8 FILLER_43_754 ();
 FILLCELL_X1 FILLER_43_778 ();
 FILLCELL_X8 FILLER_44_1 ();
 FILLCELL_X4 FILLER_44_9 ();
 FILLCELL_X2 FILLER_44_13 ();
 FILLCELL_X1 FILLER_44_15 ();
 FILLCELL_X2 FILLER_44_40 ();
 FILLCELL_X1 FILLER_44_42 ();
 FILLCELL_X4 FILLER_44_48 ();
 FILLCELL_X2 FILLER_44_52 ();
 FILLCELL_X4 FILLER_44_58 ();
 FILLCELL_X1 FILLER_44_69 ();
 FILLCELL_X1 FILLER_44_84 ();
 FILLCELL_X4 FILLER_44_92 ();
 FILLCELL_X2 FILLER_44_96 ();
 FILLCELL_X8 FILLER_44_127 ();
 FILLCELL_X4 FILLER_44_135 ();
 FILLCELL_X4 FILLER_44_143 ();
 FILLCELL_X16 FILLER_44_150 ();
 FILLCELL_X4 FILLER_44_166 ();
 FILLCELL_X1 FILLER_44_170 ();
 FILLCELL_X16 FILLER_44_178 ();
 FILLCELL_X8 FILLER_44_197 ();
 FILLCELL_X4 FILLER_44_205 ();
 FILLCELL_X4 FILLER_44_216 ();
 FILLCELL_X2 FILLER_44_220 ();
 FILLCELL_X8 FILLER_44_225 ();
 FILLCELL_X2 FILLER_44_233 ();
 FILLCELL_X2 FILLER_44_253 ();
 FILLCELL_X1 FILLER_44_266 ();
 FILLCELL_X16 FILLER_44_270 ();
 FILLCELL_X8 FILLER_44_286 ();
 FILLCELL_X1 FILLER_44_314 ();
 FILLCELL_X1 FILLER_44_322 ();
 FILLCELL_X8 FILLER_44_330 ();
 FILLCELL_X4 FILLER_44_338 ();
 FILLCELL_X1 FILLER_44_342 ();
 FILLCELL_X4 FILLER_44_360 ();
 FILLCELL_X2 FILLER_44_364 ();
 FILLCELL_X4 FILLER_44_372 ();
 FILLCELL_X2 FILLER_44_383 ();
 FILLCELL_X1 FILLER_44_385 ();
 FILLCELL_X4 FILLER_44_393 ();
 FILLCELL_X2 FILLER_44_397 ();
 FILLCELL_X1 FILLER_44_399 ();
 FILLCELL_X1 FILLER_44_407 ();
 FILLCELL_X2 FILLER_44_421 ();
 FILLCELL_X1 FILLER_44_423 ();
 FILLCELL_X2 FILLER_44_431 ();
 FILLCELL_X1 FILLER_44_433 ();
 FILLCELL_X4 FILLER_44_437 ();
 FILLCELL_X1 FILLER_44_441 ();
 FILLCELL_X1 FILLER_44_445 ();
 FILLCELL_X8 FILLER_44_469 ();
 FILLCELL_X4 FILLER_44_477 ();
 FILLCELL_X2 FILLER_44_481 ();
 FILLCELL_X1 FILLER_44_483 ();
 FILLCELL_X1 FILLER_44_487 ();
 FILLCELL_X16 FILLER_44_502 ();
 FILLCELL_X8 FILLER_44_518 ();
 FILLCELL_X2 FILLER_44_526 ();
 FILLCELL_X1 FILLER_44_528 ();
 FILLCELL_X2 FILLER_44_536 ();
 FILLCELL_X1 FILLER_44_544 ();
 FILLCELL_X1 FILLER_44_551 ();
 FILLCELL_X1 FILLER_44_563 ();
 FILLCELL_X1 FILLER_44_566 ();
 FILLCELL_X2 FILLER_44_573 ();
 FILLCELL_X1 FILLER_44_575 ();
 FILLCELL_X1 FILLER_44_584 ();
 FILLCELL_X8 FILLER_44_596 ();
 FILLCELL_X1 FILLER_44_604 ();
 FILLCELL_X4 FILLER_44_624 ();
 FILLCELL_X2 FILLER_44_628 ();
 FILLCELL_X1 FILLER_44_630 ();
 FILLCELL_X8 FILLER_44_632 ();
 FILLCELL_X4 FILLER_44_640 ();
 FILLCELL_X2 FILLER_44_644 ();
 FILLCELL_X1 FILLER_44_646 ();
 FILLCELL_X2 FILLER_44_654 ();
 FILLCELL_X8 FILLER_44_670 ();
 FILLCELL_X4 FILLER_44_678 ();
 FILLCELL_X2 FILLER_44_682 ();
 FILLCELL_X2 FILLER_44_735 ();
 FILLCELL_X2 FILLER_44_744 ();
 FILLCELL_X2 FILLER_44_749 ();
 FILLCELL_X1 FILLER_44_755 ();
 FILLCELL_X4 FILLER_44_765 ();
 FILLCELL_X2 FILLER_44_769 ();
 FILLCELL_X1 FILLER_44_771 ();
 FILLCELL_X1 FILLER_44_789 ();
 FILLCELL_X1 FILLER_44_794 ();
 FILLCELL_X1 FILLER_44_798 ();
 FILLCELL_X2 FILLER_44_812 ();
 FILLCELL_X4 FILLER_45_1 ();
 FILLCELL_X2 FILLER_45_5 ();
 FILLCELL_X1 FILLER_45_7 ();
 FILLCELL_X16 FILLER_45_12 ();
 FILLCELL_X4 FILLER_45_28 ();
 FILLCELL_X1 FILLER_45_32 ();
 FILLCELL_X4 FILLER_45_36 ();
 FILLCELL_X2 FILLER_45_40 ();
 FILLCELL_X8 FILLER_45_67 ();
 FILLCELL_X4 FILLER_45_75 ();
 FILLCELL_X2 FILLER_45_79 ();
 FILLCELL_X1 FILLER_45_81 ();
 FILLCELL_X4 FILLER_45_87 ();
 FILLCELL_X1 FILLER_45_91 ();
 FILLCELL_X4 FILLER_45_113 ();
 FILLCELL_X1 FILLER_45_117 ();
 FILLCELL_X1 FILLER_45_132 ();
 FILLCELL_X1 FILLER_45_150 ();
 FILLCELL_X4 FILLER_45_172 ();
 FILLCELL_X2 FILLER_45_176 ();
 FILLCELL_X1 FILLER_45_195 ();
 FILLCELL_X2 FILLER_45_200 ();
 FILLCELL_X2 FILLER_45_205 ();
 FILLCELL_X2 FILLER_45_224 ();
 FILLCELL_X2 FILLER_45_253 ();
 FILLCELL_X1 FILLER_45_255 ();
 FILLCELL_X8 FILLER_45_276 ();
 FILLCELL_X2 FILLER_45_284 ();
 FILLCELL_X8 FILLER_45_303 ();
 FILLCELL_X8 FILLER_45_339 ();
 FILLCELL_X1 FILLER_45_347 ();
 FILLCELL_X32 FILLER_45_372 ();
 FILLCELL_X1 FILLER_45_404 ();
 FILLCELL_X8 FILLER_45_422 ();
 FILLCELL_X1 FILLER_45_430 ();
 FILLCELL_X2 FILLER_45_445 ();
 FILLCELL_X1 FILLER_45_447 ();
 FILLCELL_X8 FILLER_45_454 ();
 FILLCELL_X4 FILLER_45_462 ();
 FILLCELL_X2 FILLER_45_466 ();
 FILLCELL_X8 FILLER_45_475 ();
 FILLCELL_X2 FILLER_45_487 ();
 FILLCELL_X1 FILLER_45_489 ();
 FILLCELL_X8 FILLER_45_502 ();
 FILLCELL_X1 FILLER_45_514 ();
 FILLCELL_X4 FILLER_45_519 ();
 FILLCELL_X8 FILLER_45_536 ();
 FILLCELL_X4 FILLER_45_544 ();
 FILLCELL_X1 FILLER_45_554 ();
 FILLCELL_X1 FILLER_45_574 ();
 FILLCELL_X1 FILLER_45_592 ();
 FILLCELL_X16 FILLER_45_602 ();
 FILLCELL_X1 FILLER_45_618 ();
 FILLCELL_X8 FILLER_45_636 ();
 FILLCELL_X1 FILLER_45_644 ();
 FILLCELL_X32 FILLER_45_662 ();
 FILLCELL_X16 FILLER_45_694 ();
 FILLCELL_X8 FILLER_45_710 ();
 FILLCELL_X4 FILLER_45_722 ();
 FILLCELL_X2 FILLER_45_726 ();
 FILLCELL_X1 FILLER_45_728 ();
 FILLCELL_X4 FILLER_45_750 ();
 FILLCELL_X2 FILLER_45_754 ();
 FILLCELL_X4 FILLER_45_776 ();
 FILLCELL_X1 FILLER_45_780 ();
 FILLCELL_X2 FILLER_45_783 ();
 FILLCELL_X4 FILLER_45_792 ();
 FILLCELL_X2 FILLER_45_796 ();
 FILLCELL_X1 FILLER_45_798 ();
 FILLCELL_X2 FILLER_45_802 ();
 FILLCELL_X1 FILLER_45_804 ();
 FILLCELL_X2 FILLER_45_811 ();
 FILLCELL_X1 FILLER_45_813 ();
 FILLCELL_X16 FILLER_46_1 ();
 FILLCELL_X1 FILLER_46_17 ();
 FILLCELL_X4 FILLER_46_35 ();
 FILLCELL_X2 FILLER_46_39 ();
 FILLCELL_X1 FILLER_46_41 ();
 FILLCELL_X2 FILLER_46_63 ();
 FILLCELL_X1 FILLER_46_69 ();
 FILLCELL_X8 FILLER_46_77 ();
 FILLCELL_X32 FILLER_46_92 ();
 FILLCELL_X8 FILLER_46_124 ();
 FILLCELL_X4 FILLER_46_132 ();
 FILLCELL_X2 FILLER_46_136 ();
 FILLCELL_X8 FILLER_46_148 ();
 FILLCELL_X16 FILLER_46_172 ();
 FILLCELL_X4 FILLER_46_188 ();
 FILLCELL_X2 FILLER_46_192 ();
 FILLCELL_X4 FILLER_46_209 ();
 FILLCELL_X2 FILLER_46_213 ();
 FILLCELL_X1 FILLER_46_215 ();
 FILLCELL_X4 FILLER_46_223 ();
 FILLCELL_X2 FILLER_46_227 ();
 FILLCELL_X1 FILLER_46_229 ();
 FILLCELL_X4 FILLER_46_238 ();
 FILLCELL_X1 FILLER_46_242 ();
 FILLCELL_X1 FILLER_46_247 ();
 FILLCELL_X32 FILLER_46_251 ();
 FILLCELL_X8 FILLER_46_283 ();
 FILLCELL_X2 FILLER_46_291 ();
 FILLCELL_X1 FILLER_46_297 ();
 FILLCELL_X4 FILLER_46_304 ();
 FILLCELL_X1 FILLER_46_308 ();
 FILLCELL_X1 FILLER_46_316 ();
 FILLCELL_X1 FILLER_46_329 ();
 FILLCELL_X32 FILLER_46_339 ();
 FILLCELL_X2 FILLER_46_371 ();
 FILLCELL_X16 FILLER_46_378 ();
 FILLCELL_X8 FILLER_46_394 ();
 FILLCELL_X8 FILLER_46_409 ();
 FILLCELL_X2 FILLER_46_417 ();
 FILLCELL_X1 FILLER_46_419 ();
 FILLCELL_X1 FILLER_46_437 ();
 FILLCELL_X4 FILLER_46_462 ();
 FILLCELL_X2 FILLER_46_466 ();
 FILLCELL_X1 FILLER_46_475 ();
 FILLCELL_X2 FILLER_46_501 ();
 FILLCELL_X4 FILLER_46_541 ();
 FILLCELL_X2 FILLER_46_545 ();
 FILLCELL_X8 FILLER_46_557 ();
 FILLCELL_X2 FILLER_46_565 ();
 FILLCELL_X16 FILLER_46_569 ();
 FILLCELL_X4 FILLER_46_585 ();
 FILLCELL_X8 FILLER_46_617 ();
 FILLCELL_X1 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_649 ();
 FILLCELL_X4 FILLER_46_661 ();
 FILLCELL_X2 FILLER_46_665 ();
 FILLCELL_X1 FILLER_46_674 ();
 FILLCELL_X1 FILLER_46_678 ();
 FILLCELL_X8 FILLER_46_686 ();
 FILLCELL_X4 FILLER_46_694 ();
 FILLCELL_X1 FILLER_46_698 ();
 FILLCELL_X8 FILLER_46_703 ();
 FILLCELL_X4 FILLER_46_711 ();
 FILLCELL_X1 FILLER_46_715 ();
 FILLCELL_X32 FILLER_46_723 ();
 FILLCELL_X8 FILLER_46_755 ();
 FILLCELL_X4 FILLER_46_763 ();
 FILLCELL_X1 FILLER_46_767 ();
 FILLCELL_X8 FILLER_46_771 ();
 FILLCELL_X1 FILLER_46_782 ();
 FILLCELL_X1 FILLER_46_793 ();
 FILLCELL_X1 FILLER_46_810 ();
 FILLCELL_X16 FILLER_47_1 ();
 FILLCELL_X8 FILLER_47_17 ();
 FILLCELL_X1 FILLER_47_25 ();
 FILLCELL_X4 FILLER_47_36 ();
 FILLCELL_X1 FILLER_47_40 ();
 FILLCELL_X8 FILLER_47_46 ();
 FILLCELL_X4 FILLER_47_54 ();
 FILLCELL_X4 FILLER_47_63 ();
 FILLCELL_X2 FILLER_47_74 ();
 FILLCELL_X8 FILLER_47_88 ();
 FILLCELL_X1 FILLER_47_100 ();
 FILLCELL_X1 FILLER_47_110 ();
 FILLCELL_X2 FILLER_47_115 ();
 FILLCELL_X2 FILLER_47_120 ();
 FILLCELL_X2 FILLER_47_129 ();
 FILLCELL_X1 FILLER_47_131 ();
 FILLCELL_X2 FILLER_47_149 ();
 FILLCELL_X1 FILLER_47_151 ();
 FILLCELL_X1 FILLER_47_159 ();
 FILLCELL_X16 FILLER_47_167 ();
 FILLCELL_X8 FILLER_47_183 ();
 FILLCELL_X4 FILLER_47_191 ();
 FILLCELL_X2 FILLER_47_195 ();
 FILLCELL_X1 FILLER_47_197 ();
 FILLCELL_X8 FILLER_47_218 ();
 FILLCELL_X4 FILLER_47_231 ();
 FILLCELL_X2 FILLER_47_252 ();
 FILLCELL_X4 FILLER_47_271 ();
 FILLCELL_X16 FILLER_47_282 ();
 FILLCELL_X4 FILLER_47_298 ();
 FILLCELL_X1 FILLER_47_302 ();
 FILLCELL_X2 FILLER_47_310 ();
 FILLCELL_X2 FILLER_47_333 ();
 FILLCELL_X2 FILLER_47_358 ();
 FILLCELL_X1 FILLER_47_367 ();
 FILLCELL_X1 FILLER_47_372 ();
 FILLCELL_X1 FILLER_47_383 ();
 FILLCELL_X16 FILLER_47_391 ();
 FILLCELL_X2 FILLER_47_407 ();
 FILLCELL_X1 FILLER_47_409 ();
 FILLCELL_X1 FILLER_47_414 ();
 FILLCELL_X2 FILLER_47_423 ();
 FILLCELL_X4 FILLER_47_432 ();
 FILLCELL_X2 FILLER_47_436 ();
 FILLCELL_X1 FILLER_47_438 ();
 FILLCELL_X8 FILLER_47_442 ();
 FILLCELL_X1 FILLER_47_450 ();
 FILLCELL_X16 FILLER_47_468 ();
 FILLCELL_X1 FILLER_47_484 ();
 FILLCELL_X32 FILLER_47_495 ();
 FILLCELL_X16 FILLER_47_531 ();
 FILLCELL_X4 FILLER_47_547 ();
 FILLCELL_X1 FILLER_47_551 ();
 FILLCELL_X4 FILLER_47_569 ();
 FILLCELL_X2 FILLER_47_573 ();
 FILLCELL_X1 FILLER_47_575 ();
 FILLCELL_X2 FILLER_47_580 ();
 FILLCELL_X4 FILLER_47_589 ();
 FILLCELL_X4 FILLER_47_609 ();
 FILLCELL_X1 FILLER_47_613 ();
 FILLCELL_X2 FILLER_47_622 ();
 FILLCELL_X1 FILLER_47_624 ();
 FILLCELL_X1 FILLER_47_632 ();
 FILLCELL_X16 FILLER_47_638 ();
 FILLCELL_X1 FILLER_47_658 ();
 FILLCELL_X2 FILLER_47_663 ();
 FILLCELL_X2 FILLER_47_689 ();
 FILLCELL_X4 FILLER_47_712 ();
 FILLCELL_X1 FILLER_47_735 ();
 FILLCELL_X1 FILLER_47_739 ();
 FILLCELL_X4 FILLER_47_747 ();
 FILLCELL_X2 FILLER_47_751 ();
 FILLCELL_X1 FILLER_47_753 ();
 FILLCELL_X4 FILLER_47_757 ();
 FILLCELL_X1 FILLER_47_761 ();
 FILLCELL_X1 FILLER_47_766 ();
 FILLCELL_X2 FILLER_47_795 ();
 FILLCELL_X4 FILLER_48_1 ();
 FILLCELL_X1 FILLER_48_5 ();
 FILLCELL_X16 FILLER_48_10 ();
 FILLCELL_X8 FILLER_48_26 ();
 FILLCELL_X1 FILLER_48_34 ();
 FILLCELL_X4 FILLER_48_38 ();
 FILLCELL_X2 FILLER_48_42 ();
 FILLCELL_X1 FILLER_48_44 ();
 FILLCELL_X4 FILLER_48_66 ();
 FILLCELL_X2 FILLER_48_70 ();
 FILLCELL_X1 FILLER_48_86 ();
 FILLCELL_X4 FILLER_48_133 ();
 FILLCELL_X2 FILLER_48_137 ();
 FILLCELL_X1 FILLER_48_172 ();
 FILLCELL_X8 FILLER_48_194 ();
 FILLCELL_X2 FILLER_48_209 ();
 FILLCELL_X8 FILLER_48_235 ();
 FILLCELL_X4 FILLER_48_246 ();
 FILLCELL_X2 FILLER_48_250 ();
 FILLCELL_X2 FILLER_48_259 ();
 FILLCELL_X4 FILLER_48_264 ();
 FILLCELL_X2 FILLER_48_316 ();
 FILLCELL_X8 FILLER_48_323 ();
 FILLCELL_X4 FILLER_48_331 ();
 FILLCELL_X2 FILLER_48_335 ();
 FILLCELL_X1 FILLER_48_358 ();
 FILLCELL_X2 FILLER_48_383 ();
 FILLCELL_X4 FILLER_48_399 ();
 FILLCELL_X1 FILLER_48_420 ();
 FILLCELL_X1 FILLER_48_445 ();
 FILLCELL_X4 FILLER_48_453 ();
 FILLCELL_X2 FILLER_48_457 ();
 FILLCELL_X2 FILLER_48_463 ();
 FILLCELL_X4 FILLER_48_482 ();
 FILLCELL_X2 FILLER_48_490 ();
 FILLCELL_X1 FILLER_48_492 ();
 FILLCELL_X4 FILLER_48_500 ();
 FILLCELL_X1 FILLER_48_514 ();
 FILLCELL_X2 FILLER_48_519 ();
 FILLCELL_X1 FILLER_48_521 ();
 FILLCELL_X1 FILLER_48_539 ();
 FILLCELL_X1 FILLER_48_557 ();
 FILLCELL_X4 FILLER_48_560 ();
 FILLCELL_X2 FILLER_48_564 ();
 FILLCELL_X2 FILLER_48_600 ();
 FILLCELL_X4 FILLER_48_619 ();
 FILLCELL_X1 FILLER_48_628 ();
 FILLCELL_X1 FILLER_48_632 ();
 FILLCELL_X1 FILLER_48_650 ();
 FILLCELL_X1 FILLER_48_668 ();
 FILLCELL_X4 FILLER_48_673 ();
 FILLCELL_X1 FILLER_48_677 ();
 FILLCELL_X8 FILLER_48_681 ();
 FILLCELL_X4 FILLER_48_689 ();
 FILLCELL_X2 FILLER_48_693 ();
 FILLCELL_X2 FILLER_48_711 ();
 FILLCELL_X1 FILLER_48_713 ();
 FILLCELL_X1 FILLER_48_721 ();
 FILLCELL_X2 FILLER_48_731 ();
 FILLCELL_X4 FILLER_48_737 ();
 FILLCELL_X2 FILLER_48_741 ();
 FILLCELL_X2 FILLER_48_757 ();
 FILLCELL_X1 FILLER_48_759 ();
 FILLCELL_X4 FILLER_48_780 ();
 FILLCELL_X2 FILLER_48_794 ();
 FILLCELL_X1 FILLER_48_796 ();
 FILLCELL_X4 FILLER_48_800 ();
 FILLCELL_X1 FILLER_48_804 ();
 FILLCELL_X1 FILLER_48_808 ();
 FILLCELL_X2 FILLER_48_812 ();
 FILLCELL_X16 FILLER_49_1 ();
 FILLCELL_X16 FILLER_49_41 ();
 FILLCELL_X1 FILLER_49_57 ();
 FILLCELL_X2 FILLER_49_66 ();
 FILLCELL_X1 FILLER_49_68 ();
 FILLCELL_X16 FILLER_49_81 ();
 FILLCELL_X8 FILLER_49_97 ();
 FILLCELL_X4 FILLER_49_105 ();
 FILLCELL_X2 FILLER_49_109 ();
 FILLCELL_X1 FILLER_49_111 ();
 FILLCELL_X16 FILLER_49_115 ();
 FILLCELL_X2 FILLER_49_131 ();
 FILLCELL_X2 FILLER_49_137 ();
 FILLCELL_X4 FILLER_49_142 ();
 FILLCELL_X2 FILLER_49_146 ();
 FILLCELL_X8 FILLER_49_155 ();
 FILLCELL_X4 FILLER_49_163 ();
 FILLCELL_X2 FILLER_49_167 ();
 FILLCELL_X1 FILLER_49_169 ();
 FILLCELL_X4 FILLER_49_178 ();
 FILLCELL_X2 FILLER_49_182 ();
 FILLCELL_X1 FILLER_49_184 ();
 FILLCELL_X1 FILLER_49_188 ();
 FILLCELL_X1 FILLER_49_192 ();
 FILLCELL_X1 FILLER_49_196 ();
 FILLCELL_X1 FILLER_49_204 ();
 FILLCELL_X1 FILLER_49_209 ();
 FILLCELL_X1 FILLER_49_213 ();
 FILLCELL_X1 FILLER_49_217 ();
 FILLCELL_X2 FILLER_49_222 ();
 FILLCELL_X16 FILLER_49_235 ();
 FILLCELL_X2 FILLER_49_255 ();
 FILLCELL_X16 FILLER_49_260 ();
 FILLCELL_X4 FILLER_49_276 ();
 FILLCELL_X32 FILLER_49_287 ();
 FILLCELL_X4 FILLER_49_319 ();
 FILLCELL_X1 FILLER_49_323 ();
 FILLCELL_X8 FILLER_49_331 ();
 FILLCELL_X4 FILLER_49_339 ();
 FILLCELL_X2 FILLER_49_343 ();
 FILLCELL_X1 FILLER_49_345 ();
 FILLCELL_X2 FILLER_49_350 ();
 FILLCELL_X8 FILLER_49_356 ();
 FILLCELL_X4 FILLER_49_364 ();
 FILLCELL_X1 FILLER_49_368 ();
 FILLCELL_X2 FILLER_49_372 ();
 FILLCELL_X1 FILLER_49_374 ();
 FILLCELL_X16 FILLER_49_389 ();
 FILLCELL_X4 FILLER_49_405 ();
 FILLCELL_X2 FILLER_49_409 ();
 FILLCELL_X4 FILLER_49_414 ();
 FILLCELL_X4 FILLER_49_421 ();
 FILLCELL_X1 FILLER_49_425 ();
 FILLCELL_X1 FILLER_49_433 ();
 FILLCELL_X4 FILLER_49_475 ();
 FILLCELL_X2 FILLER_49_479 ();
 FILLCELL_X2 FILLER_49_505 ();
 FILLCELL_X1 FILLER_49_507 ();
 FILLCELL_X2 FILLER_49_532 ();
 FILLCELL_X4 FILLER_49_536 ();
 FILLCELL_X2 FILLER_49_540 ();
 FILLCELL_X1 FILLER_49_542 ();
 FILLCELL_X2 FILLER_49_565 ();
 FILLCELL_X4 FILLER_49_600 ();
 FILLCELL_X1 FILLER_49_604 ();
 FILLCELL_X16 FILLER_49_621 ();
 FILLCELL_X8 FILLER_49_637 ();
 FILLCELL_X4 FILLER_49_645 ();
 FILLCELL_X1 FILLER_49_649 ();
 FILLCELL_X1 FILLER_49_654 ();
 FILLCELL_X2 FILLER_49_659 ();
 FILLCELL_X1 FILLER_49_661 ();
 FILLCELL_X2 FILLER_49_689 ();
 FILLCELL_X4 FILLER_49_695 ();
 FILLCELL_X2 FILLER_49_699 ();
 FILLCELL_X2 FILLER_49_718 ();
 FILLCELL_X1 FILLER_49_720 ();
 FILLCELL_X8 FILLER_49_727 ();
 FILLCELL_X4 FILLER_49_735 ();
 FILLCELL_X2 FILLER_49_739 ();
 FILLCELL_X1 FILLER_49_741 ();
 FILLCELL_X8 FILLER_49_766 ();
 FILLCELL_X4 FILLER_49_774 ();
 FILLCELL_X4 FILLER_49_783 ();
 FILLCELL_X4 FILLER_49_790 ();
 FILLCELL_X2 FILLER_49_794 ();
 FILLCELL_X4 FILLER_49_799 ();
 FILLCELL_X2 FILLER_49_803 ();
 FILLCELL_X1 FILLER_49_805 ();
 FILLCELL_X4 FILLER_49_809 ();
 FILLCELL_X1 FILLER_49_813 ();
 FILLCELL_X4 FILLER_50_1 ();
 FILLCELL_X2 FILLER_50_5 ();
 FILLCELL_X1 FILLER_50_7 ();
 FILLCELL_X8 FILLER_50_12 ();
 FILLCELL_X2 FILLER_50_20 ();
 FILLCELL_X2 FILLER_50_25 ();
 FILLCELL_X1 FILLER_50_27 ();
 FILLCELL_X2 FILLER_50_34 ();
 FILLCELL_X2 FILLER_50_41 ();
 FILLCELL_X1 FILLER_50_43 ();
 FILLCELL_X2 FILLER_50_65 ();
 FILLCELL_X2 FILLER_50_74 ();
 FILLCELL_X2 FILLER_50_83 ();
 FILLCELL_X8 FILLER_50_90 ();
 FILLCELL_X2 FILLER_50_106 ();
 FILLCELL_X1 FILLER_50_108 ();
 FILLCELL_X2 FILLER_50_113 ();
 FILLCELL_X8 FILLER_50_159 ();
 FILLCELL_X4 FILLER_50_167 ();
 FILLCELL_X2 FILLER_50_171 ();
 FILLCELL_X2 FILLER_50_194 ();
 FILLCELL_X8 FILLER_50_233 ();
 FILLCELL_X4 FILLER_50_241 ();
 FILLCELL_X1 FILLER_50_262 ();
 FILLCELL_X2 FILLER_50_271 ();
 FILLCELL_X8 FILLER_50_287 ();
 FILLCELL_X4 FILLER_50_295 ();
 FILLCELL_X1 FILLER_50_299 ();
 FILLCELL_X8 FILLER_50_308 ();
 FILLCELL_X2 FILLER_50_316 ();
 FILLCELL_X8 FILLER_50_335 ();
 FILLCELL_X2 FILLER_50_343 ();
 FILLCELL_X2 FILLER_50_352 ();
 FILLCELL_X2 FILLER_50_357 ();
 FILLCELL_X1 FILLER_50_359 ();
 FILLCELL_X4 FILLER_50_374 ();
 FILLCELL_X1 FILLER_50_378 ();
 FILLCELL_X2 FILLER_50_386 ();
 FILLCELL_X1 FILLER_50_388 ();
 FILLCELL_X16 FILLER_50_396 ();
 FILLCELL_X1 FILLER_50_412 ();
 FILLCELL_X1 FILLER_50_420 ();
 FILLCELL_X2 FILLER_50_444 ();
 FILLCELL_X1 FILLER_50_446 ();
 FILLCELL_X2 FILLER_50_450 ();
 FILLCELL_X1 FILLER_50_452 ();
 FILLCELL_X8 FILLER_50_456 ();
 FILLCELL_X2 FILLER_50_464 ();
 FILLCELL_X1 FILLER_50_466 ();
 FILLCELL_X16 FILLER_50_472 ();
 FILLCELL_X1 FILLER_50_488 ();
 FILLCELL_X4 FILLER_50_492 ();
 FILLCELL_X2 FILLER_50_496 ();
 FILLCELL_X8 FILLER_50_503 ();
 FILLCELL_X4 FILLER_50_511 ();
 FILLCELL_X1 FILLER_50_515 ();
 FILLCELL_X16 FILLER_50_520 ();
 FILLCELL_X8 FILLER_50_536 ();
 FILLCELL_X4 FILLER_50_544 ();
 FILLCELL_X2 FILLER_50_548 ();
 FILLCELL_X1 FILLER_50_550 ();
 FILLCELL_X32 FILLER_50_557 ();
 FILLCELL_X2 FILLER_50_589 ();
 FILLCELL_X8 FILLER_50_596 ();
 FILLCELL_X4 FILLER_50_604 ();
 FILLCELL_X8 FILLER_50_621 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X8 FILLER_50_632 ();
 FILLCELL_X4 FILLER_50_640 ();
 FILLCELL_X8 FILLER_50_661 ();
 FILLCELL_X2 FILLER_50_669 ();
 FILLCELL_X4 FILLER_50_679 ();
 FILLCELL_X1 FILLER_50_690 ();
 FILLCELL_X16 FILLER_50_699 ();
 FILLCELL_X4 FILLER_50_715 ();
 FILLCELL_X2 FILLER_50_719 ();
 FILLCELL_X1 FILLER_50_721 ();
 FILLCELL_X8 FILLER_50_725 ();
 FILLCELL_X4 FILLER_50_733 ();
 FILLCELL_X1 FILLER_50_737 ();
 FILLCELL_X1 FILLER_50_796 ();
 FILLCELL_X4 FILLER_51_1 ();
 FILLCELL_X4 FILLER_51_26 ();
 FILLCELL_X1 FILLER_51_34 ();
 FILLCELL_X1 FILLER_51_38 ();
 FILLCELL_X8 FILLER_51_46 ();
 FILLCELL_X4 FILLER_51_54 ();
 FILLCELL_X2 FILLER_51_58 ();
 FILLCELL_X16 FILLER_51_126 ();
 FILLCELL_X4 FILLER_51_167 ();
 FILLCELL_X1 FILLER_51_171 ();
 FILLCELL_X16 FILLER_51_186 ();
 FILLCELL_X4 FILLER_51_202 ();
 FILLCELL_X2 FILLER_51_206 ();
 FILLCELL_X1 FILLER_51_208 ();
 FILLCELL_X4 FILLER_51_213 ();
 FILLCELL_X4 FILLER_51_220 ();
 FILLCELL_X2 FILLER_51_224 ();
 FILLCELL_X1 FILLER_51_226 ();
 FILLCELL_X2 FILLER_51_232 ();
 FILLCELL_X1 FILLER_51_234 ();
 FILLCELL_X1 FILLER_51_242 ();
 FILLCELL_X4 FILLER_51_246 ();
 FILLCELL_X2 FILLER_51_250 ();
 FILLCELL_X1 FILLER_51_252 ();
 FILLCELL_X4 FILLER_51_256 ();
 FILLCELL_X1 FILLER_51_281 ();
 FILLCELL_X4 FILLER_51_289 ();
 FILLCELL_X8 FILLER_51_310 ();
 FILLCELL_X4 FILLER_51_318 ();
 FILLCELL_X2 FILLER_51_322 ();
 FILLCELL_X1 FILLER_51_324 ();
 FILLCELL_X8 FILLER_51_328 ();
 FILLCELL_X1 FILLER_51_336 ();
 FILLCELL_X2 FILLER_51_341 ();
 FILLCELL_X1 FILLER_51_343 ();
 FILLCELL_X8 FILLER_51_396 ();
 FILLCELL_X4 FILLER_51_404 ();
 FILLCELL_X2 FILLER_51_408 ();
 FILLCELL_X1 FILLER_51_434 ();
 FILLCELL_X1 FILLER_51_439 ();
 FILLCELL_X2 FILLER_51_443 ();
 FILLCELL_X1 FILLER_51_445 ();
 FILLCELL_X2 FILLER_51_461 ();
 FILLCELL_X2 FILLER_51_466 ();
 FILLCELL_X8 FILLER_51_475 ();
 FILLCELL_X4 FILLER_51_487 ();
 FILLCELL_X16 FILLER_51_501 ();
 FILLCELL_X2 FILLER_51_528 ();
 FILLCELL_X1 FILLER_51_532 ();
 FILLCELL_X4 FILLER_51_538 ();
 FILLCELL_X2 FILLER_51_553 ();
 FILLCELL_X1 FILLER_51_560 ();
 FILLCELL_X4 FILLER_51_563 ();
 FILLCELL_X1 FILLER_51_567 ();
 FILLCELL_X8 FILLER_51_572 ();
 FILLCELL_X1 FILLER_51_580 ();
 FILLCELL_X1 FILLER_51_585 ();
 FILLCELL_X2 FILLER_51_595 ();
 FILLCELL_X2 FILLER_51_599 ();
 FILLCELL_X4 FILLER_51_612 ();
 FILLCELL_X1 FILLER_51_616 ();
 FILLCELL_X4 FILLER_51_641 ();
 FILLCELL_X2 FILLER_51_645 ();
 FILLCELL_X1 FILLER_51_647 ();
 FILLCELL_X1 FILLER_51_656 ();
 FILLCELL_X8 FILLER_51_664 ();
 FILLCELL_X4 FILLER_51_672 ();
 FILLCELL_X4 FILLER_51_680 ();
 FILLCELL_X2 FILLER_51_684 ();
 FILLCELL_X4 FILLER_51_697 ();
 FILLCELL_X1 FILLER_51_704 ();
 FILLCELL_X2 FILLER_51_709 ();
 FILLCELL_X1 FILLER_51_720 ();
 FILLCELL_X2 FILLER_51_735 ();
 FILLCELL_X2 FILLER_51_754 ();
 FILLCELL_X1 FILLER_51_756 ();
 FILLCELL_X16 FILLER_51_761 ();
 FILLCELL_X1 FILLER_51_777 ();
 FILLCELL_X1 FILLER_51_785 ();
 FILLCELL_X1 FILLER_51_796 ();
 FILLCELL_X4 FILLER_51_810 ();
 FILLCELL_X16 FILLER_52_1 ();
 FILLCELL_X4 FILLER_52_17 ();
 FILLCELL_X1 FILLER_52_21 ();
 FILLCELL_X8 FILLER_52_39 ();
 FILLCELL_X2 FILLER_52_47 ();
 FILLCELL_X2 FILLER_52_70 ();
 FILLCELL_X1 FILLER_52_72 ();
 FILLCELL_X16 FILLER_52_80 ();
 FILLCELL_X8 FILLER_52_96 ();
 FILLCELL_X4 FILLER_52_104 ();
 FILLCELL_X2 FILLER_52_108 ();
 FILLCELL_X1 FILLER_52_110 ();
 FILLCELL_X16 FILLER_52_114 ();
 FILLCELL_X2 FILLER_52_130 ();
 FILLCELL_X1 FILLER_52_132 ();
 FILLCELL_X16 FILLER_52_137 ();
 FILLCELL_X4 FILLER_52_153 ();
 FILLCELL_X1 FILLER_52_157 ();
 FILLCELL_X16 FILLER_52_172 ();
 FILLCELL_X4 FILLER_52_188 ();
 FILLCELL_X1 FILLER_52_192 ();
 FILLCELL_X2 FILLER_52_197 ();
 FILLCELL_X1 FILLER_52_199 ();
 FILLCELL_X8 FILLER_52_220 ();
 FILLCELL_X4 FILLER_52_228 ();
 FILLCELL_X2 FILLER_52_232 ();
 FILLCELL_X4 FILLER_52_258 ();
 FILLCELL_X1 FILLER_52_262 ();
 FILLCELL_X32 FILLER_52_270 ();
 FILLCELL_X2 FILLER_52_302 ();
 FILLCELL_X1 FILLER_52_304 ();
 FILLCELL_X16 FILLER_52_342 ();
 FILLCELL_X2 FILLER_52_358 ();
 FILLCELL_X1 FILLER_52_360 ();
 FILLCELL_X32 FILLER_52_368 ();
 FILLCELL_X2 FILLER_52_400 ();
 FILLCELL_X4 FILLER_52_416 ();
 FILLCELL_X2 FILLER_52_420 ();
 FILLCELL_X1 FILLER_52_422 ();
 FILLCELL_X2 FILLER_52_447 ();
 FILLCELL_X1 FILLER_52_449 ();
 FILLCELL_X2 FILLER_52_467 ();
 FILLCELL_X2 FILLER_52_505 ();
 FILLCELL_X4 FILLER_52_530 ();
 FILLCELL_X1 FILLER_52_538 ();
 FILLCELL_X1 FILLER_52_544 ();
 FILLCELL_X1 FILLER_52_554 ();
 FILLCELL_X1 FILLER_52_572 ();
 FILLCELL_X1 FILLER_52_590 ();
 FILLCELL_X1 FILLER_52_595 ();
 FILLCELL_X1 FILLER_52_607 ();
 FILLCELL_X16 FILLER_52_612 ();
 FILLCELL_X2 FILLER_52_628 ();
 FILLCELL_X1 FILLER_52_630 ();
 FILLCELL_X1 FILLER_52_632 ();
 FILLCELL_X4 FILLER_52_638 ();
 FILLCELL_X1 FILLER_52_642 ();
 FILLCELL_X8 FILLER_52_660 ();
 FILLCELL_X4 FILLER_52_668 ();
 FILLCELL_X1 FILLER_52_672 ();
 FILLCELL_X2 FILLER_52_690 ();
 FILLCELL_X1 FILLER_52_692 ();
 FILLCELL_X2 FILLER_52_700 ();
 FILLCELL_X8 FILLER_52_706 ();
 FILLCELL_X2 FILLER_52_714 ();
 FILLCELL_X2 FILLER_52_733 ();
 FILLCELL_X1 FILLER_52_742 ();
 FILLCELL_X4 FILLER_52_753 ();
 FILLCELL_X4 FILLER_52_762 ();
 FILLCELL_X2 FILLER_52_766 ();
 FILLCELL_X8 FILLER_52_775 ();
 FILLCELL_X4 FILLER_52_783 ();
 FILLCELL_X2 FILLER_52_787 ();
 FILLCELL_X1 FILLER_52_789 ();
 FILLCELL_X8 FILLER_52_793 ();
 FILLCELL_X1 FILLER_52_810 ();
 FILLCELL_X8 FILLER_53_1 ();
 FILLCELL_X4 FILLER_53_9 ();
 FILLCELL_X2 FILLER_53_13 ();
 FILLCELL_X1 FILLER_53_38 ();
 FILLCELL_X8 FILLER_53_44 ();
 FILLCELL_X2 FILLER_53_52 ();
 FILLCELL_X1 FILLER_53_54 ();
 FILLCELL_X2 FILLER_53_59 ();
 FILLCELL_X2 FILLER_53_69 ();
 FILLCELL_X1 FILLER_53_71 ();
 FILLCELL_X8 FILLER_53_79 ();
 FILLCELL_X4 FILLER_53_87 ();
 FILLCELL_X1 FILLER_53_91 ();
 FILLCELL_X2 FILLER_53_101 ();
 FILLCELL_X16 FILLER_53_107 ();
 FILLCELL_X2 FILLER_53_123 ();
 FILLCELL_X1 FILLER_53_125 ();
 FILLCELL_X1 FILLER_53_150 ();
 FILLCELL_X8 FILLER_53_172 ();
 FILLCELL_X1 FILLER_53_180 ();
 FILLCELL_X1 FILLER_53_211 ();
 FILLCELL_X4 FILLER_53_219 ();
 FILLCELL_X8 FILLER_53_226 ();
 FILLCELL_X4 FILLER_53_234 ();
 FILLCELL_X2 FILLER_53_238 ();
 FILLCELL_X2 FILLER_53_247 ();
 FILLCELL_X1 FILLER_53_249 ();
 FILLCELL_X8 FILLER_53_277 ();
 FILLCELL_X4 FILLER_53_285 ();
 FILLCELL_X1 FILLER_53_293 ();
 FILLCELL_X1 FILLER_53_297 ();
 FILLCELL_X1 FILLER_53_301 ();
 FILLCELL_X1 FILLER_53_309 ();
 FILLCELL_X2 FILLER_53_320 ();
 FILLCELL_X8 FILLER_53_329 ();
 FILLCELL_X4 FILLER_53_337 ();
 FILLCELL_X1 FILLER_53_341 ();
 FILLCELL_X2 FILLER_53_350 ();
 FILLCELL_X8 FILLER_53_360 ();
 FILLCELL_X2 FILLER_53_368 ();
 FILLCELL_X2 FILLER_53_380 ();
 FILLCELL_X4 FILLER_53_402 ();
 FILLCELL_X2 FILLER_53_406 ();
 FILLCELL_X32 FILLER_53_440 ();
 FILLCELL_X8 FILLER_53_472 ();
 FILLCELL_X4 FILLER_53_480 ();
 FILLCELL_X8 FILLER_53_487 ();
 FILLCELL_X1 FILLER_53_495 ();
 FILLCELL_X16 FILLER_53_501 ();
 FILLCELL_X2 FILLER_53_517 ();
 FILLCELL_X1 FILLER_53_526 ();
 FILLCELL_X1 FILLER_53_531 ();
 FILLCELL_X4 FILLER_53_539 ();
 FILLCELL_X1 FILLER_53_543 ();
 FILLCELL_X1 FILLER_53_549 ();
 FILLCELL_X1 FILLER_53_555 ();
 FILLCELL_X16 FILLER_53_563 ();
 FILLCELL_X8 FILLER_53_579 ();
 FILLCELL_X1 FILLER_53_602 ();
 FILLCELL_X8 FILLER_53_641 ();
 FILLCELL_X2 FILLER_53_656 ();
 FILLCELL_X4 FILLER_53_665 ();
 FILLCELL_X2 FILLER_53_669 ();
 FILLCELL_X1 FILLER_53_671 ();
 FILLCELL_X4 FILLER_53_693 ();
 FILLCELL_X1 FILLER_53_697 ();
 FILLCELL_X1 FILLER_53_702 ();
 FILLCELL_X8 FILLER_53_707 ();
 FILLCELL_X4 FILLER_53_729 ();
 FILLCELL_X2 FILLER_53_733 ();
 FILLCELL_X1 FILLER_53_754 ();
 FILLCELL_X4 FILLER_53_757 ();
 FILLCELL_X4 FILLER_53_781 ();
 FILLCELL_X2 FILLER_53_785 ();
 FILLCELL_X4 FILLER_53_807 ();
 FILLCELL_X16 FILLER_54_1 ();
 FILLCELL_X8 FILLER_54_17 ();
 FILLCELL_X4 FILLER_54_25 ();
 FILLCELL_X8 FILLER_54_40 ();
 FILLCELL_X2 FILLER_54_48 ();
 FILLCELL_X1 FILLER_54_50 ();
 FILLCELL_X2 FILLER_54_68 ();
 FILLCELL_X4 FILLER_54_84 ();
 FILLCELL_X2 FILLER_54_88 ();
 FILLCELL_X1 FILLER_54_90 ();
 FILLCELL_X2 FILLER_54_108 ();
 FILLCELL_X2 FILLER_54_133 ();
 FILLCELL_X1 FILLER_54_138 ();
 FILLCELL_X2 FILLER_54_142 ();
 FILLCELL_X8 FILLER_54_151 ();
 FILLCELL_X2 FILLER_54_166 ();
 FILLCELL_X1 FILLER_54_168 ();
 FILLCELL_X32 FILLER_54_176 ();
 FILLCELL_X2 FILLER_54_208 ();
 FILLCELL_X1 FILLER_54_210 ();
 FILLCELL_X1 FILLER_54_228 ();
 FILLCELL_X2 FILLER_54_327 ();
 FILLCELL_X8 FILLER_54_336 ();
 FILLCELL_X2 FILLER_54_344 ();
 FILLCELL_X4 FILLER_54_363 ();
 FILLCELL_X1 FILLER_54_367 ();
 FILLCELL_X16 FILLER_54_378 ();
 FILLCELL_X8 FILLER_54_401 ();
 FILLCELL_X2 FILLER_54_409 ();
 FILLCELL_X1 FILLER_54_411 ();
 FILLCELL_X2 FILLER_54_431 ();
 FILLCELL_X4 FILLER_54_437 ();
 FILLCELL_X1 FILLER_54_441 ();
 FILLCELL_X4 FILLER_54_448 ();
 FILLCELL_X8 FILLER_54_459 ();
 FILLCELL_X2 FILLER_54_467 ();
 FILLCELL_X1 FILLER_54_483 ();
 FILLCELL_X2 FILLER_54_488 ();
 FILLCELL_X4 FILLER_54_505 ();
 FILLCELL_X2 FILLER_54_509 ();
 FILLCELL_X1 FILLER_54_511 ();
 FILLCELL_X2 FILLER_54_523 ();
 FILLCELL_X2 FILLER_54_527 ();
 FILLCELL_X8 FILLER_54_533 ();
 FILLCELL_X1 FILLER_54_548 ();
 FILLCELL_X2 FILLER_54_574 ();
 FILLCELL_X1 FILLER_54_576 ();
 FILLCELL_X4 FILLER_54_591 ();
 FILLCELL_X4 FILLER_54_612 ();
 FILLCELL_X1 FILLER_54_632 ();
 FILLCELL_X4 FILLER_54_640 ();
 FILLCELL_X16 FILLER_54_661 ();
 FILLCELL_X1 FILLER_54_677 ();
 FILLCELL_X8 FILLER_54_682 ();
 FILLCELL_X2 FILLER_54_690 ();
 FILLCELL_X1 FILLER_54_692 ();
 FILLCELL_X4 FILLER_54_718 ();
 FILLCELL_X1 FILLER_54_722 ();
 FILLCELL_X8 FILLER_54_727 ();
 FILLCELL_X4 FILLER_54_735 ();
 FILLCELL_X2 FILLER_54_739 ();
 FILLCELL_X2 FILLER_54_748 ();
 FILLCELL_X8 FILLER_54_753 ();
 FILLCELL_X1 FILLER_54_765 ();
 FILLCELL_X16 FILLER_54_769 ();
 FILLCELL_X2 FILLER_54_795 ();
 FILLCELL_X4 FILLER_55_1 ();
 FILLCELL_X4 FILLER_55_9 ();
 FILLCELL_X4 FILLER_55_18 ();
 FILLCELL_X1 FILLER_55_22 ();
 FILLCELL_X1 FILLER_55_43 ();
 FILLCELL_X2 FILLER_55_61 ();
 FILLCELL_X1 FILLER_55_77 ();
 FILLCELL_X4 FILLER_55_92 ();
 FILLCELL_X2 FILLER_55_96 ();
 FILLCELL_X1 FILLER_55_98 ();
 FILLCELL_X16 FILLER_55_123 ();
 FILLCELL_X4 FILLER_55_139 ();
 FILLCELL_X1 FILLER_55_143 ();
 FILLCELL_X8 FILLER_55_156 ();
 FILLCELL_X4 FILLER_55_164 ();
 FILLCELL_X1 FILLER_55_168 ();
 FILLCELL_X1 FILLER_55_176 ();
 FILLCELL_X16 FILLER_55_190 ();
 FILLCELL_X4 FILLER_55_206 ();
 FILLCELL_X1 FILLER_55_210 ();
 FILLCELL_X16 FILLER_55_214 ();
 FILLCELL_X4 FILLER_55_230 ();
 FILLCELL_X2 FILLER_55_244 ();
 FILLCELL_X16 FILLER_55_263 ();
 FILLCELL_X1 FILLER_55_279 ();
 FILLCELL_X16 FILLER_55_287 ();
 FILLCELL_X4 FILLER_55_303 ();
 FILLCELL_X2 FILLER_55_307 ();
 FILLCELL_X1 FILLER_55_309 ();
 FILLCELL_X1 FILLER_55_334 ();
 FILLCELL_X16 FILLER_55_338 ();
 FILLCELL_X4 FILLER_55_354 ();
 FILLCELL_X8 FILLER_55_379 ();
 FILLCELL_X1 FILLER_55_387 ();
 FILLCELL_X1 FILLER_55_406 ();
 FILLCELL_X2 FILLER_55_424 ();
 FILLCELL_X1 FILLER_55_426 ();
 FILLCELL_X1 FILLER_55_447 ();
 FILLCELL_X8 FILLER_55_465 ();
 FILLCELL_X4 FILLER_55_473 ();
 FILLCELL_X2 FILLER_55_501 ();
 FILLCELL_X1 FILLER_55_519 ();
 FILLCELL_X2 FILLER_55_524 ();
 FILLCELL_X1 FILLER_55_530 ();
 FILLCELL_X2 FILLER_55_535 ();
 FILLCELL_X1 FILLER_55_537 ();
 FILLCELL_X2 FILLER_55_551 ();
 FILLCELL_X1 FILLER_55_553 ();
 FILLCELL_X4 FILLER_55_559 ();
 FILLCELL_X2 FILLER_55_569 ();
 FILLCELL_X1 FILLER_55_571 ();
 FILLCELL_X8 FILLER_55_589 ();
 FILLCELL_X2 FILLER_55_597 ();
 FILLCELL_X1 FILLER_55_599 ();
 FILLCELL_X2 FILLER_55_604 ();
 FILLCELL_X32 FILLER_55_610 ();
 FILLCELL_X8 FILLER_55_642 ();
 FILLCELL_X4 FILLER_55_650 ();
 FILLCELL_X1 FILLER_55_654 ();
 FILLCELL_X2 FILLER_55_675 ();
 FILLCELL_X1 FILLER_55_677 ();
 FILLCELL_X4 FILLER_55_685 ();
 FILLCELL_X4 FILLER_55_696 ();
 FILLCELL_X2 FILLER_55_700 ();
 FILLCELL_X1 FILLER_55_723 ();
 FILLCELL_X1 FILLER_55_731 ();
 FILLCELL_X4 FILLER_55_775 ();
 FILLCELL_X2 FILLER_55_779 ();
 FILLCELL_X1 FILLER_55_781 ();
 FILLCELL_X2 FILLER_55_809 ();
 FILLCELL_X4 FILLER_56_32 ();
 FILLCELL_X2 FILLER_56_36 ();
 FILLCELL_X8 FILLER_56_51 ();
 FILLCELL_X8 FILLER_56_63 ();
 FILLCELL_X1 FILLER_56_71 ();
 FILLCELL_X16 FILLER_56_82 ();
 FILLCELL_X8 FILLER_56_98 ();
 FILLCELL_X1 FILLER_56_106 ();
 FILLCELL_X1 FILLER_56_114 ();
 FILLCELL_X16 FILLER_56_118 ();
 FILLCELL_X4 FILLER_56_144 ();
 FILLCELL_X2 FILLER_56_148 ();
 FILLCELL_X4 FILLER_56_172 ();
 FILLCELL_X1 FILLER_56_176 ();
 FILLCELL_X1 FILLER_56_216 ();
 FILLCELL_X2 FILLER_56_221 ();
 FILLCELL_X1 FILLER_56_223 ();
 FILLCELL_X8 FILLER_56_227 ();
 FILLCELL_X2 FILLER_56_235 ();
 FILLCELL_X1 FILLER_56_241 ();
 FILLCELL_X1 FILLER_56_249 ();
 FILLCELL_X2 FILLER_56_254 ();
 FILLCELL_X2 FILLER_56_259 ();
 FILLCELL_X8 FILLER_56_264 ();
 FILLCELL_X4 FILLER_56_272 ();
 FILLCELL_X2 FILLER_56_276 ();
 FILLCELL_X1 FILLER_56_278 ();
 FILLCELL_X8 FILLER_56_291 ();
 FILLCELL_X4 FILLER_56_299 ();
 FILLCELL_X1 FILLER_56_307 ();
 FILLCELL_X2 FILLER_56_312 ();
 FILLCELL_X1 FILLER_56_314 ();
 FILLCELL_X2 FILLER_56_329 ();
 FILLCELL_X1 FILLER_56_331 ();
 FILLCELL_X16 FILLER_56_335 ();
 FILLCELL_X8 FILLER_56_351 ();
 FILLCELL_X1 FILLER_56_359 ();
 FILLCELL_X4 FILLER_56_367 ();
 FILLCELL_X2 FILLER_56_371 ();
 FILLCELL_X1 FILLER_56_373 ();
 FILLCELL_X1 FILLER_56_393 ();
 FILLCELL_X1 FILLER_56_413 ();
 FILLCELL_X16 FILLER_56_417 ();
 FILLCELL_X1 FILLER_56_433 ();
 FILLCELL_X8 FILLER_56_437 ();
 FILLCELL_X4 FILLER_56_445 ();
 FILLCELL_X1 FILLER_56_449 ();
 FILLCELL_X8 FILLER_56_474 ();
 FILLCELL_X2 FILLER_56_482 ();
 FILLCELL_X1 FILLER_56_484 ();
 FILLCELL_X1 FILLER_56_488 ();
 FILLCELL_X2 FILLER_56_492 ();
 FILLCELL_X8 FILLER_56_499 ();
 FILLCELL_X1 FILLER_56_507 ();
 FILLCELL_X2 FILLER_56_522 ();
 FILLCELL_X8 FILLER_56_541 ();
 FILLCELL_X4 FILLER_56_549 ();
 FILLCELL_X4 FILLER_56_570 ();
 FILLCELL_X2 FILLER_56_574 ();
 FILLCELL_X32 FILLER_56_589 ();
 FILLCELL_X2 FILLER_56_621 ();
 FILLCELL_X1 FILLER_56_623 ();
 FILLCELL_X8 FILLER_56_632 ();
 FILLCELL_X4 FILLER_56_640 ();
 FILLCELL_X2 FILLER_56_644 ();
 FILLCELL_X1 FILLER_56_646 ();
 FILLCELL_X1 FILLER_56_651 ();
 FILLCELL_X1 FILLER_56_664 ();
 FILLCELL_X2 FILLER_56_682 ();
 FILLCELL_X16 FILLER_56_705 ();
 FILLCELL_X8 FILLER_56_721 ();
 FILLCELL_X2 FILLER_56_729 ();
 FILLCELL_X1 FILLER_56_731 ();
 FILLCELL_X4 FILLER_56_745 ();
 FILLCELL_X2 FILLER_56_749 ();
 FILLCELL_X4 FILLER_56_756 ();
 FILLCELL_X2 FILLER_56_760 ();
 FILLCELL_X16 FILLER_56_770 ();
 FILLCELL_X2 FILLER_56_786 ();
 FILLCELL_X1 FILLER_56_788 ();
 FILLCELL_X8 FILLER_56_798 ();
 FILLCELL_X4 FILLER_56_806 ();
 FILLCELL_X1 FILLER_56_810 ();
 FILLCELL_X2 FILLER_57_1 ();
 FILLCELL_X4 FILLER_57_10 ();
 FILLCELL_X4 FILLER_57_18 ();
 FILLCELL_X2 FILLER_57_22 ();
 FILLCELL_X2 FILLER_57_27 ();
 FILLCELL_X4 FILLER_57_33 ();
 FILLCELL_X2 FILLER_57_57 ();
 FILLCELL_X1 FILLER_57_59 ();
 FILLCELL_X16 FILLER_57_74 ();
 FILLCELL_X1 FILLER_57_90 ();
 FILLCELL_X2 FILLER_57_102 ();
 FILLCELL_X1 FILLER_57_108 ();
 FILLCELL_X1 FILLER_57_113 ();
 FILLCELL_X8 FILLER_57_117 ();
 FILLCELL_X2 FILLER_57_125 ();
 FILLCELL_X2 FILLER_57_174 ();
 FILLCELL_X1 FILLER_57_176 ();
 FILLCELL_X2 FILLER_57_181 ();
 FILLCELL_X4 FILLER_57_189 ();
 FILLCELL_X1 FILLER_57_250 ();
 FILLCELL_X2 FILLER_57_275 ();
 FILLCELL_X2 FILLER_57_280 ();
 FILLCELL_X1 FILLER_57_282 ();
 FILLCELL_X1 FILLER_57_289 ();
 FILLCELL_X2 FILLER_57_295 ();
 FILLCELL_X2 FILLER_57_328 ();
 FILLCELL_X8 FILLER_57_337 ();
 FILLCELL_X4 FILLER_57_345 ();
 FILLCELL_X1 FILLER_57_349 ();
 FILLCELL_X1 FILLER_57_364 ();
 FILLCELL_X1 FILLER_57_368 ();
 FILLCELL_X2 FILLER_57_430 ();
 FILLCELL_X1 FILLER_57_432 ();
 FILLCELL_X1 FILLER_57_437 ();
 FILLCELL_X8 FILLER_57_444 ();
 FILLCELL_X2 FILLER_57_452 ();
 FILLCELL_X8 FILLER_57_459 ();
 FILLCELL_X2 FILLER_57_467 ();
 FILLCELL_X4 FILLER_57_472 ();
 FILLCELL_X2 FILLER_57_476 ();
 FILLCELL_X1 FILLER_57_490 ();
 FILLCELL_X8 FILLER_57_494 ();
 FILLCELL_X2 FILLER_57_502 ();
 FILLCELL_X4 FILLER_57_509 ();
 FILLCELL_X1 FILLER_57_513 ();
 FILLCELL_X16 FILLER_57_521 ();
 FILLCELL_X8 FILLER_57_537 ();
 FILLCELL_X1 FILLER_57_545 ();
 FILLCELL_X4 FILLER_57_551 ();
 FILLCELL_X16 FILLER_57_560 ();
 FILLCELL_X4 FILLER_57_576 ();
 FILLCELL_X1 FILLER_57_584 ();
 FILLCELL_X4 FILLER_57_592 ();
 FILLCELL_X2 FILLER_57_596 ();
 FILLCELL_X1 FILLER_57_598 ();
 FILLCELL_X2 FILLER_57_607 ();
 FILLCELL_X4 FILLER_57_664 ();
 FILLCELL_X1 FILLER_57_668 ();
 FILLCELL_X2 FILLER_57_681 ();
 FILLCELL_X1 FILLER_57_683 ();
 FILLCELL_X4 FILLER_57_701 ();
 FILLCELL_X1 FILLER_57_705 ();
 FILLCELL_X2 FILLER_57_709 ();
 FILLCELL_X8 FILLER_57_718 ();
 FILLCELL_X1 FILLER_57_726 ();
 FILLCELL_X8 FILLER_57_734 ();
 FILLCELL_X2 FILLER_57_742 ();
 FILLCELL_X1 FILLER_57_744 ();
 FILLCELL_X16 FILLER_57_752 ();
 FILLCELL_X8 FILLER_57_768 ();
 FILLCELL_X2 FILLER_57_776 ();
 FILLCELL_X1 FILLER_57_778 ();
 FILLCELL_X4 FILLER_57_796 ();
 FILLCELL_X1 FILLER_57_800 ();
 FILLCELL_X2 FILLER_57_804 ();
 FILLCELL_X1 FILLER_57_806 ();
 FILLCELL_X4 FILLER_57_810 ();
 FILLCELL_X4 FILLER_58_6 ();
 FILLCELL_X2 FILLER_58_10 ();
 FILLCELL_X1 FILLER_58_12 ();
 FILLCELL_X2 FILLER_58_20 ();
 FILLCELL_X1 FILLER_58_22 ();
 FILLCELL_X1 FILLER_58_40 ();
 FILLCELL_X2 FILLER_58_48 ();
 FILLCELL_X1 FILLER_58_50 ();
 FILLCELL_X2 FILLER_58_55 ();
 FILLCELL_X4 FILLER_58_61 ();
 FILLCELL_X2 FILLER_58_79 ();
 FILLCELL_X2 FILLER_58_88 ();
 FILLCELL_X1 FILLER_58_90 ();
 FILLCELL_X1 FILLER_58_108 ();
 FILLCELL_X2 FILLER_58_126 ();
 FILLCELL_X4 FILLER_58_144 ();
 FILLCELL_X4 FILLER_58_175 ();
 FILLCELL_X2 FILLER_58_191 ();
 FILLCELL_X1 FILLER_58_193 ();
 FILLCELL_X1 FILLER_58_204 ();
 FILLCELL_X2 FILLER_58_209 ();
 FILLCELL_X16 FILLER_58_214 ();
 FILLCELL_X8 FILLER_58_230 ();
 FILLCELL_X1 FILLER_58_238 ();
 FILLCELL_X2 FILLER_58_249 ();
 FILLCELL_X1 FILLER_58_251 ();
 FILLCELL_X8 FILLER_58_259 ();
 FILLCELL_X2 FILLER_58_267 ();
 FILLCELL_X1 FILLER_58_269 ();
 FILLCELL_X2 FILLER_58_277 ();
 FILLCELL_X1 FILLER_58_286 ();
 FILLCELL_X1 FILLER_58_294 ();
 FILLCELL_X1 FILLER_58_302 ();
 FILLCELL_X8 FILLER_58_310 ();
 FILLCELL_X1 FILLER_58_325 ();
 FILLCELL_X1 FILLER_58_333 ();
 FILLCELL_X1 FILLER_58_341 ();
 FILLCELL_X2 FILLER_58_354 ();
 FILLCELL_X2 FILLER_58_369 ();
 FILLCELL_X4 FILLER_58_376 ();
 FILLCELL_X1 FILLER_58_380 ();
 FILLCELL_X2 FILLER_58_404 ();
 FILLCELL_X1 FILLER_58_406 ();
 FILLCELL_X1 FILLER_58_431 ();
 FILLCELL_X1 FILLER_58_437 ();
 FILLCELL_X1 FILLER_58_441 ();
 FILLCELL_X1 FILLER_58_447 ();
 FILLCELL_X1 FILLER_58_452 ();
 FILLCELL_X4 FILLER_58_456 ();
 FILLCELL_X2 FILLER_58_460 ();
 FILLCELL_X1 FILLER_58_462 ();
 FILLCELL_X2 FILLER_58_467 ();
 FILLCELL_X8 FILLER_58_494 ();
 FILLCELL_X1 FILLER_58_502 ();
 FILLCELL_X4 FILLER_58_535 ();
 FILLCELL_X2 FILLER_58_539 ();
 FILLCELL_X4 FILLER_58_546 ();
 FILLCELL_X8 FILLER_58_556 ();
 FILLCELL_X4 FILLER_58_569 ();
 FILLCELL_X1 FILLER_58_573 ();
 FILLCELL_X1 FILLER_58_593 ();
 FILLCELL_X1 FILLER_58_611 ();
 FILLCELL_X1 FILLER_58_617 ();
 FILLCELL_X2 FILLER_58_628 ();
 FILLCELL_X1 FILLER_58_630 ();
 FILLCELL_X8 FILLER_58_632 ();
 FILLCELL_X2 FILLER_58_640 ();
 FILLCELL_X16 FILLER_58_647 ();
 FILLCELL_X8 FILLER_58_675 ();
 FILLCELL_X2 FILLER_58_683 ();
 FILLCELL_X1 FILLER_58_685 ();
 FILLCELL_X8 FILLER_58_690 ();
 FILLCELL_X1 FILLER_58_706 ();
 FILLCELL_X2 FILLER_58_718 ();
 FILLCELL_X2 FILLER_58_723 ();
 FILLCELL_X4 FILLER_58_728 ();
 FILLCELL_X2 FILLER_58_732 ();
 FILLCELL_X1 FILLER_58_734 ();
 FILLCELL_X4 FILLER_58_742 ();
 FILLCELL_X8 FILLER_58_753 ();
 FILLCELL_X4 FILLER_58_761 ();
 FILLCELL_X1 FILLER_58_765 ();
 FILLCELL_X1 FILLER_58_777 ();
 FILLCELL_X2 FILLER_58_795 ();
 FILLCELL_X8 FILLER_58_803 ();
 FILLCELL_X2 FILLER_58_811 ();
 FILLCELL_X1 FILLER_58_813 ();
 FILLCELL_X16 FILLER_59_1 ();
 FILLCELL_X4 FILLER_59_17 ();
 FILLCELL_X2 FILLER_59_28 ();
 FILLCELL_X1 FILLER_59_30 ();
 FILLCELL_X4 FILLER_59_38 ();
 FILLCELL_X2 FILLER_59_42 ();
 FILLCELL_X4 FILLER_59_65 ();
 FILLCELL_X1 FILLER_59_69 ();
 FILLCELL_X8 FILLER_59_77 ();
 FILLCELL_X4 FILLER_59_85 ();
 FILLCELL_X1 FILLER_59_89 ();
 FILLCELL_X4 FILLER_59_104 ();
 FILLCELL_X2 FILLER_59_108 ();
 FILLCELL_X1 FILLER_59_110 ();
 FILLCELL_X2 FILLER_59_114 ();
 FILLCELL_X1 FILLER_59_123 ();
 FILLCELL_X2 FILLER_59_131 ();
 FILLCELL_X2 FILLER_59_140 ();
 FILLCELL_X8 FILLER_59_149 ();
 FILLCELL_X2 FILLER_59_157 ();
 FILLCELL_X4 FILLER_59_198 ();
 FILLCELL_X1 FILLER_59_202 ();
 FILLCELL_X1 FILLER_59_211 ();
 FILLCELL_X32 FILLER_59_215 ();
 FILLCELL_X4 FILLER_59_247 ();
 FILLCELL_X1 FILLER_59_251 ();
 FILLCELL_X4 FILLER_59_256 ();
 FILLCELL_X2 FILLER_59_260 ();
 FILLCELL_X4 FILLER_59_265 ();
 FILLCELL_X1 FILLER_59_269 ();
 FILLCELL_X16 FILLER_59_275 ();
 FILLCELL_X4 FILLER_59_291 ();
 FILLCELL_X2 FILLER_59_295 ();
 FILLCELL_X1 FILLER_59_297 ();
 FILLCELL_X4 FILLER_59_315 ();
 FILLCELL_X1 FILLER_59_319 ();
 FILLCELL_X8 FILLER_59_340 ();
 FILLCELL_X4 FILLER_59_351 ();
 FILLCELL_X4 FILLER_59_359 ();
 FILLCELL_X1 FILLER_59_363 ();
 FILLCELL_X16 FILLER_59_374 ();
 FILLCELL_X8 FILLER_59_390 ();
 FILLCELL_X1 FILLER_59_398 ();
 FILLCELL_X4 FILLER_59_418 ();
 FILLCELL_X1 FILLER_59_422 ();
 FILLCELL_X1 FILLER_59_435 ();
 FILLCELL_X1 FILLER_59_443 ();
 FILLCELL_X8 FILLER_59_478 ();
 FILLCELL_X4 FILLER_59_486 ();
 FILLCELL_X1 FILLER_59_490 ();
 FILLCELL_X1 FILLER_59_505 ();
 FILLCELL_X2 FILLER_59_543 ();
 FILLCELL_X2 FILLER_59_551 ();
 FILLCELL_X2 FILLER_59_558 ();
 FILLCELL_X2 FILLER_59_562 ();
 FILLCELL_X8 FILLER_59_568 ();
 FILLCELL_X2 FILLER_59_576 ();
 FILLCELL_X1 FILLER_59_578 ();
 FILLCELL_X2 FILLER_59_583 ();
 FILLCELL_X1 FILLER_59_585 ();
 FILLCELL_X1 FILLER_59_601 ();
 FILLCELL_X8 FILLER_59_621 ();
 FILLCELL_X4 FILLER_59_629 ();
 FILLCELL_X4 FILLER_59_687 ();
 FILLCELL_X2 FILLER_59_691 ();
 FILLCELL_X1 FILLER_59_693 ();
 FILLCELL_X8 FILLER_59_699 ();
 FILLCELL_X2 FILLER_59_707 ();
 FILLCELL_X1 FILLER_59_727 ();
 FILLCELL_X1 FILLER_59_732 ();
 FILLCELL_X1 FILLER_59_753 ();
 FILLCELL_X1 FILLER_59_778 ();
 FILLCELL_X1 FILLER_59_796 ();
 FILLCELL_X8 FILLER_60_1 ();
 FILLCELL_X4 FILLER_60_9 ();
 FILLCELL_X1 FILLER_60_13 ();
 FILLCELL_X8 FILLER_60_18 ();
 FILLCELL_X4 FILLER_60_26 ();
 FILLCELL_X1 FILLER_60_30 ();
 FILLCELL_X2 FILLER_60_35 ();
 FILLCELL_X4 FILLER_60_49 ();
 FILLCELL_X2 FILLER_60_57 ();
 FILLCELL_X1 FILLER_60_59 ();
 FILLCELL_X1 FILLER_60_64 ();
 FILLCELL_X4 FILLER_60_69 ();
 FILLCELL_X32 FILLER_60_78 ();
 FILLCELL_X4 FILLER_60_110 ();
 FILLCELL_X2 FILLER_60_114 ();
 FILLCELL_X1 FILLER_60_116 ();
 FILLCELL_X8 FILLER_60_124 ();
 FILLCELL_X2 FILLER_60_132 ();
 FILLCELL_X16 FILLER_60_148 ();
 FILLCELL_X2 FILLER_60_164 ();
 FILLCELL_X1 FILLER_60_166 ();
 FILLCELL_X2 FILLER_60_225 ();
 FILLCELL_X1 FILLER_60_227 ();
 FILLCELL_X2 FILLER_60_231 ();
 FILLCELL_X1 FILLER_60_233 ();
 FILLCELL_X1 FILLER_60_249 ();
 FILLCELL_X4 FILLER_60_267 ();
 FILLCELL_X4 FILLER_60_278 ();
 FILLCELL_X8 FILLER_60_289 ();
 FILLCELL_X1 FILLER_60_301 ();
 FILLCELL_X16 FILLER_60_308 ();
 FILLCELL_X1 FILLER_60_324 ();
 FILLCELL_X2 FILLER_60_329 ();
 FILLCELL_X8 FILLER_60_334 ();
 FILLCELL_X2 FILLER_60_342 ();
 FILLCELL_X1 FILLER_60_344 ();
 FILLCELL_X4 FILLER_60_349 ();
 FILLCELL_X4 FILLER_60_356 ();
 FILLCELL_X8 FILLER_60_374 ();
 FILLCELL_X8 FILLER_60_395 ();
 FILLCELL_X4 FILLER_60_403 ();
 FILLCELL_X2 FILLER_60_407 ();
 FILLCELL_X1 FILLER_60_409 ();
 FILLCELL_X1 FILLER_60_417 ();
 FILLCELL_X2 FILLER_60_422 ();
 FILLCELL_X1 FILLER_60_447 ();
 FILLCELL_X1 FILLER_60_451 ();
 FILLCELL_X16 FILLER_60_455 ();
 FILLCELL_X8 FILLER_60_471 ();
 FILLCELL_X2 FILLER_60_493 ();
 FILLCELL_X1 FILLER_60_495 ();
 FILLCELL_X2 FILLER_60_507 ();
 FILLCELL_X1 FILLER_60_509 ();
 FILLCELL_X2 FILLER_60_514 ();
 FILLCELL_X8 FILLER_60_520 ();
 FILLCELL_X2 FILLER_60_528 ();
 FILLCELL_X2 FILLER_60_538 ();
 FILLCELL_X1 FILLER_60_540 ();
 FILLCELL_X1 FILLER_60_544 ();
 FILLCELL_X2 FILLER_60_562 ();
 FILLCELL_X4 FILLER_60_573 ();
 FILLCELL_X1 FILLER_60_577 ();
 FILLCELL_X2 FILLER_60_585 ();
 FILLCELL_X4 FILLER_60_591 ();
 FILLCELL_X4 FILLER_60_600 ();
 FILLCELL_X2 FILLER_60_604 ();
 FILLCELL_X8 FILLER_60_617 ();
 FILLCELL_X4 FILLER_60_625 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X8 FILLER_60_640 ();
 FILLCELL_X4 FILLER_60_648 ();
 FILLCELL_X1 FILLER_60_652 ();
 FILLCELL_X8 FILLER_60_661 ();
 FILLCELL_X2 FILLER_60_672 ();
 FILLCELL_X4 FILLER_60_681 ();
 FILLCELL_X4 FILLER_60_689 ();
 FILLCELL_X1 FILLER_60_707 ();
 FILLCELL_X4 FILLER_60_717 ();
 FILLCELL_X1 FILLER_60_721 ();
 FILLCELL_X4 FILLER_60_729 ();
 FILLCELL_X2 FILLER_60_733 ();
 FILLCELL_X1 FILLER_60_735 ();
 FILLCELL_X4 FILLER_60_739 ();
 FILLCELL_X2 FILLER_60_743 ();
 FILLCELL_X1 FILLER_60_745 ();
 FILLCELL_X8 FILLER_60_757 ();
 FILLCELL_X2 FILLER_60_765 ();
 FILLCELL_X16 FILLER_60_773 ();
 FILLCELL_X4 FILLER_60_789 ();
 FILLCELL_X2 FILLER_60_799 ();
 FILLCELL_X16 FILLER_61_1 ();
 FILLCELL_X8 FILLER_61_17 ();
 FILLCELL_X8 FILLER_61_45 ();
 FILLCELL_X2 FILLER_61_53 ();
 FILLCELL_X1 FILLER_61_79 ();
 FILLCELL_X8 FILLER_61_104 ();
 FILLCELL_X1 FILLER_61_112 ();
 FILLCELL_X2 FILLER_61_120 ();
 FILLCELL_X8 FILLER_61_125 ();
 FILLCELL_X4 FILLER_61_133 ();
 FILLCELL_X2 FILLER_61_137 ();
 FILLCELL_X8 FILLER_61_146 ();
 FILLCELL_X4 FILLER_61_154 ();
 FILLCELL_X2 FILLER_61_158 ();
 FILLCELL_X16 FILLER_61_167 ();
 FILLCELL_X1 FILLER_61_183 ();
 FILLCELL_X16 FILLER_61_188 ();
 FILLCELL_X2 FILLER_61_211 ();
 FILLCELL_X4 FILLER_61_230 ();
 FILLCELL_X2 FILLER_61_251 ();
 FILLCELL_X1 FILLER_61_256 ();
 FILLCELL_X1 FILLER_61_260 ();
 FILLCELL_X1 FILLER_61_264 ();
 FILLCELL_X2 FILLER_61_272 ();
 FILLCELL_X2 FILLER_61_281 ();
 FILLCELL_X1 FILLER_61_283 ();
 FILLCELL_X2 FILLER_61_291 ();
 FILLCELL_X1 FILLER_61_293 ();
 FILLCELL_X2 FILLER_61_326 ();
 FILLCELL_X1 FILLER_61_328 ();
 FILLCELL_X2 FILLER_61_332 ();
 FILLCELL_X1 FILLER_61_334 ();
 FILLCELL_X4 FILLER_61_342 ();
 FILLCELL_X4 FILLER_61_363 ();
 FILLCELL_X2 FILLER_61_367 ();
 FILLCELL_X2 FILLER_61_390 ();
 FILLCELL_X1 FILLER_61_392 ();
 FILLCELL_X2 FILLER_61_423 ();
 FILLCELL_X8 FILLER_61_432 ();
 FILLCELL_X4 FILLER_61_440 ();
 FILLCELL_X1 FILLER_61_447 ();
 FILLCELL_X2 FILLER_61_451 ();
 FILLCELL_X1 FILLER_61_456 ();
 FILLCELL_X2 FILLER_61_461 ();
 FILLCELL_X16 FILLER_61_466 ();
 FILLCELL_X2 FILLER_61_482 ();
 FILLCELL_X1 FILLER_61_491 ();
 FILLCELL_X8 FILLER_61_495 ();
 FILLCELL_X1 FILLER_61_520 ();
 FILLCELL_X4 FILLER_61_542 ();
 FILLCELL_X2 FILLER_61_571 ();
 FILLCELL_X1 FILLER_61_573 ();
 FILLCELL_X2 FILLER_61_582 ();
 FILLCELL_X1 FILLER_61_584 ();
 FILLCELL_X16 FILLER_61_602 ();
 FILLCELL_X8 FILLER_61_635 ();
 FILLCELL_X2 FILLER_61_643 ();
 FILLCELL_X1 FILLER_61_645 ();
 FILLCELL_X16 FILLER_61_654 ();
 FILLCELL_X8 FILLER_61_670 ();
 FILLCELL_X2 FILLER_61_682 ();
 FILLCELL_X1 FILLER_61_695 ();
 FILLCELL_X1 FILLER_61_699 ();
 FILLCELL_X1 FILLER_61_704 ();
 FILLCELL_X1 FILLER_61_709 ();
 FILLCELL_X1 FILLER_61_713 ();
 FILLCELL_X4 FILLER_61_718 ();
 FILLCELL_X2 FILLER_61_722 ();
 FILLCELL_X1 FILLER_61_724 ();
 FILLCELL_X4 FILLER_61_732 ();
 FILLCELL_X1 FILLER_61_736 ();
 FILLCELL_X8 FILLER_61_751 ();
 FILLCELL_X2 FILLER_61_759 ();
 FILLCELL_X2 FILLER_61_768 ();
 FILLCELL_X1 FILLER_61_770 ();
 FILLCELL_X8 FILLER_61_773 ();
 FILLCELL_X4 FILLER_61_781 ();
 FILLCELL_X1 FILLER_61_795 ();
 FILLCELL_X4 FILLER_61_803 ();
 FILLCELL_X16 FILLER_62_1 ();
 FILLCELL_X8 FILLER_62_17 ();
 FILLCELL_X4 FILLER_62_28 ();
 FILLCELL_X1 FILLER_62_32 ();
 FILLCELL_X2 FILLER_62_41 ();
 FILLCELL_X1 FILLER_62_43 ();
 FILLCELL_X2 FILLER_62_61 ();
 FILLCELL_X4 FILLER_62_70 ();
 FILLCELL_X2 FILLER_62_74 ();
 FILLCELL_X1 FILLER_62_76 ();
 FILLCELL_X8 FILLER_62_84 ();
 FILLCELL_X2 FILLER_62_92 ();
 FILLCELL_X4 FILLER_62_98 ();
 FILLCELL_X4 FILLER_62_106 ();
 FILLCELL_X1 FILLER_62_113 ();
 FILLCELL_X8 FILLER_62_131 ();
 FILLCELL_X1 FILLER_62_146 ();
 FILLCELL_X2 FILLER_62_168 ();
 FILLCELL_X2 FILLER_62_194 ();
 FILLCELL_X4 FILLER_62_199 ();
 FILLCELL_X16 FILLER_62_216 ();
 FILLCELL_X4 FILLER_62_232 ();
 FILLCELL_X2 FILLER_62_236 ();
 FILLCELL_X2 FILLER_62_262 ();
 FILLCELL_X8 FILLER_62_285 ();
 FILLCELL_X4 FILLER_62_293 ();
 FILLCELL_X1 FILLER_62_297 ();
 FILLCELL_X1 FILLER_62_301 ();
 FILLCELL_X2 FILLER_62_322 ();
 FILLCELL_X4 FILLER_62_327 ();
 FILLCELL_X2 FILLER_62_331 ();
 FILLCELL_X8 FILLER_62_350 ();
 FILLCELL_X1 FILLER_62_358 ();
 FILLCELL_X8 FILLER_62_366 ();
 FILLCELL_X2 FILLER_62_374 ();
 FILLCELL_X2 FILLER_62_379 ();
 FILLCELL_X2 FILLER_62_394 ();
 FILLCELL_X1 FILLER_62_396 ();
 FILLCELL_X2 FILLER_62_401 ();
 FILLCELL_X1 FILLER_62_410 ();
 FILLCELL_X2 FILLER_62_414 ();
 FILLCELL_X1 FILLER_62_416 ();
 FILLCELL_X2 FILLER_62_424 ();
 FILLCELL_X2 FILLER_62_447 ();
 FILLCELL_X4 FILLER_62_473 ();
 FILLCELL_X2 FILLER_62_477 ();
 FILLCELL_X16 FILLER_62_496 ();
 FILLCELL_X2 FILLER_62_512 ();
 FILLCELL_X8 FILLER_62_521 ();
 FILLCELL_X4 FILLER_62_529 ();
 FILLCELL_X4 FILLER_62_542 ();
 FILLCELL_X2 FILLER_62_546 ();
 FILLCELL_X1 FILLER_62_554 ();
 FILLCELL_X4 FILLER_62_560 ();
 FILLCELL_X2 FILLER_62_596 ();
 FILLCELL_X16 FILLER_62_614 ();
 FILLCELL_X1 FILLER_62_630 ();
 FILLCELL_X4 FILLER_62_634 ();
 FILLCELL_X2 FILLER_62_638 ();
 FILLCELL_X1 FILLER_62_640 ();
 FILLCELL_X4 FILLER_62_658 ();
 FILLCELL_X2 FILLER_62_662 ();
 FILLCELL_X2 FILLER_62_667 ();
 FILLCELL_X2 FILLER_62_713 ();
 FILLCELL_X8 FILLER_62_720 ();
 FILLCELL_X1 FILLER_62_728 ();
 FILLCELL_X4 FILLER_62_777 ();
 FILLCELL_X1 FILLER_62_781 ();
 FILLCELL_X4 FILLER_63_1 ();
 FILLCELL_X2 FILLER_63_5 ();
 FILLCELL_X8 FILLER_63_44 ();
 FILLCELL_X2 FILLER_63_52 ();
 FILLCELL_X2 FILLER_63_62 ();
 FILLCELL_X1 FILLER_63_64 ();
 FILLCELL_X2 FILLER_63_72 ();
 FILLCELL_X4 FILLER_63_79 ();
 FILLCELL_X8 FILLER_63_90 ();
 FILLCELL_X2 FILLER_63_106 ();
 FILLCELL_X1 FILLER_63_108 ();
 FILLCELL_X1 FILLER_63_116 ();
 FILLCELL_X4 FILLER_63_124 ();
 FILLCELL_X2 FILLER_63_128 ();
 FILLCELL_X16 FILLER_63_139 ();
 FILLCELL_X2 FILLER_63_155 ();
 FILLCELL_X16 FILLER_63_171 ();
 FILLCELL_X8 FILLER_63_187 ();
 FILLCELL_X2 FILLER_63_195 ();
 FILLCELL_X1 FILLER_63_197 ();
 FILLCELL_X4 FILLER_63_201 ();
 FILLCELL_X2 FILLER_63_205 ();
 FILLCELL_X1 FILLER_63_211 ();
 FILLCELL_X2 FILLER_63_215 ();
 FILLCELL_X1 FILLER_63_221 ();
 FILLCELL_X8 FILLER_63_227 ();
 FILLCELL_X2 FILLER_63_235 ();
 FILLCELL_X1 FILLER_63_241 ();
 FILLCELL_X1 FILLER_63_245 ();
 FILLCELL_X4 FILLER_63_253 ();
 FILLCELL_X2 FILLER_63_257 ();
 FILLCELL_X8 FILLER_63_266 ();
 FILLCELL_X1 FILLER_63_274 ();
 FILLCELL_X8 FILLER_63_282 ();
 FILLCELL_X4 FILLER_63_290 ();
 FILLCELL_X2 FILLER_63_294 ();
 FILLCELL_X1 FILLER_63_296 ();
 FILLCELL_X2 FILLER_63_310 ();
 FILLCELL_X1 FILLER_63_312 ();
 FILLCELL_X8 FILLER_63_324 ();
 FILLCELL_X2 FILLER_63_332 ();
 FILLCELL_X16 FILLER_63_337 ();
 FILLCELL_X8 FILLER_63_353 ();
 FILLCELL_X4 FILLER_63_361 ();
 FILLCELL_X4 FILLER_63_372 ();
 FILLCELL_X2 FILLER_63_376 ();
 FILLCELL_X16 FILLER_63_391 ();
 FILLCELL_X8 FILLER_63_407 ();
 FILLCELL_X4 FILLER_63_418 ();
 FILLCELL_X1 FILLER_63_422 ();
 FILLCELL_X8 FILLER_63_426 ();
 FILLCELL_X4 FILLER_63_434 ();
 FILLCELL_X2 FILLER_63_438 ();
 FILLCELL_X8 FILLER_63_443 ();
 FILLCELL_X2 FILLER_63_451 ();
 FILLCELL_X8 FILLER_63_477 ();
 FILLCELL_X1 FILLER_63_488 ();
 FILLCELL_X2 FILLER_63_503 ();
 FILLCELL_X1 FILLER_63_505 ();
 FILLCELL_X8 FILLER_63_516 ();
 FILLCELL_X4 FILLER_63_526 ();
 FILLCELL_X2 FILLER_63_530 ();
 FILLCELL_X1 FILLER_63_532 ();
 FILLCELL_X32 FILLER_63_546 ();
 FILLCELL_X16 FILLER_63_578 ();
 FILLCELL_X4 FILLER_63_615 ();
 FILLCELL_X1 FILLER_63_619 ();
 FILLCELL_X4 FILLER_63_625 ();
 FILLCELL_X2 FILLER_63_629 ();
 FILLCELL_X8 FILLER_63_638 ();
 FILLCELL_X4 FILLER_63_646 ();
 FILLCELL_X2 FILLER_63_650 ();
 FILLCELL_X2 FILLER_63_659 ();
 FILLCELL_X8 FILLER_63_672 ();
 FILLCELL_X2 FILLER_63_684 ();
 FILLCELL_X1 FILLER_63_686 ();
 FILLCELL_X4 FILLER_63_691 ();
 FILLCELL_X2 FILLER_63_695 ();
 FILLCELL_X2 FILLER_63_701 ();
 FILLCELL_X2 FILLER_63_707 ();
 FILLCELL_X1 FILLER_63_709 ();
 FILLCELL_X2 FILLER_63_717 ();
 FILLCELL_X1 FILLER_63_719 ();
 FILLCELL_X2 FILLER_63_727 ();
 FILLCELL_X1 FILLER_63_729 ();
 FILLCELL_X4 FILLER_63_743 ();
 FILLCELL_X8 FILLER_63_753 ();
 FILLCELL_X2 FILLER_63_761 ();
 FILLCELL_X1 FILLER_63_763 ();
 FILLCELL_X4 FILLER_63_767 ();
 FILLCELL_X2 FILLER_63_771 ();
 FILLCELL_X1 FILLER_63_773 ();
 FILLCELL_X1 FILLER_63_791 ();
 FILLCELL_X16 FILLER_64_1 ();
 FILLCELL_X8 FILLER_64_17 ();
 FILLCELL_X1 FILLER_64_42 ();
 FILLCELL_X1 FILLER_64_48 ();
 FILLCELL_X4 FILLER_64_70 ();
 FILLCELL_X2 FILLER_64_81 ();
 FILLCELL_X1 FILLER_64_83 ();
 FILLCELL_X2 FILLER_64_125 ();
 FILLCELL_X4 FILLER_64_153 ();
 FILLCELL_X2 FILLER_64_173 ();
 FILLCELL_X1 FILLER_64_175 ();
 FILLCELL_X4 FILLER_64_191 ();
 FILLCELL_X1 FILLER_64_195 ();
 FILLCELL_X1 FILLER_64_213 ();
 FILLCELL_X2 FILLER_64_231 ();
 FILLCELL_X1 FILLER_64_257 ();
 FILLCELL_X4 FILLER_64_265 ();
 FILLCELL_X1 FILLER_64_274 ();
 FILLCELL_X4 FILLER_64_288 ();
 FILLCELL_X2 FILLER_64_292 ();
 FILLCELL_X1 FILLER_64_294 ();
 FILLCELL_X2 FILLER_64_306 ();
 FILLCELL_X1 FILLER_64_308 ();
 FILLCELL_X2 FILLER_64_330 ();
 FILLCELL_X1 FILLER_64_332 ();
 FILLCELL_X8 FILLER_64_337 ();
 FILLCELL_X2 FILLER_64_345 ();
 FILLCELL_X2 FILLER_64_352 ();
 FILLCELL_X4 FILLER_64_358 ();
 FILLCELL_X2 FILLER_64_362 ();
 FILLCELL_X1 FILLER_64_371 ();
 FILLCELL_X16 FILLER_64_379 ();
 FILLCELL_X8 FILLER_64_395 ();
 FILLCELL_X2 FILLER_64_403 ();
 FILLCELL_X8 FILLER_64_426 ();
 FILLCELL_X1 FILLER_64_434 ();
 FILLCELL_X2 FILLER_64_445 ();
 FILLCELL_X2 FILLER_64_450 ();
 FILLCELL_X16 FILLER_64_455 ();
 FILLCELL_X2 FILLER_64_471 ();
 FILLCELL_X4 FILLER_64_487 ();
 FILLCELL_X1 FILLER_64_491 ();
 FILLCELL_X4 FILLER_64_497 ();
 FILLCELL_X4 FILLER_64_504 ();
 FILLCELL_X2 FILLER_64_532 ();
 FILLCELL_X4 FILLER_64_539 ();
 FILLCELL_X1 FILLER_64_543 ();
 FILLCELL_X1 FILLER_64_548 ();
 FILLCELL_X1 FILLER_64_555 ();
 FILLCELL_X2 FILLER_64_561 ();
 FILLCELL_X2 FILLER_64_576 ();
 FILLCELL_X2 FILLER_64_585 ();
 FILLCELL_X2 FILLER_64_602 ();
 FILLCELL_X4 FILLER_64_608 ();
 FILLCELL_X2 FILLER_64_629 ();
 FILLCELL_X2 FILLER_64_632 ();
 FILLCELL_X1 FILLER_64_641 ();
 FILLCELL_X2 FILLER_64_644 ();
 FILLCELL_X1 FILLER_64_675 ();
 FILLCELL_X2 FILLER_64_729 ();
 FILLCELL_X8 FILLER_64_752 ();
 FILLCELL_X4 FILLER_64_760 ();
 FILLCELL_X1 FILLER_64_766 ();
 FILLCELL_X4 FILLER_64_770 ();
 FILLCELL_X2 FILLER_64_774 ();
 FILLCELL_X1 FILLER_64_776 ();
 FILLCELL_X4 FILLER_64_787 ();
 FILLCELL_X4 FILLER_64_807 ();
 FILLCELL_X2 FILLER_64_811 ();
 FILLCELL_X1 FILLER_64_813 ();
 FILLCELL_X8 FILLER_65_1 ();
 FILLCELL_X4 FILLER_65_9 ();
 FILLCELL_X2 FILLER_65_13 ();
 FILLCELL_X1 FILLER_65_15 ();
 FILLCELL_X16 FILLER_65_21 ();
 FILLCELL_X2 FILLER_65_37 ();
 FILLCELL_X8 FILLER_65_43 ();
 FILLCELL_X1 FILLER_65_51 ();
 FILLCELL_X1 FILLER_65_60 ();
 FILLCELL_X8 FILLER_65_65 ();
 FILLCELL_X1 FILLER_65_73 ();
 FILLCELL_X2 FILLER_65_88 ();
 FILLCELL_X16 FILLER_65_97 ();
 FILLCELL_X8 FILLER_65_113 ();
 FILLCELL_X1 FILLER_65_121 ();
 FILLCELL_X4 FILLER_65_129 ();
 FILLCELL_X2 FILLER_65_133 ();
 FILLCELL_X2 FILLER_65_145 ();
 FILLCELL_X1 FILLER_65_147 ();
 FILLCELL_X2 FILLER_65_152 ();
 FILLCELL_X1 FILLER_65_154 ();
 FILLCELL_X4 FILLER_65_158 ();
 FILLCELL_X2 FILLER_65_169 ();
 FILLCELL_X16 FILLER_65_195 ();
 FILLCELL_X4 FILLER_65_211 ();
 FILLCELL_X1 FILLER_65_215 ();
 FILLCELL_X4 FILLER_65_221 ();
 FILLCELL_X16 FILLER_65_228 ();
 FILLCELL_X2 FILLER_65_244 ();
 FILLCELL_X1 FILLER_65_246 ();
 FILLCELL_X16 FILLER_65_268 ();
 FILLCELL_X4 FILLER_65_284 ();
 FILLCELL_X1 FILLER_65_288 ();
 FILLCELL_X1 FILLER_65_313 ();
 FILLCELL_X4 FILLER_65_350 ();
 FILLCELL_X4 FILLER_65_358 ();
 FILLCELL_X2 FILLER_65_362 ();
 FILLCELL_X1 FILLER_65_364 ();
 FILLCELL_X2 FILLER_65_382 ();
 FILLCELL_X8 FILLER_65_397 ();
 FILLCELL_X4 FILLER_65_405 ();
 FILLCELL_X2 FILLER_65_409 ();
 FILLCELL_X4 FILLER_65_418 ();
 FILLCELL_X2 FILLER_65_425 ();
 FILLCELL_X2 FILLER_65_432 ();
 FILLCELL_X1 FILLER_65_434 ();
 FILLCELL_X4 FILLER_65_452 ();
 FILLCELL_X1 FILLER_65_456 ();
 FILLCELL_X16 FILLER_65_469 ();
 FILLCELL_X4 FILLER_65_489 ();
 FILLCELL_X2 FILLER_65_493 ();
 FILLCELL_X1 FILLER_65_495 ();
 FILLCELL_X8 FILLER_65_501 ();
 FILLCELL_X1 FILLER_65_509 ();
 FILLCELL_X4 FILLER_65_514 ();
 FILLCELL_X2 FILLER_65_518 ();
 FILLCELL_X4 FILLER_65_524 ();
 FILLCELL_X1 FILLER_65_532 ();
 FILLCELL_X2 FILLER_65_537 ();
 FILLCELL_X1 FILLER_65_539 ();
 FILLCELL_X2 FILLER_65_547 ();
 FILLCELL_X1 FILLER_65_549 ();
 FILLCELL_X2 FILLER_65_556 ();
 FILLCELL_X2 FILLER_65_575 ();
 FILLCELL_X2 FILLER_65_584 ();
 FILLCELL_X8 FILLER_65_590 ();
 FILLCELL_X1 FILLER_65_598 ();
 FILLCELL_X8 FILLER_65_608 ();
 FILLCELL_X1 FILLER_65_616 ();
 FILLCELL_X2 FILLER_65_624 ();
 FILLCELL_X1 FILLER_65_630 ();
 FILLCELL_X16 FILLER_65_644 ();
 FILLCELL_X4 FILLER_65_660 ();
 FILLCELL_X1 FILLER_65_664 ();
 FILLCELL_X16 FILLER_65_672 ();
 FILLCELL_X2 FILLER_65_688 ();
 FILLCELL_X1 FILLER_65_697 ();
 FILLCELL_X2 FILLER_65_705 ();
 FILLCELL_X4 FILLER_65_711 ();
 FILLCELL_X1 FILLER_65_724 ();
 FILLCELL_X4 FILLER_65_732 ();
 FILLCELL_X2 FILLER_65_736 ();
 FILLCELL_X1 FILLER_65_738 ();
 FILLCELL_X4 FILLER_65_756 ();
 FILLCELL_X2 FILLER_65_760 ();
 FILLCELL_X8 FILLER_65_769 ();
 FILLCELL_X1 FILLER_65_777 ();
 FILLCELL_X2 FILLER_65_792 ();
 FILLCELL_X16 FILLER_66_1 ();
 FILLCELL_X2 FILLER_66_22 ();
 FILLCELL_X1 FILLER_66_24 ();
 FILLCELL_X2 FILLER_66_45 ();
 FILLCELL_X2 FILLER_66_69 ();
 FILLCELL_X1 FILLER_66_71 ();
 FILLCELL_X8 FILLER_66_93 ();
 FILLCELL_X4 FILLER_66_101 ();
 FILLCELL_X2 FILLER_66_105 ();
 FILLCELL_X1 FILLER_66_107 ();
 FILLCELL_X4 FILLER_66_113 ();
 FILLCELL_X2 FILLER_66_117 ();
 FILLCELL_X1 FILLER_66_119 ();
 FILLCELL_X2 FILLER_66_141 ();
 FILLCELL_X32 FILLER_66_160 ();
 FILLCELL_X8 FILLER_66_192 ();
 FILLCELL_X4 FILLER_66_200 ();
 FILLCELL_X16 FILLER_66_208 ();
 FILLCELL_X8 FILLER_66_224 ();
 FILLCELL_X4 FILLER_66_232 ();
 FILLCELL_X4 FILLER_66_249 ();
 FILLCELL_X2 FILLER_66_253 ();
 FILLCELL_X32 FILLER_66_267 ();
 FILLCELL_X8 FILLER_66_299 ();
 FILLCELL_X1 FILLER_66_311 ();
 FILLCELL_X4 FILLER_66_319 ();
 FILLCELL_X1 FILLER_66_323 ();
 FILLCELL_X1 FILLER_66_331 ();
 FILLCELL_X2 FILLER_66_335 ();
 FILLCELL_X1 FILLER_66_337 ();
 FILLCELL_X2 FILLER_66_368 ();
 FILLCELL_X1 FILLER_66_370 ();
 FILLCELL_X8 FILLER_66_426 ();
 FILLCELL_X2 FILLER_66_434 ();
 FILLCELL_X1 FILLER_66_436 ();
 FILLCELL_X8 FILLER_66_441 ();
 FILLCELL_X1 FILLER_66_449 ();
 FILLCELL_X2 FILLER_66_470 ();
 FILLCELL_X1 FILLER_66_472 ();
 FILLCELL_X8 FILLER_66_504 ();
 FILLCELL_X16 FILLER_66_524 ();
 FILLCELL_X8 FILLER_66_557 ();
 FILLCELL_X2 FILLER_66_565 ();
 FILLCELL_X2 FILLER_66_572 ();
 FILLCELL_X4 FILLER_66_598 ();
 FILLCELL_X2 FILLER_66_602 ();
 FILLCELL_X1 FILLER_66_604 ();
 FILLCELL_X4 FILLER_66_612 ();
 FILLCELL_X1 FILLER_66_616 ();
 FILLCELL_X1 FILLER_66_632 ();
 FILLCELL_X4 FILLER_66_652 ();
 FILLCELL_X2 FILLER_66_656 ();
 FILLCELL_X2 FILLER_66_663 ();
 FILLCELL_X1 FILLER_66_665 ();
 FILLCELL_X4 FILLER_66_673 ();
 FILLCELL_X2 FILLER_66_677 ();
 FILLCELL_X1 FILLER_66_679 ();
 FILLCELL_X8 FILLER_66_685 ();
 FILLCELL_X1 FILLER_66_693 ();
 FILLCELL_X8 FILLER_66_701 ();
 FILLCELL_X8 FILLER_66_728 ();
 FILLCELL_X4 FILLER_66_736 ();
 FILLCELL_X1 FILLER_66_740 ();
 FILLCELL_X8 FILLER_66_748 ();
 FILLCELL_X4 FILLER_66_756 ();
 FILLCELL_X2 FILLER_66_797 ();
 FILLCELL_X8 FILLER_66_803 ();
 FILLCELL_X2 FILLER_67_1 ();
 FILLCELL_X1 FILLER_67_3 ();
 FILLCELL_X16 FILLER_67_11 ();
 FILLCELL_X2 FILLER_67_27 ();
 FILLCELL_X2 FILLER_67_34 ();
 FILLCELL_X1 FILLER_67_36 ();
 FILLCELL_X16 FILLER_67_42 ();
 FILLCELL_X4 FILLER_67_58 ();
 FILLCELL_X16 FILLER_67_67 ();
 FILLCELL_X8 FILLER_67_83 ();
 FILLCELL_X4 FILLER_67_91 ();
 FILLCELL_X2 FILLER_67_95 ();
 FILLCELL_X1 FILLER_67_97 ();
 FILLCELL_X2 FILLER_67_120 ();
 FILLCELL_X1 FILLER_67_122 ();
 FILLCELL_X4 FILLER_67_128 ();
 FILLCELL_X2 FILLER_67_132 ();
 FILLCELL_X8 FILLER_67_137 ();
 FILLCELL_X2 FILLER_67_145 ();
 FILLCELL_X1 FILLER_67_147 ();
 FILLCELL_X8 FILLER_67_158 ();
 FILLCELL_X2 FILLER_67_166 ();
 FILLCELL_X8 FILLER_67_189 ();
 FILLCELL_X8 FILLER_67_200 ();
 FILLCELL_X2 FILLER_67_211 ();
 FILLCELL_X2 FILLER_67_220 ();
 FILLCELL_X1 FILLER_67_222 ();
 FILLCELL_X4 FILLER_67_226 ();
 FILLCELL_X1 FILLER_67_230 ();
 FILLCELL_X2 FILLER_67_251 ();
 FILLCELL_X1 FILLER_67_253 ();
 FILLCELL_X2 FILLER_67_288 ();
 FILLCELL_X1 FILLER_67_290 ();
 FILLCELL_X16 FILLER_67_308 ();
 FILLCELL_X4 FILLER_67_324 ();
 FILLCELL_X1 FILLER_67_328 ();
 FILLCELL_X4 FILLER_67_342 ();
 FILLCELL_X1 FILLER_67_346 ();
 FILLCELL_X32 FILLER_67_352 ();
 FILLCELL_X4 FILLER_67_384 ();
 FILLCELL_X1 FILLER_67_388 ();
 FILLCELL_X1 FILLER_67_418 ();
 FILLCELL_X8 FILLER_67_422 ();
 FILLCELL_X16 FILLER_67_460 ();
 FILLCELL_X1 FILLER_67_476 ();
 FILLCELL_X4 FILLER_67_484 ();
 FILLCELL_X2 FILLER_67_488 ();
 FILLCELL_X1 FILLER_67_490 ();
 FILLCELL_X4 FILLER_67_506 ();
 FILLCELL_X2 FILLER_67_513 ();
 FILLCELL_X2 FILLER_67_527 ();
 FILLCELL_X16 FILLER_67_538 ();
 FILLCELL_X8 FILLER_67_554 ();
 FILLCELL_X16 FILLER_67_569 ();
 FILLCELL_X2 FILLER_67_585 ();
 FILLCELL_X4 FILLER_67_591 ();
 FILLCELL_X2 FILLER_67_616 ();
 FILLCELL_X1 FILLER_67_618 ();
 FILLCELL_X2 FILLER_67_633 ();
 FILLCELL_X1 FILLER_67_635 ();
 FILLCELL_X4 FILLER_67_643 ();
 FILLCELL_X2 FILLER_67_647 ();
 FILLCELL_X2 FILLER_67_662 ();
 FILLCELL_X1 FILLER_67_664 ();
 FILLCELL_X8 FILLER_67_672 ();
 FILLCELL_X1 FILLER_67_680 ();
 FILLCELL_X4 FILLER_67_688 ();
 FILLCELL_X2 FILLER_67_692 ();
 FILLCELL_X1 FILLER_67_694 ();
 FILLCELL_X8 FILLER_67_707 ();
 FILLCELL_X4 FILLER_67_715 ();
 FILLCELL_X2 FILLER_67_719 ();
 FILLCELL_X1 FILLER_67_721 ();
 FILLCELL_X16 FILLER_67_727 ();
 FILLCELL_X8 FILLER_67_743 ();
 FILLCELL_X4 FILLER_67_751 ();
 FILLCELL_X2 FILLER_67_755 ();
 FILLCELL_X16 FILLER_67_762 ();
 FILLCELL_X8 FILLER_67_778 ();
 FILLCELL_X4 FILLER_67_794 ();
 FILLCELL_X2 FILLER_67_798 ();
 FILLCELL_X1 FILLER_67_800 ();
 FILLCELL_X8 FILLER_67_804 ();
 FILLCELL_X2 FILLER_67_812 ();
 FILLCELL_X16 FILLER_68_37 ();
 FILLCELL_X4 FILLER_68_72 ();
 FILLCELL_X1 FILLER_68_76 ();
 FILLCELL_X4 FILLER_68_84 ();
 FILLCELL_X1 FILLER_68_88 ();
 FILLCELL_X2 FILLER_68_110 ();
 FILLCELL_X8 FILLER_68_123 ();
 FILLCELL_X1 FILLER_68_131 ();
 FILLCELL_X4 FILLER_68_146 ();
 FILLCELL_X1 FILLER_68_150 ();
 FILLCELL_X1 FILLER_68_158 ();
 FILLCELL_X1 FILLER_68_166 ();
 FILLCELL_X8 FILLER_68_188 ();
 FILLCELL_X1 FILLER_68_196 ();
 FILLCELL_X8 FILLER_68_231 ();
 FILLCELL_X4 FILLER_68_239 ();
 FILLCELL_X2 FILLER_68_243 ();
 FILLCELL_X8 FILLER_68_249 ();
 FILLCELL_X2 FILLER_68_257 ();
 FILLCELL_X1 FILLER_68_259 ();
 FILLCELL_X2 FILLER_68_264 ();
 FILLCELL_X8 FILLER_68_287 ();
 FILLCELL_X4 FILLER_68_295 ();
 FILLCELL_X32 FILLER_68_316 ();
 FILLCELL_X2 FILLER_68_348 ();
 FILLCELL_X1 FILLER_68_350 ();
 FILLCELL_X4 FILLER_68_355 ();
 FILLCELL_X2 FILLER_68_363 ();
 FILLCELL_X1 FILLER_68_365 ();
 FILLCELL_X32 FILLER_68_373 ();
 FILLCELL_X8 FILLER_68_405 ();
 FILLCELL_X1 FILLER_68_413 ();
 FILLCELL_X16 FILLER_68_419 ();
 FILLCELL_X4 FILLER_68_435 ();
 FILLCELL_X4 FILLER_68_449 ();
 FILLCELL_X1 FILLER_68_453 ();
 FILLCELL_X4 FILLER_68_471 ();
 FILLCELL_X2 FILLER_68_475 ();
 FILLCELL_X1 FILLER_68_477 ();
 FILLCELL_X4 FILLER_68_490 ();
 FILLCELL_X8 FILLER_68_499 ();
 FILLCELL_X2 FILLER_68_507 ();
 FILLCELL_X1 FILLER_68_509 ();
 FILLCELL_X1 FILLER_68_514 ();
 FILLCELL_X4 FILLER_68_519 ();
 FILLCELL_X1 FILLER_68_559 ();
 FILLCELL_X8 FILLER_68_579 ();
 FILLCELL_X1 FILLER_68_587 ();
 FILLCELL_X2 FILLER_68_598 ();
 FILLCELL_X4 FILLER_68_626 ();
 FILLCELL_X1 FILLER_68_630 ();
 FILLCELL_X8 FILLER_68_632 ();
 FILLCELL_X4 FILLER_68_640 ();
 FILLCELL_X1 FILLER_68_644 ();
 FILLCELL_X1 FILLER_68_653 ();
 FILLCELL_X2 FILLER_68_671 ();
 FILLCELL_X4 FILLER_68_676 ();
 FILLCELL_X2 FILLER_68_680 ();
 FILLCELL_X1 FILLER_68_682 ();
 FILLCELL_X8 FILLER_68_695 ();
 FILLCELL_X4 FILLER_68_703 ();
 FILLCELL_X1 FILLER_68_707 ();
 FILLCELL_X4 FILLER_68_715 ();
 FILLCELL_X1 FILLER_68_719 ();
 FILLCELL_X16 FILLER_68_730 ();
 FILLCELL_X4 FILLER_68_746 ();
 FILLCELL_X2 FILLER_68_757 ();
 FILLCELL_X2 FILLER_68_776 ();
 FILLCELL_X1 FILLER_68_778 ();
 FILLCELL_X4 FILLER_68_788 ();
 FILLCELL_X2 FILLER_68_792 ();
 FILLCELL_X8 FILLER_68_801 ();
 FILLCELL_X4 FILLER_68_809 ();
 FILLCELL_X1 FILLER_68_813 ();
 FILLCELL_X16 FILLER_69_1 ();
 FILLCELL_X4 FILLER_69_17 ();
 FILLCELL_X2 FILLER_69_21 ();
 FILLCELL_X1 FILLER_69_47 ();
 FILLCELL_X2 FILLER_69_57 ();
 FILLCELL_X2 FILLER_69_64 ();
 FILLCELL_X4 FILLER_69_74 ();
 FILLCELL_X1 FILLER_69_85 ();
 FILLCELL_X4 FILLER_69_93 ();
 FILLCELL_X1 FILLER_69_97 ();
 FILLCELL_X4 FILLER_69_107 ();
 FILLCELL_X2 FILLER_69_111 ();
 FILLCELL_X16 FILLER_69_139 ();
 FILLCELL_X1 FILLER_69_155 ();
 FILLCELL_X1 FILLER_69_165 ();
 FILLCELL_X16 FILLER_69_175 ();
 FILLCELL_X1 FILLER_69_191 ();
 FILLCELL_X2 FILLER_69_201 ();
 FILLCELL_X1 FILLER_69_210 ();
 FILLCELL_X2 FILLER_69_215 ();
 FILLCELL_X1 FILLER_69_220 ();
 FILLCELL_X4 FILLER_69_252 ();
 FILLCELL_X2 FILLER_69_259 ();
 FILLCELL_X1 FILLER_69_261 ();
 FILLCELL_X8 FILLER_69_265 ();
 FILLCELL_X4 FILLER_69_287 ();
 FILLCELL_X1 FILLER_69_305 ();
 FILLCELL_X2 FILLER_69_330 ();
 FILLCELL_X8 FILLER_69_336 ();
 FILLCELL_X2 FILLER_69_344 ();
 FILLCELL_X2 FILLER_69_370 ();
 FILLCELL_X1 FILLER_69_372 ();
 FILLCELL_X16 FILLER_69_380 ();
 FILLCELL_X8 FILLER_69_396 ();
 FILLCELL_X4 FILLER_69_404 ();
 FILLCELL_X2 FILLER_69_408 ();
 FILLCELL_X1 FILLER_69_427 ();
 FILLCELL_X2 FILLER_69_445 ();
 FILLCELL_X2 FILLER_69_450 ();
 FILLCELL_X2 FILLER_69_455 ();
 FILLCELL_X2 FILLER_69_461 ();
 FILLCELL_X8 FILLER_69_466 ();
 FILLCELL_X4 FILLER_69_474 ();
 FILLCELL_X1 FILLER_69_478 ();
 FILLCELL_X16 FILLER_69_493 ();
 FILLCELL_X2 FILLER_69_509 ();
 FILLCELL_X1 FILLER_69_532 ();
 FILLCELL_X2 FILLER_69_546 ();
 FILLCELL_X2 FILLER_69_559 ();
 FILLCELL_X2 FILLER_69_566 ();
 FILLCELL_X1 FILLER_69_568 ();
 FILLCELL_X2 FILLER_69_578 ();
 FILLCELL_X2 FILLER_69_604 ();
 FILLCELL_X8 FILLER_69_617 ();
 FILLCELL_X4 FILLER_69_625 ();
 FILLCELL_X2 FILLER_69_629 ();
 FILLCELL_X1 FILLER_69_631 ();
 FILLCELL_X2 FILLER_69_665 ();
 FILLCELL_X2 FILLER_69_695 ();
 FILLCELL_X1 FILLER_69_701 ();
 FILLCELL_X1 FILLER_69_706 ();
 FILLCELL_X1 FILLER_69_716 ();
 FILLCELL_X2 FILLER_69_726 ();
 FILLCELL_X1 FILLER_69_732 ();
 FILLCELL_X2 FILLER_69_736 ();
 FILLCELL_X8 FILLER_69_741 ();
 FILLCELL_X1 FILLER_69_749 ();
 FILLCELL_X4 FILLER_69_762 ();
 FILLCELL_X1 FILLER_69_766 ();
 FILLCELL_X2 FILLER_69_774 ();
 FILLCELL_X16 FILLER_70_1 ();
 FILLCELL_X8 FILLER_70_17 ();
 FILLCELL_X4 FILLER_70_25 ();
 FILLCELL_X1 FILLER_70_32 ();
 FILLCELL_X8 FILLER_70_36 ();
 FILLCELL_X2 FILLER_70_44 ();
 FILLCELL_X4 FILLER_70_89 ();
 FILLCELL_X2 FILLER_70_93 ();
 FILLCELL_X4 FILLER_70_102 ();
 FILLCELL_X1 FILLER_70_106 ();
 FILLCELL_X2 FILLER_70_111 ();
 FILLCELL_X1 FILLER_70_116 ();
 FILLCELL_X16 FILLER_70_127 ();
 FILLCELL_X2 FILLER_70_150 ();
 FILLCELL_X1 FILLER_70_152 ();
 FILLCELL_X8 FILLER_70_167 ();
 FILLCELL_X2 FILLER_70_175 ();
 FILLCELL_X1 FILLER_70_177 ();
 FILLCELL_X1 FILLER_70_195 ();
 FILLCELL_X2 FILLER_70_203 ();
 FILLCELL_X2 FILLER_70_225 ();
 FILLCELL_X2 FILLER_70_230 ();
 FILLCELL_X8 FILLER_70_268 ();
 FILLCELL_X4 FILLER_70_281 ();
 FILLCELL_X2 FILLER_70_285 ();
 FILLCELL_X4 FILLER_70_294 ();
 FILLCELL_X1 FILLER_70_298 ();
 FILLCELL_X8 FILLER_70_313 ();
 FILLCELL_X1 FILLER_70_321 ();
 FILLCELL_X1 FILLER_70_327 ();
 FILLCELL_X8 FILLER_70_331 ();
 FILLCELL_X2 FILLER_70_339 ();
 FILLCELL_X8 FILLER_70_344 ();
 FILLCELL_X8 FILLER_70_383 ();
 FILLCELL_X2 FILLER_70_391 ();
 FILLCELL_X16 FILLER_70_400 ();
 FILLCELL_X2 FILLER_70_416 ();
 FILLCELL_X1 FILLER_70_418 ();
 FILLCELL_X4 FILLER_70_426 ();
 FILLCELL_X1 FILLER_70_430 ();
 FILLCELL_X1 FILLER_70_444 ();
 FILLCELL_X2 FILLER_70_449 ();
 FILLCELL_X2 FILLER_70_454 ();
 FILLCELL_X4 FILLER_70_460 ();
 FILLCELL_X2 FILLER_70_464 ();
 FILLCELL_X8 FILLER_70_469 ();
 FILLCELL_X4 FILLER_70_477 ();
 FILLCELL_X2 FILLER_70_481 ();
 FILLCELL_X1 FILLER_70_490 ();
 FILLCELL_X8 FILLER_70_496 ();
 FILLCELL_X2 FILLER_70_504 ();
 FILLCELL_X32 FILLER_70_520 ();
 FILLCELL_X8 FILLER_70_573 ();
 FILLCELL_X4 FILLER_70_581 ();
 FILLCELL_X2 FILLER_70_585 ();
 FILLCELL_X8 FILLER_70_603 ();
 FILLCELL_X2 FILLER_70_618 ();
 FILLCELL_X1 FILLER_70_630 ();
 FILLCELL_X4 FILLER_70_650 ();
 FILLCELL_X4 FILLER_70_661 ();
 FILLCELL_X2 FILLER_70_665 ();
 FILLCELL_X1 FILLER_70_667 ();
 FILLCELL_X4 FILLER_70_671 ();
 FILLCELL_X2 FILLER_70_675 ();
 FILLCELL_X8 FILLER_70_681 ();
 FILLCELL_X4 FILLER_70_689 ();
 FILLCELL_X1 FILLER_70_693 ();
 FILLCELL_X1 FILLER_70_699 ();
 FILLCELL_X1 FILLER_70_704 ();
 FILLCELL_X1 FILLER_70_715 ();
 FILLCELL_X8 FILLER_70_725 ();
 FILLCELL_X4 FILLER_70_753 ();
 FILLCELL_X4 FILLER_70_771 ();
 FILLCELL_X1 FILLER_70_775 ();
 FILLCELL_X2 FILLER_70_778 ();
 FILLCELL_X2 FILLER_70_783 ();
 FILLCELL_X2 FILLER_70_788 ();
 FILLCELL_X1 FILLER_70_790 ();
 FILLCELL_X8 FILLER_70_804 ();
 FILLCELL_X2 FILLER_70_812 ();
 FILLCELL_X4 FILLER_71_1 ();
 FILLCELL_X1 FILLER_71_5 ();
 FILLCELL_X16 FILLER_71_11 ();
 FILLCELL_X1 FILLER_71_27 ();
 FILLCELL_X1 FILLER_71_32 ();
 FILLCELL_X2 FILLER_71_38 ();
 FILLCELL_X1 FILLER_71_40 ();
 FILLCELL_X2 FILLER_71_58 ();
 FILLCELL_X1 FILLER_71_60 ();
 FILLCELL_X8 FILLER_71_65 ();
 FILLCELL_X2 FILLER_71_73 ();
 FILLCELL_X1 FILLER_71_75 ();
 FILLCELL_X2 FILLER_71_97 ();
 FILLCELL_X1 FILLER_71_135 ();
 FILLCELL_X1 FILLER_71_143 ();
 FILLCELL_X1 FILLER_71_161 ();
 FILLCELL_X8 FILLER_71_165 ();
 FILLCELL_X1 FILLER_71_194 ();
 FILLCELL_X2 FILLER_71_198 ();
 FILLCELL_X2 FILLER_71_203 ();
 FILLCELL_X32 FILLER_71_208 ();
 FILLCELL_X8 FILLER_71_254 ();
 FILLCELL_X2 FILLER_71_271 ();
 FILLCELL_X2 FILLER_71_276 ();
 FILLCELL_X1 FILLER_71_278 ();
 FILLCELL_X1 FILLER_71_286 ();
 FILLCELL_X4 FILLER_71_294 ();
 FILLCELL_X2 FILLER_71_305 ();
 FILLCELL_X1 FILLER_71_307 ();
 FILLCELL_X4 FILLER_71_318 ();
 FILLCELL_X1 FILLER_71_322 ();
 FILLCELL_X4 FILLER_71_347 ();
 FILLCELL_X2 FILLER_71_351 ();
 FILLCELL_X1 FILLER_71_353 ();
 FILLCELL_X1 FILLER_71_370 ();
 FILLCELL_X16 FILLER_71_388 ();
 FILLCELL_X8 FILLER_71_404 ();
 FILLCELL_X1 FILLER_71_412 ();
 FILLCELL_X4 FILLER_71_421 ();
 FILLCELL_X2 FILLER_71_450 ();
 FILLCELL_X1 FILLER_71_452 ();
 FILLCELL_X2 FILLER_71_477 ();
 FILLCELL_X2 FILLER_71_483 ();
 FILLCELL_X1 FILLER_71_485 ();
 FILLCELL_X8 FILLER_71_489 ();
 FILLCELL_X1 FILLER_71_497 ();
 FILLCELL_X2 FILLER_71_505 ();
 FILLCELL_X4 FILLER_71_529 ();
 FILLCELL_X1 FILLER_71_533 ();
 FILLCELL_X8 FILLER_71_540 ();
 FILLCELL_X4 FILLER_71_548 ();
 FILLCELL_X2 FILLER_71_552 ();
 FILLCELL_X2 FILLER_71_567 ();
 FILLCELL_X8 FILLER_71_573 ();
 FILLCELL_X4 FILLER_71_581 ();
 FILLCELL_X2 FILLER_71_585 ();
 FILLCELL_X2 FILLER_71_591 ();
 FILLCELL_X1 FILLER_71_593 ();
 FILLCELL_X8 FILLER_71_602 ();
 FILLCELL_X4 FILLER_71_610 ();
 FILLCELL_X1 FILLER_71_614 ();
 FILLCELL_X4 FILLER_71_641 ();
 FILLCELL_X2 FILLER_71_645 ();
 FILLCELL_X2 FILLER_71_664 ();
 FILLCELL_X2 FILLER_71_720 ();
 FILLCELL_X1 FILLER_71_722 ();
 FILLCELL_X1 FILLER_71_730 ();
 FILLCELL_X2 FILLER_71_743 ();
 FILLCELL_X2 FILLER_71_749 ();
 FILLCELL_X1 FILLER_71_768 ();
 FILLCELL_X1 FILLER_71_772 ();
 FILLCELL_X2 FILLER_71_795 ();
 FILLCELL_X8 FILLER_72_1 ();
 FILLCELL_X4 FILLER_72_9 ();
 FILLCELL_X2 FILLER_72_13 ();
 FILLCELL_X4 FILLER_72_35 ();
 FILLCELL_X4 FILLER_72_42 ();
 FILLCELL_X2 FILLER_72_46 ();
 FILLCELL_X1 FILLER_72_48 ();
 FILLCELL_X4 FILLER_72_52 ();
 FILLCELL_X2 FILLER_72_56 ();
 FILLCELL_X4 FILLER_72_62 ();
 FILLCELL_X2 FILLER_72_66 ();
 FILLCELL_X1 FILLER_72_68 ();
 FILLCELL_X1 FILLER_72_73 ();
 FILLCELL_X32 FILLER_72_81 ();
 FILLCELL_X2 FILLER_72_113 ();
 FILLCELL_X4 FILLER_72_122 ();
 FILLCELL_X2 FILLER_72_126 ();
 FILLCELL_X1 FILLER_72_128 ();
 FILLCELL_X2 FILLER_72_141 ();
 FILLCELL_X16 FILLER_72_164 ();
 FILLCELL_X8 FILLER_72_180 ();
 FILLCELL_X8 FILLER_72_191 ();
 FILLCELL_X1 FILLER_72_202 ();
 FILLCELL_X4 FILLER_72_208 ();
 FILLCELL_X2 FILLER_72_212 ();
 FILLCELL_X2 FILLER_72_222 ();
 FILLCELL_X1 FILLER_72_224 ();
 FILLCELL_X4 FILLER_72_230 ();
 FILLCELL_X1 FILLER_72_234 ();
 FILLCELL_X1 FILLER_72_255 ();
 FILLCELL_X2 FILLER_72_276 ();
 FILLCELL_X2 FILLER_72_302 ();
 FILLCELL_X16 FILLER_72_326 ();
 FILLCELL_X1 FILLER_72_342 ();
 FILLCELL_X2 FILLER_72_360 ();
 FILLCELL_X1 FILLER_72_367 ();
 FILLCELL_X16 FILLER_72_375 ();
 FILLCELL_X8 FILLER_72_391 ();
 FILLCELL_X2 FILLER_72_399 ();
 FILLCELL_X1 FILLER_72_401 ();
 FILLCELL_X16 FILLER_72_422 ();
 FILLCELL_X4 FILLER_72_438 ();
 FILLCELL_X1 FILLER_72_442 ();
 FILLCELL_X1 FILLER_72_464 ();
 FILLCELL_X1 FILLER_72_493 ();
 FILLCELL_X1 FILLER_72_497 ();
 FILLCELL_X1 FILLER_72_508 ();
 FILLCELL_X2 FILLER_72_524 ();
 FILLCELL_X1 FILLER_72_526 ();
 FILLCELL_X8 FILLER_72_532 ();
 FILLCELL_X2 FILLER_72_540 ();
 FILLCELL_X1 FILLER_72_542 ();
 FILLCELL_X2 FILLER_72_547 ();
 FILLCELL_X1 FILLER_72_549 ();
 FILLCELL_X8 FILLER_72_564 ();
 FILLCELL_X1 FILLER_72_572 ();
 FILLCELL_X4 FILLER_72_618 ();
 FILLCELL_X2 FILLER_72_622 ();
 FILLCELL_X16 FILLER_72_632 ();
 FILLCELL_X2 FILLER_72_648 ();
 FILLCELL_X8 FILLER_72_658 ();
 FILLCELL_X4 FILLER_72_666 ();
 FILLCELL_X2 FILLER_72_677 ();
 FILLCELL_X1 FILLER_72_679 ();
 FILLCELL_X1 FILLER_72_684 ();
 FILLCELL_X2 FILLER_72_692 ();
 FILLCELL_X16 FILLER_72_702 ();
 FILLCELL_X8 FILLER_72_718 ();
 FILLCELL_X4 FILLER_72_726 ();
 FILLCELL_X1 FILLER_72_730 ();
 FILLCELL_X4 FILLER_72_734 ();
 FILLCELL_X16 FILLER_72_742 ();
 FILLCELL_X8 FILLER_72_758 ();
 FILLCELL_X4 FILLER_72_766 ();
 FILLCELL_X2 FILLER_72_770 ();
 FILLCELL_X4 FILLER_72_774 ();
 FILLCELL_X1 FILLER_72_778 ();
 FILLCELL_X4 FILLER_72_782 ();
 FILLCELL_X2 FILLER_72_786 ();
 FILLCELL_X1 FILLER_72_788 ();
 FILLCELL_X4 FILLER_72_796 ();
 FILLCELL_X1 FILLER_72_800 ();
 FILLCELL_X8 FILLER_72_804 ();
 FILLCELL_X2 FILLER_72_812 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X1 FILLER_73_33 ();
 FILLCELL_X2 FILLER_73_37 ();
 FILLCELL_X2 FILLER_73_69 ();
 FILLCELL_X16 FILLER_73_82 ();
 FILLCELL_X2 FILLER_73_98 ();
 FILLCELL_X1 FILLER_73_100 ();
 FILLCELL_X1 FILLER_73_112 ();
 FILLCELL_X4 FILLER_73_120 ();
 FILLCELL_X2 FILLER_73_124 ();
 FILLCELL_X8 FILLER_73_148 ();
 FILLCELL_X16 FILLER_73_161 ();
 FILLCELL_X4 FILLER_73_177 ();
 FILLCELL_X2 FILLER_73_181 ();
 FILLCELL_X4 FILLER_73_190 ();
 FILLCELL_X2 FILLER_73_201 ();
 FILLCELL_X2 FILLER_73_216 ();
 FILLCELL_X8 FILLER_73_222 ();
 FILLCELL_X16 FILLER_73_233 ();
 FILLCELL_X32 FILLER_73_256 ();
 FILLCELL_X2 FILLER_73_293 ();
 FILLCELL_X4 FILLER_73_298 ();
 FILLCELL_X1 FILLER_73_302 ();
 FILLCELL_X16 FILLER_73_311 ();
 FILLCELL_X1 FILLER_73_327 ();
 FILLCELL_X8 FILLER_73_338 ();
 FILLCELL_X2 FILLER_73_346 ();
 FILLCELL_X4 FILLER_73_355 ();
 FILLCELL_X1 FILLER_73_359 ();
 FILLCELL_X1 FILLER_73_363 ();
 FILLCELL_X4 FILLER_73_367 ();
 FILLCELL_X1 FILLER_73_371 ();
 FILLCELL_X4 FILLER_73_386 ();
 FILLCELL_X2 FILLER_73_390 ();
 FILLCELL_X1 FILLER_73_392 ();
 FILLCELL_X1 FILLER_73_400 ();
 FILLCELL_X1 FILLER_73_408 ();
 FILLCELL_X8 FILLER_73_416 ();
 FILLCELL_X16 FILLER_73_454 ();
 FILLCELL_X8 FILLER_73_470 ();
 FILLCELL_X2 FILLER_73_478 ();
 FILLCELL_X2 FILLER_73_483 ();
 FILLCELL_X8 FILLER_73_502 ();
 FILLCELL_X4 FILLER_73_510 ();
 FILLCELL_X1 FILLER_73_525 ();
 FILLCELL_X2 FILLER_73_531 ();
 FILLCELL_X1 FILLER_73_533 ();
 FILLCELL_X32 FILLER_73_599 ();
 FILLCELL_X8 FILLER_73_631 ();
 FILLCELL_X4 FILLER_73_639 ();
 FILLCELL_X2 FILLER_73_643 ();
 FILLCELL_X4 FILLER_73_652 ();
 FILLCELL_X1 FILLER_73_656 ();
 FILLCELL_X2 FILLER_73_694 ();
 FILLCELL_X1 FILLER_73_701 ();
 FILLCELL_X4 FILLER_73_719 ();
 FILLCELL_X2 FILLER_73_723 ();
 FILLCELL_X2 FILLER_73_745 ();
 FILLCELL_X2 FILLER_73_750 ();
 FILLCELL_X8 FILLER_73_759 ();
 FILLCELL_X4 FILLER_73_774 ();
 FILLCELL_X2 FILLER_73_778 ();
 FILLCELL_X1 FILLER_73_780 ();
 FILLCELL_X2 FILLER_73_798 ();
 FILLCELL_X8 FILLER_73_804 ();
 FILLCELL_X2 FILLER_73_812 ();
 FILLCELL_X16 FILLER_74_1 ();
 FILLCELL_X8 FILLER_74_17 ();
 FILLCELL_X4 FILLER_74_25 ();
 FILLCELL_X8 FILLER_74_34 ();
 FILLCELL_X1 FILLER_74_42 ();
 FILLCELL_X4 FILLER_74_46 ();
 FILLCELL_X2 FILLER_74_50 ();
 FILLCELL_X1 FILLER_74_52 ();
 FILLCELL_X4 FILLER_74_58 ();
 FILLCELL_X8 FILLER_74_79 ();
 FILLCELL_X1 FILLER_74_87 ();
 FILLCELL_X1 FILLER_74_105 ();
 FILLCELL_X2 FILLER_74_113 ();
 FILLCELL_X1 FILLER_74_115 ();
 FILLCELL_X4 FILLER_74_123 ();
 FILLCELL_X8 FILLER_74_132 ();
 FILLCELL_X4 FILLER_74_140 ();
 FILLCELL_X2 FILLER_74_144 ();
 FILLCELL_X8 FILLER_74_151 ();
 FILLCELL_X1 FILLER_74_162 ();
 FILLCELL_X4 FILLER_74_180 ();
 FILLCELL_X2 FILLER_74_207 ();
 FILLCELL_X1 FILLER_74_209 ();
 FILLCELL_X2 FILLER_74_234 ();
 FILLCELL_X1 FILLER_74_236 ();
 FILLCELL_X4 FILLER_74_240 ();
 FILLCELL_X2 FILLER_74_244 ();
 FILLCELL_X1 FILLER_74_246 ();
 FILLCELL_X4 FILLER_74_250 ();
 FILLCELL_X1 FILLER_74_254 ();
 FILLCELL_X2 FILLER_74_262 ();
 FILLCELL_X1 FILLER_74_264 ();
 FILLCELL_X8 FILLER_74_278 ();
 FILLCELL_X8 FILLER_74_306 ();
 FILLCELL_X1 FILLER_74_314 ();
 FILLCELL_X16 FILLER_74_322 ();
 FILLCELL_X1 FILLER_74_365 ();
 FILLCELL_X8 FILLER_74_390 ();
 FILLCELL_X4 FILLER_74_405 ();
 FILLCELL_X2 FILLER_74_409 ();
 FILLCELL_X4 FILLER_74_418 ();
 FILLCELL_X8 FILLER_74_425 ();
 FILLCELL_X4 FILLER_74_433 ();
 FILLCELL_X2 FILLER_74_447 ();
 FILLCELL_X8 FILLER_74_455 ();
 FILLCELL_X4 FILLER_74_463 ();
 FILLCELL_X2 FILLER_74_467 ();
 FILLCELL_X8 FILLER_74_476 ();
 FILLCELL_X8 FILLER_74_492 ();
 FILLCELL_X4 FILLER_74_500 ();
 FILLCELL_X1 FILLER_74_504 ();
 FILLCELL_X2 FILLER_74_508 ();
 FILLCELL_X2 FILLER_74_517 ();
 FILLCELL_X1 FILLER_74_530 ();
 FILLCELL_X2 FILLER_74_540 ();
 FILLCELL_X1 FILLER_74_542 ();
 FILLCELL_X2 FILLER_74_548 ();
 FILLCELL_X8 FILLER_74_552 ();
 FILLCELL_X2 FILLER_74_560 ();
 FILLCELL_X8 FILLER_74_567 ();
 FILLCELL_X4 FILLER_74_575 ();
 FILLCELL_X1 FILLER_74_579 ();
 FILLCELL_X2 FILLER_74_585 ();
 FILLCELL_X2 FILLER_74_591 ();
 FILLCELL_X2 FILLER_74_604 ();
 FILLCELL_X2 FILLER_74_627 ();
 FILLCELL_X4 FILLER_74_646 ();
 FILLCELL_X1 FILLER_74_650 ();
 FILLCELL_X4 FILLER_74_668 ();
 FILLCELL_X1 FILLER_74_672 ();
 FILLCELL_X8 FILLER_74_678 ();
 FILLCELL_X4 FILLER_74_686 ();
 FILLCELL_X2 FILLER_74_690 ();
 FILLCELL_X2 FILLER_74_709 ();
 FILLCELL_X1 FILLER_74_711 ();
 FILLCELL_X8 FILLER_74_715 ();
 FILLCELL_X4 FILLER_74_723 ();
 FILLCELL_X2 FILLER_74_727 ();
 FILLCELL_X1 FILLER_74_729 ();
 FILLCELL_X8 FILLER_74_737 ();
 FILLCELL_X4 FILLER_74_745 ();
 FILLCELL_X2 FILLER_74_749 ();
 FILLCELL_X1 FILLER_74_751 ();
 FILLCELL_X4 FILLER_74_764 ();
 FILLCELL_X2 FILLER_74_768 ();
 FILLCELL_X1 FILLER_74_770 ();
 FILLCELL_X8 FILLER_74_778 ();
 FILLCELL_X2 FILLER_74_786 ();
 FILLCELL_X1 FILLER_74_788 ();
 FILLCELL_X8 FILLER_74_799 ();
 FILLCELL_X4 FILLER_74_807 ();
 FILLCELL_X2 FILLER_74_811 ();
 FILLCELL_X1 FILLER_74_813 ();
 FILLCELL_X16 FILLER_75_1 ();
 FILLCELL_X4 FILLER_75_17 ();
 FILLCELL_X2 FILLER_75_21 ();
 FILLCELL_X1 FILLER_75_23 ();
 FILLCELL_X1 FILLER_75_45 ();
 FILLCELL_X4 FILLER_75_57 ();
 FILLCELL_X2 FILLER_75_61 ();
 FILLCELL_X4 FILLER_75_98 ();
 FILLCELL_X1 FILLER_75_102 ();
 FILLCELL_X16 FILLER_75_117 ();
 FILLCELL_X8 FILLER_75_133 ();
 FILLCELL_X4 FILLER_75_141 ();
 FILLCELL_X2 FILLER_75_145 ();
 FILLCELL_X1 FILLER_75_147 ();
 FILLCELL_X4 FILLER_75_153 ();
 FILLCELL_X2 FILLER_75_161 ();
 FILLCELL_X2 FILLER_75_173 ();
 FILLCELL_X1 FILLER_75_175 ();
 FILLCELL_X16 FILLER_75_200 ();
 FILLCELL_X4 FILLER_75_238 ();
 FILLCELL_X2 FILLER_75_273 ();
 FILLCELL_X4 FILLER_75_278 ();
 FILLCELL_X2 FILLER_75_310 ();
 FILLCELL_X8 FILLER_75_322 ();
 FILLCELL_X1 FILLER_75_343 ();
 FILLCELL_X1 FILLER_75_353 ();
 FILLCELL_X4 FILLER_75_371 ();
 FILLCELL_X2 FILLER_75_375 ();
 FILLCELL_X1 FILLER_75_384 ();
 FILLCELL_X8 FILLER_75_399 ();
 FILLCELL_X1 FILLER_75_407 ();
 FILLCELL_X1 FILLER_75_425 ();
 FILLCELL_X1 FILLER_75_431 ();
 FILLCELL_X2 FILLER_75_444 ();
 FILLCELL_X1 FILLER_75_467 ();
 FILLCELL_X16 FILLER_75_475 ();
 FILLCELL_X4 FILLER_75_491 ();
 FILLCELL_X1 FILLER_75_495 ();
 FILLCELL_X2 FILLER_75_503 ();
 FILLCELL_X2 FILLER_75_522 ();
 FILLCELL_X4 FILLER_75_547 ();
 FILLCELL_X4 FILLER_75_558 ();
 FILLCELL_X2 FILLER_75_562 ();
 FILLCELL_X1 FILLER_75_564 ();
 FILLCELL_X4 FILLER_75_574 ();
 FILLCELL_X1 FILLER_75_583 ();
 FILLCELL_X2 FILLER_75_591 ();
 FILLCELL_X1 FILLER_75_607 ();
 FILLCELL_X2 FILLER_75_647 ();
 FILLCELL_X1 FILLER_75_649 ();
 FILLCELL_X1 FILLER_75_665 ();
 FILLCELL_X8 FILLER_75_673 ();
 FILLCELL_X4 FILLER_75_708 ();
 FILLCELL_X2 FILLER_75_721 ();
 FILLCELL_X1 FILLER_75_723 ();
 FILLCELL_X1 FILLER_75_727 ();
 FILLCELL_X4 FILLER_75_760 ();
 FILLCELL_X2 FILLER_75_764 ();
 FILLCELL_X4 FILLER_75_769 ();
 FILLCELL_X2 FILLER_75_773 ();
 FILLCELL_X1 FILLER_75_775 ();
 FILLCELL_X2 FILLER_75_793 ();
 FILLCELL_X1 FILLER_75_795 ();
 FILLCELL_X8 FILLER_75_801 ();
 FILLCELL_X4 FILLER_75_809 ();
 FILLCELL_X1 FILLER_75_813 ();
 FILLCELL_X16 FILLER_76_1 ();
 FILLCELL_X8 FILLER_76_17 ();
 FILLCELL_X2 FILLER_76_30 ();
 FILLCELL_X1 FILLER_76_42 ();
 FILLCELL_X8 FILLER_76_67 ();
 FILLCELL_X1 FILLER_76_75 ();
 FILLCELL_X1 FILLER_76_92 ();
 FILLCELL_X1 FILLER_76_97 ();
 FILLCELL_X16 FILLER_76_102 ();
 FILLCELL_X4 FILLER_76_118 ();
 FILLCELL_X2 FILLER_76_148 ();
 FILLCELL_X1 FILLER_76_150 ();
 FILLCELL_X16 FILLER_76_168 ();
 FILLCELL_X8 FILLER_76_184 ();
 FILLCELL_X2 FILLER_76_192 ();
 FILLCELL_X1 FILLER_76_194 ();
 FILLCELL_X16 FILLER_76_212 ();
 FILLCELL_X4 FILLER_76_228 ();
 FILLCELL_X2 FILLER_76_232 ();
 FILLCELL_X1 FILLER_76_234 ();
 FILLCELL_X4 FILLER_76_252 ();
 FILLCELL_X2 FILLER_76_256 ();
 FILLCELL_X2 FILLER_76_263 ();
 FILLCELL_X4 FILLER_76_282 ();
 FILLCELL_X1 FILLER_76_303 ();
 FILLCELL_X8 FILLER_76_321 ();
 FILLCELL_X2 FILLER_76_353 ();
 FILLCELL_X8 FILLER_76_360 ();
 FILLCELL_X4 FILLER_76_368 ();
 FILLCELL_X1 FILLER_76_376 ();
 FILLCELL_X4 FILLER_76_391 ();
 FILLCELL_X2 FILLER_76_395 ();
 FILLCELL_X1 FILLER_76_397 ();
 FILLCELL_X4 FILLER_76_405 ();
 FILLCELL_X2 FILLER_76_412 ();
 FILLCELL_X1 FILLER_76_414 ();
 FILLCELL_X4 FILLER_76_420 ();
 FILLCELL_X2 FILLER_76_424 ();
 FILLCELL_X4 FILLER_76_429 ();
 FILLCELL_X1 FILLER_76_433 ();
 FILLCELL_X2 FILLER_76_438 ();
 FILLCELL_X1 FILLER_76_440 ();
 FILLCELL_X4 FILLER_76_444 ();
 FILLCELL_X2 FILLER_76_448 ();
 FILLCELL_X1 FILLER_76_450 ();
 FILLCELL_X2 FILLER_76_459 ();
 FILLCELL_X1 FILLER_76_461 ();
 FILLCELL_X8 FILLER_76_469 ();
 FILLCELL_X4 FILLER_76_477 ();
 FILLCELL_X1 FILLER_76_481 ();
 FILLCELL_X8 FILLER_76_507 ();
 FILLCELL_X2 FILLER_76_515 ();
 FILLCELL_X8 FILLER_76_533 ();
 FILLCELL_X4 FILLER_76_541 ();
 FILLCELL_X2 FILLER_76_545 ();
 FILLCELL_X1 FILLER_76_547 ();
 FILLCELL_X2 FILLER_76_563 ();
 FILLCELL_X4 FILLER_76_606 ();
 FILLCELL_X4 FILLER_76_620 ();
 FILLCELL_X2 FILLER_76_624 ();
 FILLCELL_X2 FILLER_76_628 ();
 FILLCELL_X1 FILLER_76_630 ();
 FILLCELL_X4 FILLER_76_639 ();
 FILLCELL_X2 FILLER_76_643 ();
 FILLCELL_X8 FILLER_76_647 ();
 FILLCELL_X1 FILLER_76_655 ();
 FILLCELL_X16 FILLER_76_661 ();
 FILLCELL_X2 FILLER_76_677 ();
 FILLCELL_X2 FILLER_76_683 ();
 FILLCELL_X1 FILLER_76_697 ();
 FILLCELL_X4 FILLER_76_702 ();
 FILLCELL_X8 FILLER_76_713 ();
 FILLCELL_X2 FILLER_76_721 ();
 FILLCELL_X1 FILLER_76_723 ();
 FILLCELL_X8 FILLER_76_741 ();
 FILLCELL_X16 FILLER_76_795 ();
 FILLCELL_X2 FILLER_76_811 ();
 FILLCELL_X1 FILLER_76_813 ();
 FILLCELL_X16 FILLER_77_1 ();
 FILLCELL_X2 FILLER_77_17 ();
 FILLCELL_X1 FILLER_77_19 ();
 FILLCELL_X2 FILLER_77_42 ();
 FILLCELL_X1 FILLER_77_44 ();
 FILLCELL_X8 FILLER_77_55 ();
 FILLCELL_X4 FILLER_77_63 ();
 FILLCELL_X2 FILLER_77_67 ();
 FILLCELL_X8 FILLER_77_74 ();
 FILLCELL_X1 FILLER_77_82 ();
 FILLCELL_X1 FILLER_77_87 ();
 FILLCELL_X4 FILLER_77_112 ();
 FILLCELL_X2 FILLER_77_116 ();
 FILLCELL_X1 FILLER_77_118 ();
 FILLCELL_X8 FILLER_77_124 ();
 FILLCELL_X4 FILLER_77_132 ();
 FILLCELL_X8 FILLER_77_143 ();
 FILLCELL_X2 FILLER_77_151 ();
 FILLCELL_X1 FILLER_77_157 ();
 FILLCELL_X1 FILLER_77_162 ();
 FILLCELL_X4 FILLER_77_184 ();
 FILLCELL_X1 FILLER_77_188 ();
 FILLCELL_X2 FILLER_77_199 ();
 FILLCELL_X4 FILLER_77_212 ();
 FILLCELL_X2 FILLER_77_216 ();
 FILLCELL_X1 FILLER_77_218 ();
 FILLCELL_X4 FILLER_77_226 ();
 FILLCELL_X8 FILLER_77_233 ();
 FILLCELL_X4 FILLER_77_241 ();
 FILLCELL_X2 FILLER_77_245 ();
 FILLCELL_X1 FILLER_77_247 ();
 FILLCELL_X1 FILLER_77_253 ();
 FILLCELL_X8 FILLER_77_259 ();
 FILLCELL_X16 FILLER_77_270 ();
 FILLCELL_X8 FILLER_77_286 ();
 FILLCELL_X2 FILLER_77_294 ();
 FILLCELL_X1 FILLER_77_296 ();
 FILLCELL_X1 FILLER_77_300 ();
 FILLCELL_X16 FILLER_77_304 ();
 FILLCELL_X4 FILLER_77_320 ();
 FILLCELL_X8 FILLER_77_331 ();
 FILLCELL_X2 FILLER_77_339 ();
 FILLCELL_X1 FILLER_77_341 ();
 FILLCELL_X2 FILLER_77_349 ();
 FILLCELL_X4 FILLER_77_358 ();
 FILLCELL_X2 FILLER_77_362 ();
 FILLCELL_X1 FILLER_77_364 ();
 FILLCELL_X4 FILLER_77_392 ();
 FILLCELL_X1 FILLER_77_396 ();
 FILLCELL_X8 FILLER_77_404 ();
 FILLCELL_X2 FILLER_77_416 ();
 FILLCELL_X1 FILLER_77_418 ();
 FILLCELL_X8 FILLER_77_422 ();
 FILLCELL_X1 FILLER_77_450 ();
 FILLCELL_X4 FILLER_77_454 ();
 FILLCELL_X2 FILLER_77_458 ();
 FILLCELL_X4 FILLER_77_482 ();
 FILLCELL_X1 FILLER_77_486 ();
 FILLCELL_X1 FILLER_77_491 ();
 FILLCELL_X2 FILLER_77_495 ();
 FILLCELL_X1 FILLER_77_497 ();
 FILLCELL_X8 FILLER_77_505 ();
 FILLCELL_X1 FILLER_77_513 ();
 FILLCELL_X2 FILLER_77_518 ();
 FILLCELL_X1 FILLER_77_520 ();
 FILLCELL_X16 FILLER_77_525 ();
 FILLCELL_X4 FILLER_77_541 ();
 FILLCELL_X1 FILLER_77_545 ();
 FILLCELL_X2 FILLER_77_576 ();
 FILLCELL_X4 FILLER_77_583 ();
 FILLCELL_X1 FILLER_77_587 ();
 FILLCELL_X1 FILLER_77_592 ();
 FILLCELL_X4 FILLER_77_607 ();
 FILLCELL_X16 FILLER_77_619 ();
 FILLCELL_X8 FILLER_77_635 ();
 FILLCELL_X2 FILLER_77_653 ();
 FILLCELL_X8 FILLER_77_663 ();
 FILLCELL_X4 FILLER_77_671 ();
 FILLCELL_X2 FILLER_77_675 ();
 FILLCELL_X1 FILLER_77_677 ();
 FILLCELL_X2 FILLER_77_695 ();
 FILLCELL_X1 FILLER_77_697 ();
 FILLCELL_X2 FILLER_77_705 ();
 FILLCELL_X1 FILLER_77_707 ();
 FILLCELL_X4 FILLER_77_715 ();
 FILLCELL_X2 FILLER_77_719 ();
 FILLCELL_X1 FILLER_77_721 ();
 FILLCELL_X4 FILLER_77_737 ();
 FILLCELL_X1 FILLER_77_741 ();
 FILLCELL_X2 FILLER_77_747 ();
 FILLCELL_X1 FILLER_77_749 ();
 FILLCELL_X2 FILLER_77_777 ();
 FILLCELL_X16 FILLER_77_787 ();
 FILLCELL_X8 FILLER_77_803 ();
 FILLCELL_X2 FILLER_77_811 ();
 FILLCELL_X1 FILLER_77_813 ();
 FILLCELL_X16 FILLER_78_1 ();
 FILLCELL_X8 FILLER_78_17 ();
 FILLCELL_X1 FILLER_78_25 ();
 FILLCELL_X4 FILLER_78_33 ();
 FILLCELL_X2 FILLER_78_37 ();
 FILLCELL_X1 FILLER_78_39 ();
 FILLCELL_X8 FILLER_78_57 ();
 FILLCELL_X4 FILLER_78_65 ();
 FILLCELL_X1 FILLER_78_86 ();
 FILLCELL_X8 FILLER_78_108 ();
 FILLCELL_X4 FILLER_78_116 ();
 FILLCELL_X2 FILLER_78_120 ();
 FILLCELL_X1 FILLER_78_122 ();
 FILLCELL_X1 FILLER_78_147 ();
 FILLCELL_X4 FILLER_78_179 ();
 FILLCELL_X1 FILLER_78_183 ();
 FILLCELL_X2 FILLER_78_201 ();
 FILLCELL_X1 FILLER_78_203 ();
 FILLCELL_X8 FILLER_78_208 ();
 FILLCELL_X1 FILLER_78_216 ();
 FILLCELL_X4 FILLER_78_234 ();
 FILLCELL_X1 FILLER_78_242 ();
 FILLCELL_X4 FILLER_78_277 ();
 FILLCELL_X4 FILLER_78_288 ();
 FILLCELL_X2 FILLER_78_292 ();
 FILLCELL_X1 FILLER_78_294 ();
 FILLCELL_X4 FILLER_78_305 ();
 FILLCELL_X2 FILLER_78_316 ();
 FILLCELL_X16 FILLER_78_335 ();
 FILLCELL_X2 FILLER_78_351 ();
 FILLCELL_X1 FILLER_78_353 ();
 FILLCELL_X16 FILLER_78_357 ();
 FILLCELL_X8 FILLER_78_373 ();
 FILLCELL_X1 FILLER_78_381 ();
 FILLCELL_X16 FILLER_78_385 ();
 FILLCELL_X4 FILLER_78_401 ();
 FILLCELL_X1 FILLER_78_405 ();
 FILLCELL_X4 FILLER_78_423 ();
 FILLCELL_X1 FILLER_78_427 ();
 FILLCELL_X1 FILLER_78_440 ();
 FILLCELL_X2 FILLER_78_458 ();
 FILLCELL_X1 FILLER_78_460 ();
 FILLCELL_X2 FILLER_78_464 ();
 FILLCELL_X8 FILLER_78_480 ();
 FILLCELL_X8 FILLER_78_498 ();
 FILLCELL_X1 FILLER_78_523 ();
 FILLCELL_X1 FILLER_78_538 ();
 FILLCELL_X4 FILLER_78_563 ();
 FILLCELL_X8 FILLER_78_574 ();
 FILLCELL_X4 FILLER_78_582 ();
 FILLCELL_X8 FILLER_78_595 ();
 FILLCELL_X1 FILLER_78_603 ();
 FILLCELL_X8 FILLER_78_677 ();
 FILLCELL_X1 FILLER_78_685 ();
 FILLCELL_X1 FILLER_78_691 ();
 FILLCELL_X1 FILLER_78_700 ();
 FILLCELL_X2 FILLER_78_718 ();
 FILLCELL_X4 FILLER_78_724 ();
 FILLCELL_X2 FILLER_78_728 ();
 FILLCELL_X1 FILLER_78_730 ();
 FILLCELL_X1 FILLER_78_734 ();
 FILLCELL_X2 FILLER_78_744 ();
 FILLCELL_X1 FILLER_78_746 ();
 FILLCELL_X8 FILLER_78_763 ();
 FILLCELL_X4 FILLER_78_771 ();
 FILLCELL_X2 FILLER_78_775 ();
 FILLCELL_X1 FILLER_78_777 ();
 FILLCELL_X8 FILLER_78_802 ();
 FILLCELL_X4 FILLER_78_810 ();
 FILLCELL_X16 FILLER_79_1 ();
 FILLCELL_X4 FILLER_79_17 ();
 FILLCELL_X1 FILLER_79_21 ();
 FILLCELL_X16 FILLER_79_27 ();
 FILLCELL_X4 FILLER_79_43 ();
 FILLCELL_X4 FILLER_79_50 ();
 FILLCELL_X2 FILLER_79_54 ();
 FILLCELL_X4 FILLER_79_73 ();
 FILLCELL_X2 FILLER_79_77 ();
 FILLCELL_X1 FILLER_79_79 ();
 FILLCELL_X2 FILLER_79_84 ();
 FILLCELL_X16 FILLER_79_93 ();
 FILLCELL_X16 FILLER_79_116 ();
 FILLCELL_X4 FILLER_79_132 ();
 FILLCELL_X2 FILLER_79_136 ();
 FILLCELL_X4 FILLER_79_145 ();
 FILLCELL_X1 FILLER_79_149 ();
 FILLCELL_X8 FILLER_79_157 ();
 FILLCELL_X4 FILLER_79_165 ();
 FILLCELL_X16 FILLER_79_183 ();
 FILLCELL_X8 FILLER_79_215 ();
 FILLCELL_X2 FILLER_79_223 ();
 FILLCELL_X1 FILLER_79_225 ();
 FILLCELL_X2 FILLER_79_250 ();
 FILLCELL_X4 FILLER_79_266 ();
 FILLCELL_X2 FILLER_79_290 ();
 FILLCELL_X4 FILLER_79_309 ();
 FILLCELL_X2 FILLER_79_313 ();
 FILLCELL_X1 FILLER_79_329 ();
 FILLCELL_X2 FILLER_79_344 ();
 FILLCELL_X1 FILLER_79_346 ();
 FILLCELL_X2 FILLER_79_371 ();
 FILLCELL_X1 FILLER_79_373 ();
 FILLCELL_X4 FILLER_79_381 ();
 FILLCELL_X4 FILLER_79_395 ();
 FILLCELL_X2 FILLER_79_399 ();
 FILLCELL_X1 FILLER_79_401 ();
 FILLCELL_X2 FILLER_79_444 ();
 FILLCELL_X2 FILLER_79_463 ();
 FILLCELL_X1 FILLER_79_465 ();
 FILLCELL_X8 FILLER_79_473 ();
 FILLCELL_X2 FILLER_79_481 ();
 FILLCELL_X1 FILLER_79_514 ();
 FILLCELL_X2 FILLER_79_518 ();
 FILLCELL_X1 FILLER_79_520 ();
 FILLCELL_X1 FILLER_79_529 ();
 FILLCELL_X2 FILLER_79_533 ();
 FILLCELL_X2 FILLER_79_555 ();
 FILLCELL_X4 FILLER_79_561 ();
 FILLCELL_X2 FILLER_79_565 ();
 FILLCELL_X4 FILLER_79_574 ();
 FILLCELL_X2 FILLER_79_578 ();
 FILLCELL_X8 FILLER_79_597 ();
 FILLCELL_X4 FILLER_79_605 ();
 FILLCELL_X2 FILLER_79_609 ();
 FILLCELL_X2 FILLER_79_616 ();
 FILLCELL_X4 FILLER_79_637 ();
 FILLCELL_X2 FILLER_79_641 ();
 FILLCELL_X1 FILLER_79_643 ();
 FILLCELL_X2 FILLER_79_647 ();
 FILLCELL_X1 FILLER_79_649 ();
 FILLCELL_X2 FILLER_79_653 ();
 FILLCELL_X1 FILLER_79_655 ();
 FILLCELL_X4 FILLER_79_670 ();
 FILLCELL_X8 FILLER_79_679 ();
 FILLCELL_X1 FILLER_79_687 ();
 FILLCELL_X8 FILLER_79_713 ();
 FILLCELL_X2 FILLER_79_721 ();
 FILLCELL_X2 FILLER_79_747 ();
 FILLCELL_X1 FILLER_79_749 ();
 FILLCELL_X4 FILLER_79_757 ();
 FILLCELL_X4 FILLER_79_778 ();
 FILLCELL_X4 FILLER_79_785 ();
 FILLCELL_X2 FILLER_79_789 ();
 FILLCELL_X4 FILLER_79_808 ();
 FILLCELL_X2 FILLER_79_812 ();
 FILLCELL_X16 FILLER_80_1 ();
 FILLCELL_X8 FILLER_80_17 ();
 FILLCELL_X4 FILLER_80_25 ();
 FILLCELL_X1 FILLER_80_29 ();
 FILLCELL_X4 FILLER_80_37 ();
 FILLCELL_X1 FILLER_80_48 ();
 FILLCELL_X4 FILLER_80_56 ();
 FILLCELL_X2 FILLER_80_60 ();
 FILLCELL_X1 FILLER_80_62 ();
 FILLCELL_X2 FILLER_80_76 ();
 FILLCELL_X4 FILLER_80_85 ();
 FILLCELL_X1 FILLER_80_89 ();
 FILLCELL_X4 FILLER_80_95 ();
 FILLCELL_X2 FILLER_80_99 ();
 FILLCELL_X2 FILLER_80_133 ();
 FILLCELL_X1 FILLER_80_135 ();
 FILLCELL_X1 FILLER_80_143 ();
 FILLCELL_X1 FILLER_80_161 ();
 FILLCELL_X8 FILLER_80_165 ();
 FILLCELL_X2 FILLER_80_173 ();
 FILLCELL_X8 FILLER_80_180 ();
 FILLCELL_X4 FILLER_80_188 ();
 FILLCELL_X2 FILLER_80_192 ();
 FILLCELL_X1 FILLER_80_194 ();
 FILLCELL_X4 FILLER_80_212 ();
 FILLCELL_X1 FILLER_80_216 ();
 FILLCELL_X8 FILLER_80_227 ();
 FILLCELL_X2 FILLER_80_235 ();
 FILLCELL_X1 FILLER_80_237 ();
 FILLCELL_X32 FILLER_80_241 ();
 FILLCELL_X2 FILLER_80_273 ();
 FILLCELL_X8 FILLER_80_285 ();
 FILLCELL_X4 FILLER_80_293 ();
 FILLCELL_X2 FILLER_80_297 ();
 FILLCELL_X1 FILLER_80_299 ();
 FILLCELL_X8 FILLER_80_314 ();
 FILLCELL_X2 FILLER_80_322 ();
 FILLCELL_X1 FILLER_80_324 ();
 FILLCELL_X2 FILLER_80_335 ();
 FILLCELL_X1 FILLER_80_337 ();
 FILLCELL_X1 FILLER_80_342 ();
 FILLCELL_X8 FILLER_80_348 ();
 FILLCELL_X4 FILLER_80_356 ();
 FILLCELL_X2 FILLER_80_360 ();
 FILLCELL_X1 FILLER_80_366 ();
 FILLCELL_X2 FILLER_80_370 ();
 FILLCELL_X2 FILLER_80_389 ();
 FILLCELL_X16 FILLER_80_398 ();
 FILLCELL_X4 FILLER_80_414 ();
 FILLCELL_X2 FILLER_80_418 ();
 FILLCELL_X4 FILLER_80_429 ();
 FILLCELL_X1 FILLER_80_433 ();
 FILLCELL_X4 FILLER_80_437 ();
 FILLCELL_X8 FILLER_80_446 ();
 FILLCELL_X4 FILLER_80_454 ();
 FILLCELL_X2 FILLER_80_458 ();
 FILLCELL_X32 FILLER_80_477 ();
 FILLCELL_X8 FILLER_80_509 ();
 FILLCELL_X16 FILLER_80_542 ();
 FILLCELL_X4 FILLER_80_558 ();
 FILLCELL_X2 FILLER_80_562 ();
 FILLCELL_X2 FILLER_80_589 ();
 FILLCELL_X2 FILLER_80_596 ();
 FILLCELL_X4 FILLER_80_619 ();
 FILLCELL_X1 FILLER_80_623 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X2 FILLER_80_632 ();
 FILLCELL_X2 FILLER_80_636 ();
 FILLCELL_X1 FILLER_80_645 ();
 FILLCELL_X2 FILLER_80_659 ();
 FILLCELL_X1 FILLER_80_668 ();
 FILLCELL_X16 FILLER_80_672 ();
 FILLCELL_X8 FILLER_80_688 ();
 FILLCELL_X8 FILLER_80_713 ();
 FILLCELL_X2 FILLER_80_728 ();
 FILLCELL_X16 FILLER_80_737 ();
 FILLCELL_X8 FILLER_80_753 ();
 FILLCELL_X2 FILLER_80_761 ();
 FILLCELL_X1 FILLER_80_773 ();
 FILLCELL_X1 FILLER_80_788 ();
 FILLCELL_X1 FILLER_80_793 ();
 FILLCELL_X16 FILLER_80_797 ();
 FILLCELL_X1 FILLER_80_813 ();
 FILLCELL_X16 FILLER_81_1 ();
 FILLCELL_X8 FILLER_81_17 ();
 FILLCELL_X8 FILLER_81_28 ();
 FILLCELL_X2 FILLER_81_36 ();
 FILLCELL_X8 FILLER_81_55 ();
 FILLCELL_X1 FILLER_81_63 ();
 FILLCELL_X16 FILLER_81_89 ();
 FILLCELL_X4 FILLER_81_105 ();
 FILLCELL_X2 FILLER_81_109 ();
 FILLCELL_X4 FILLER_81_144 ();
 FILLCELL_X2 FILLER_81_148 ();
 FILLCELL_X1 FILLER_81_150 ();
 FILLCELL_X8 FILLER_81_154 ();
 FILLCELL_X32 FILLER_81_186 ();
 FILLCELL_X4 FILLER_81_221 ();
 FILLCELL_X1 FILLER_81_229 ();
 FILLCELL_X4 FILLER_81_233 ();
 FILLCELL_X4 FILLER_81_261 ();
 FILLCELL_X8 FILLER_81_272 ();
 FILLCELL_X4 FILLER_81_280 ();
 FILLCELL_X2 FILLER_81_284 ();
 FILLCELL_X1 FILLER_81_293 ();
 FILLCELL_X16 FILLER_81_297 ();
 FILLCELL_X1 FILLER_81_313 ();
 FILLCELL_X8 FILLER_81_321 ();
 FILLCELL_X2 FILLER_81_329 ();
 FILLCELL_X1 FILLER_81_331 ();
 FILLCELL_X4 FILLER_81_349 ();
 FILLCELL_X2 FILLER_81_353 ();
 FILLCELL_X1 FILLER_81_355 ();
 FILLCELL_X32 FILLER_81_380 ();
 FILLCELL_X4 FILLER_81_412 ();
 FILLCELL_X2 FILLER_81_416 ();
 FILLCELL_X1 FILLER_81_418 ();
 FILLCELL_X8 FILLER_81_422 ();
 FILLCELL_X4 FILLER_81_430 ();
 FILLCELL_X2 FILLER_81_434 ();
 FILLCELL_X1 FILLER_81_436 ();
 FILLCELL_X4 FILLER_81_464 ();
 FILLCELL_X8 FILLER_81_475 ();
 FILLCELL_X4 FILLER_81_483 ();
 FILLCELL_X2 FILLER_81_487 ();
 FILLCELL_X1 FILLER_81_489 ();
 FILLCELL_X4 FILLER_81_497 ();
 FILLCELL_X2 FILLER_81_501 ();
 FILLCELL_X1 FILLER_81_503 ();
 FILLCELL_X1 FILLER_81_525 ();
 FILLCELL_X2 FILLER_81_537 ();
 FILLCELL_X1 FILLER_81_543 ();
 FILLCELL_X8 FILLER_81_549 ();
 FILLCELL_X2 FILLER_81_557 ();
 FILLCELL_X8 FILLER_81_582 ();
 FILLCELL_X2 FILLER_81_590 ();
 FILLCELL_X1 FILLER_81_597 ();
 FILLCELL_X2 FILLER_81_609 ();
 FILLCELL_X16 FILLER_81_632 ();
 FILLCELL_X2 FILLER_81_665 ();
 FILLCELL_X1 FILLER_81_667 ();
 FILLCELL_X2 FILLER_81_672 ();
 FILLCELL_X4 FILLER_81_677 ();
 FILLCELL_X1 FILLER_81_681 ();
 FILLCELL_X16 FILLER_81_689 ();
 FILLCELL_X8 FILLER_81_705 ();
 FILLCELL_X4 FILLER_81_713 ();
 FILLCELL_X1 FILLER_81_717 ();
 FILLCELL_X16 FILLER_81_729 ();
 FILLCELL_X2 FILLER_81_745 ();
 FILLCELL_X1 FILLER_81_758 ();
 FILLCELL_X2 FILLER_81_762 ();
 FILLCELL_X1 FILLER_81_767 ();
 FILLCELL_X2 FILLER_81_772 ();
 FILLCELL_X16 FILLER_81_797 ();
 FILLCELL_X1 FILLER_81_813 ();
 FILLCELL_X1 FILLER_82_1 ();
 FILLCELL_X1 FILLER_82_31 ();
 FILLCELL_X2 FILLER_82_42 ();
 FILLCELL_X1 FILLER_82_72 ();
 FILLCELL_X4 FILLER_82_80 ();
 FILLCELL_X2 FILLER_82_84 ();
 FILLCELL_X1 FILLER_82_86 ();
 FILLCELL_X16 FILLER_82_118 ();
 FILLCELL_X8 FILLER_82_134 ();
 FILLCELL_X1 FILLER_82_142 ();
 FILLCELL_X8 FILLER_82_150 ();
 FILLCELL_X4 FILLER_82_158 ();
 FILLCELL_X8 FILLER_82_165 ();
 FILLCELL_X4 FILLER_82_173 ();
 FILLCELL_X1 FILLER_82_177 ();
 FILLCELL_X4 FILLER_82_202 ();
 FILLCELL_X2 FILLER_82_206 ();
 FILLCELL_X4 FILLER_82_218 ();
 FILLCELL_X1 FILLER_82_222 ();
 FILLCELL_X2 FILLER_82_240 ();
 FILLCELL_X1 FILLER_82_242 ();
 FILLCELL_X4 FILLER_82_253 ();
 FILLCELL_X1 FILLER_82_271 ();
 FILLCELL_X4 FILLER_82_279 ();
 FILLCELL_X1 FILLER_82_283 ();
 FILLCELL_X4 FILLER_82_301 ();
 FILLCELL_X2 FILLER_82_305 ();
 FILLCELL_X8 FILLER_82_331 ();
 FILLCELL_X16 FILLER_82_345 ();
 FILLCELL_X2 FILLER_82_361 ();
 FILLCELL_X2 FILLER_82_366 ();
 FILLCELL_X1 FILLER_82_368 ();
 FILLCELL_X8 FILLER_82_376 ();
 FILLCELL_X2 FILLER_82_384 ();
 FILLCELL_X1 FILLER_82_400 ();
 FILLCELL_X8 FILLER_82_453 ();
 FILLCELL_X4 FILLER_82_461 ();
 FILLCELL_X2 FILLER_82_465 ();
 FILLCELL_X8 FILLER_82_474 ();
 FILLCELL_X1 FILLER_82_482 ();
 FILLCELL_X16 FILLER_82_507 ();
 FILLCELL_X2 FILLER_82_523 ();
 FILLCELL_X1 FILLER_82_525 ();
 FILLCELL_X1 FILLER_82_530 ();
 FILLCELL_X4 FILLER_82_538 ();
 FILLCELL_X2 FILLER_82_553 ();
 FILLCELL_X4 FILLER_82_574 ();
 FILLCELL_X2 FILLER_82_578 ();
 FILLCELL_X1 FILLER_82_580 ();
 FILLCELL_X8 FILLER_82_602 ();
 FILLCELL_X2 FILLER_82_610 ();
 FILLCELL_X2 FILLER_82_617 ();
 FILLCELL_X1 FILLER_82_619 ();
 FILLCELL_X4 FILLER_82_632 ();
 FILLCELL_X1 FILLER_82_636 ();
 FILLCELL_X1 FILLER_82_641 ();
 FILLCELL_X2 FILLER_82_646 ();
 FILLCELL_X1 FILLER_82_655 ();
 FILLCELL_X2 FILLER_82_663 ();
 FILLCELL_X4 FILLER_82_689 ();
 FILLCELL_X2 FILLER_82_693 ();
 FILLCELL_X1 FILLER_82_695 ();
 FILLCELL_X8 FILLER_82_700 ();
 FILLCELL_X4 FILLER_82_708 ();
 FILLCELL_X8 FILLER_82_724 ();
 FILLCELL_X4 FILLER_82_732 ();
 FILLCELL_X4 FILLER_82_781 ();
 FILLCELL_X1 FILLER_82_785 ();
 FILLCELL_X4 FILLER_82_810 ();
 FILLCELL_X16 FILLER_83_1 ();
 FILLCELL_X8 FILLER_83_17 ();
 FILLCELL_X4 FILLER_83_25 ();
 FILLCELL_X1 FILLER_83_29 ();
 FILLCELL_X16 FILLER_83_47 ();
 FILLCELL_X8 FILLER_83_63 ();
 FILLCELL_X2 FILLER_83_71 ();
 FILLCELL_X1 FILLER_83_73 ();
 FILLCELL_X16 FILLER_83_91 ();
 FILLCELL_X2 FILLER_83_107 ();
 FILLCELL_X1 FILLER_83_109 ();
 FILLCELL_X1 FILLER_83_114 ();
 FILLCELL_X4 FILLER_83_118 ();
 FILLCELL_X1 FILLER_83_122 ();
 FILLCELL_X1 FILLER_83_127 ();
 FILLCELL_X1 FILLER_83_132 ();
 FILLCELL_X4 FILLER_83_140 ();
 FILLCELL_X2 FILLER_83_144 ();
 FILLCELL_X1 FILLER_83_146 ();
 FILLCELL_X4 FILLER_83_185 ();
 FILLCELL_X2 FILLER_83_189 ();
 FILLCELL_X4 FILLER_83_195 ();
 FILLCELL_X2 FILLER_83_202 ();
 FILLCELL_X16 FILLER_83_243 ();
 FILLCELL_X4 FILLER_83_259 ();
 FILLCELL_X2 FILLER_83_263 ();
 FILLCELL_X8 FILLER_83_272 ();
 FILLCELL_X2 FILLER_83_304 ();
 FILLCELL_X2 FILLER_83_313 ();
 FILLCELL_X1 FILLER_83_315 ();
 FILLCELL_X1 FILLER_83_319 ();
 FILLCELL_X2 FILLER_83_323 ();
 FILLCELL_X1 FILLER_83_332 ();
 FILLCELL_X4 FILLER_83_347 ();
 FILLCELL_X2 FILLER_83_351 ();
 FILLCELL_X1 FILLER_83_353 ();
 FILLCELL_X8 FILLER_83_357 ();
 FILLCELL_X2 FILLER_83_365 ();
 FILLCELL_X4 FILLER_83_374 ();
 FILLCELL_X8 FILLER_83_406 ();
 FILLCELL_X2 FILLER_83_414 ();
 FILLCELL_X4 FILLER_83_420 ();
 FILLCELL_X8 FILLER_83_427 ();
 FILLCELL_X2 FILLER_83_435 ();
 FILLCELL_X4 FILLER_83_440 ();
 FILLCELL_X2 FILLER_83_444 ();
 FILLCELL_X8 FILLER_83_452 ();
 FILLCELL_X2 FILLER_83_460 ();
 FILLCELL_X2 FILLER_83_466 ();
 FILLCELL_X1 FILLER_83_468 ();
 FILLCELL_X8 FILLER_83_472 ();
 FILLCELL_X4 FILLER_83_480 ();
 FILLCELL_X2 FILLER_83_488 ();
 FILLCELL_X16 FILLER_83_502 ();
 FILLCELL_X2 FILLER_83_518 ();
 FILLCELL_X8 FILLER_83_537 ();
 FILLCELL_X2 FILLER_83_545 ();
 FILLCELL_X8 FILLER_83_559 ();
 FILLCELL_X4 FILLER_83_571 ();
 FILLCELL_X2 FILLER_83_575 ();
 FILLCELL_X1 FILLER_83_577 ();
 FILLCELL_X16 FILLER_83_580 ();
 FILLCELL_X2 FILLER_83_596 ();
 FILLCELL_X8 FILLER_83_609 ();
 FILLCELL_X4 FILLER_83_617 ();
 FILLCELL_X4 FILLER_83_625 ();
 FILLCELL_X2 FILLER_83_629 ();
 FILLCELL_X1 FILLER_83_631 ();
 FILLCELL_X16 FILLER_83_671 ();
 FILLCELL_X8 FILLER_83_687 ();
 FILLCELL_X4 FILLER_83_695 ();
 FILLCELL_X2 FILLER_83_711 ();
 FILLCELL_X8 FILLER_83_722 ();
 FILLCELL_X4 FILLER_83_730 ();
 FILLCELL_X2 FILLER_83_734 ();
 FILLCELL_X8 FILLER_83_739 ();
 FILLCELL_X1 FILLER_83_747 ();
 FILLCELL_X2 FILLER_83_750 ();
 FILLCELL_X8 FILLER_83_756 ();
 FILLCELL_X4 FILLER_83_764 ();
 FILLCELL_X2 FILLER_83_768 ();
 FILLCELL_X4 FILLER_83_773 ();
 FILLCELL_X2 FILLER_83_777 ();
 FILLCELL_X1 FILLER_83_793 ();
 FILLCELL_X2 FILLER_83_797 ();
 FILLCELL_X8 FILLER_83_806 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X2 FILLER_84_43 ();
 FILLCELL_X1 FILLER_84_45 ();
 FILLCELL_X1 FILLER_84_53 ();
 FILLCELL_X8 FILLER_84_89 ();
 FILLCELL_X2 FILLER_84_97 ();
 FILLCELL_X1 FILLER_84_99 ();
 FILLCELL_X4 FILLER_84_148 ();
 FILLCELL_X2 FILLER_84_152 ();
 FILLCELL_X1 FILLER_84_154 ();
 FILLCELL_X16 FILLER_84_162 ();
 FILLCELL_X2 FILLER_84_178 ();
 FILLCELL_X1 FILLER_84_180 ();
 FILLCELL_X2 FILLER_84_198 ();
 FILLCELL_X1 FILLER_84_200 ();
 FILLCELL_X4 FILLER_84_218 ();
 FILLCELL_X2 FILLER_84_222 ();
 FILLCELL_X4 FILLER_84_231 ();
 FILLCELL_X4 FILLER_84_240 ();
 FILLCELL_X2 FILLER_84_254 ();
 FILLCELL_X8 FILLER_84_280 ();
 FILLCELL_X1 FILLER_84_288 ();
 FILLCELL_X8 FILLER_84_299 ();
 FILLCELL_X4 FILLER_84_307 ();
 FILLCELL_X4 FILLER_84_349 ();
 FILLCELL_X2 FILLER_84_353 ();
 FILLCELL_X1 FILLER_84_359 ();
 FILLCELL_X2 FILLER_84_370 ();
 FILLCELL_X1 FILLER_84_372 ();
 FILLCELL_X4 FILLER_84_380 ();
 FILLCELL_X2 FILLER_84_384 ();
 FILLCELL_X1 FILLER_84_386 ();
 FILLCELL_X2 FILLER_84_394 ();
 FILLCELL_X1 FILLER_84_396 ();
 FILLCELL_X4 FILLER_84_404 ();
 FILLCELL_X2 FILLER_84_408 ();
 FILLCELL_X1 FILLER_84_410 ();
 FILLCELL_X2 FILLER_84_428 ();
 FILLCELL_X1 FILLER_84_430 ();
 FILLCELL_X4 FILLER_84_450 ();
 FILLCELL_X2 FILLER_84_454 ();
 FILLCELL_X1 FILLER_84_456 ();
 FILLCELL_X4 FILLER_84_484 ();
 FILLCELL_X2 FILLER_84_488 ();
 FILLCELL_X1 FILLER_84_490 ();
 FILLCELL_X4 FILLER_84_508 ();
 FILLCELL_X2 FILLER_84_512 ();
 FILLCELL_X1 FILLER_84_521 ();
 FILLCELL_X2 FILLER_84_531 ();
 FILLCELL_X1 FILLER_84_533 ();
 FILLCELL_X2 FILLER_84_551 ();
 FILLCELL_X4 FILLER_84_583 ();
 FILLCELL_X2 FILLER_84_587 ();
 FILLCELL_X2 FILLER_84_596 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X16 FILLER_84_632 ();
 FILLCELL_X4 FILLER_84_648 ();
 FILLCELL_X2 FILLER_84_652 ();
 FILLCELL_X2 FILLER_84_658 ();
 FILLCELL_X4 FILLER_84_667 ();
 FILLCELL_X1 FILLER_84_671 ();
 FILLCELL_X1 FILLER_84_676 ();
 FILLCELL_X1 FILLER_84_685 ();
 FILLCELL_X2 FILLER_84_702 ();
 FILLCELL_X2 FILLER_84_719 ();
 FILLCELL_X1 FILLER_84_721 ();
 FILLCELL_X8 FILLER_84_739 ();
 FILLCELL_X4 FILLER_84_747 ();
 FILLCELL_X2 FILLER_84_751 ();
 FILLCELL_X1 FILLER_84_753 ();
 FILLCELL_X16 FILLER_84_764 ();
 FILLCELL_X4 FILLER_84_780 ();
 FILLCELL_X2 FILLER_84_784 ();
 FILLCELL_X16 FILLER_84_793 ();
 FILLCELL_X4 FILLER_84_809 ();
 FILLCELL_X1 FILLER_84_813 ();
 FILLCELL_X16 FILLER_85_1 ();
 FILLCELL_X8 FILLER_85_17 ();
 FILLCELL_X8 FILLER_85_45 ();
 FILLCELL_X2 FILLER_85_53 ();
 FILLCELL_X4 FILLER_85_72 ();
 FILLCELL_X1 FILLER_85_76 ();
 FILLCELL_X2 FILLER_85_84 ();
 FILLCELL_X16 FILLER_85_93 ();
 FILLCELL_X2 FILLER_85_109 ();
 FILLCELL_X16 FILLER_85_114 ();
 FILLCELL_X4 FILLER_85_130 ();
 FILLCELL_X16 FILLER_85_172 ();
 FILLCELL_X4 FILLER_85_188 ();
 FILLCELL_X32 FILLER_85_195 ();
 FILLCELL_X4 FILLER_85_227 ();
 FILLCELL_X2 FILLER_85_231 ();
 FILLCELL_X1 FILLER_85_233 ();
 FILLCELL_X2 FILLER_85_258 ();
 FILLCELL_X1 FILLER_85_260 ();
 FILLCELL_X8 FILLER_85_271 ();
 FILLCELL_X4 FILLER_85_279 ();
 FILLCELL_X8 FILLER_85_290 ();
 FILLCELL_X4 FILLER_85_298 ();
 FILLCELL_X2 FILLER_85_302 ();
 FILLCELL_X4 FILLER_85_328 ();
 FILLCELL_X2 FILLER_85_332 ();
 FILLCELL_X4 FILLER_85_344 ();
 FILLCELL_X2 FILLER_85_348 ();
 FILLCELL_X1 FILLER_85_350 ();
 FILLCELL_X1 FILLER_85_368 ();
 FILLCELL_X1 FILLER_85_374 ();
 FILLCELL_X32 FILLER_85_380 ();
 FILLCELL_X4 FILLER_85_412 ();
 FILLCELL_X4 FILLER_85_419 ();
 FILLCELL_X2 FILLER_85_423 ();
 FILLCELL_X1 FILLER_85_425 ();
 FILLCELL_X8 FILLER_85_460 ();
 FILLCELL_X4 FILLER_85_468 ();
 FILLCELL_X2 FILLER_85_472 ();
 FILLCELL_X1 FILLER_85_474 ();
 FILLCELL_X2 FILLER_85_482 ();
 FILLCELL_X1 FILLER_85_484 ();
 FILLCELL_X1 FILLER_85_488 ();
 FILLCELL_X2 FILLER_85_493 ();
 FILLCELL_X1 FILLER_85_495 ();
 FILLCELL_X4 FILLER_85_511 ();
 FILLCELL_X2 FILLER_85_518 ();
 FILLCELL_X4 FILLER_85_534 ();
 FILLCELL_X8 FILLER_85_545 ();
 FILLCELL_X2 FILLER_85_553 ();
 FILLCELL_X1 FILLER_85_555 ();
 FILLCELL_X8 FILLER_85_571 ();
 FILLCELL_X4 FILLER_85_579 ();
 FILLCELL_X1 FILLER_85_583 ();
 FILLCELL_X4 FILLER_85_591 ();
 FILLCELL_X1 FILLER_85_599 ();
 FILLCELL_X1 FILLER_85_602 ();
 FILLCELL_X1 FILLER_85_608 ();
 FILLCELL_X4 FILLER_85_615 ();
 FILLCELL_X8 FILLER_85_630 ();
 FILLCELL_X4 FILLER_85_645 ();
 FILLCELL_X2 FILLER_85_649 ();
 FILLCELL_X1 FILLER_85_651 ();
 FILLCELL_X8 FILLER_85_659 ();
 FILLCELL_X4 FILLER_85_667 ();
 FILLCELL_X2 FILLER_85_671 ();
 FILLCELL_X1 FILLER_85_687 ();
 FILLCELL_X1 FILLER_85_695 ();
 FILLCELL_X2 FILLER_85_708 ();
 FILLCELL_X2 FILLER_85_722 ();
 FILLCELL_X1 FILLER_85_724 ();
 FILLCELL_X2 FILLER_85_735 ();
 FILLCELL_X1 FILLER_85_737 ();
 FILLCELL_X1 FILLER_85_745 ();
 FILLCELL_X4 FILLER_85_748 ();
 FILLCELL_X2 FILLER_85_752 ();
 FILLCELL_X1 FILLER_85_754 ();
 FILLCELL_X4 FILLER_85_772 ();
 FILLCELL_X1 FILLER_85_776 ();
 FILLCELL_X8 FILLER_85_802 ();
 FILLCELL_X4 FILLER_85_810 ();
 FILLCELL_X16 FILLER_86_1 ();
 FILLCELL_X1 FILLER_86_17 ();
 FILLCELL_X2 FILLER_86_27 ();
 FILLCELL_X8 FILLER_86_54 ();
 FILLCELL_X1 FILLER_86_62 ();
 FILLCELL_X4 FILLER_86_71 ();
 FILLCELL_X2 FILLER_86_75 ();
 FILLCELL_X2 FILLER_86_84 ();
 FILLCELL_X8 FILLER_86_93 ();
 FILLCELL_X4 FILLER_86_101 ();
 FILLCELL_X2 FILLER_86_105 ();
 FILLCELL_X1 FILLER_86_107 ();
 FILLCELL_X16 FILLER_86_125 ();
 FILLCELL_X2 FILLER_86_148 ();
 FILLCELL_X1 FILLER_86_164 ();
 FILLCELL_X2 FILLER_86_174 ();
 FILLCELL_X2 FILLER_86_197 ();
 FILLCELL_X16 FILLER_86_219 ();
 FILLCELL_X8 FILLER_86_235 ();
 FILLCELL_X1 FILLER_86_243 ();
 FILLCELL_X4 FILLER_86_258 ();
 FILLCELL_X8 FILLER_86_267 ();
 FILLCELL_X8 FILLER_86_278 ();
 FILLCELL_X1 FILLER_86_286 ();
 FILLCELL_X8 FILLER_86_300 ();
 FILLCELL_X1 FILLER_86_308 ();
 FILLCELL_X8 FILLER_86_316 ();
 FILLCELL_X1 FILLER_86_324 ();
 FILLCELL_X16 FILLER_86_332 ();
 FILLCELL_X2 FILLER_86_348 ();
 FILLCELL_X1 FILLER_86_350 ();
 FILLCELL_X8 FILLER_86_355 ();
 FILLCELL_X4 FILLER_86_363 ();
 FILLCELL_X2 FILLER_86_367 ();
 FILLCELL_X1 FILLER_86_371 ();
 FILLCELL_X16 FILLER_86_381 ();
 FILLCELL_X2 FILLER_86_397 ();
 FILLCELL_X4 FILLER_86_406 ();
 FILLCELL_X4 FILLER_86_417 ();
 FILLCELL_X1 FILLER_86_421 ();
 FILLCELL_X4 FILLER_86_425 ();
 FILLCELL_X2 FILLER_86_429 ();
 FILLCELL_X1 FILLER_86_431 ();
 FILLCELL_X8 FILLER_86_435 ();
 FILLCELL_X2 FILLER_86_443 ();
 FILLCELL_X1 FILLER_86_445 ();
 FILLCELL_X8 FILLER_86_449 ();
 FILLCELL_X1 FILLER_86_457 ();
 FILLCELL_X4 FILLER_86_461 ();
 FILLCELL_X2 FILLER_86_465 ();
 FILLCELL_X1 FILLER_86_467 ();
 FILLCELL_X16 FILLER_86_501 ();
 FILLCELL_X1 FILLER_86_517 ();
 FILLCELL_X4 FILLER_86_523 ();
 FILLCELL_X1 FILLER_86_527 ();
 FILLCELL_X1 FILLER_86_541 ();
 FILLCELL_X8 FILLER_86_546 ();
 FILLCELL_X2 FILLER_86_554 ();
 FILLCELL_X16 FILLER_86_571 ();
 FILLCELL_X2 FILLER_86_602 ();
 FILLCELL_X2 FILLER_86_628 ();
 FILLCELL_X1 FILLER_86_630 ();
 FILLCELL_X2 FILLER_86_649 ();
 FILLCELL_X16 FILLER_86_671 ();
 FILLCELL_X8 FILLER_86_687 ();
 FILLCELL_X2 FILLER_86_695 ();
 FILLCELL_X4 FILLER_86_700 ();
 FILLCELL_X2 FILLER_86_704 ();
 FILLCELL_X1 FILLER_86_706 ();
 FILLCELL_X4 FILLER_86_714 ();
 FILLCELL_X8 FILLER_86_745 ();
 FILLCELL_X4 FILLER_86_753 ();
 FILLCELL_X2 FILLER_86_757 ();
 FILLCELL_X8 FILLER_86_803 ();
 FILLCELL_X2 FILLER_86_811 ();
 FILLCELL_X1 FILLER_86_813 ();
 FILLCELL_X2 FILLER_87_1 ();
 FILLCELL_X2 FILLER_87_35 ();
 FILLCELL_X16 FILLER_87_47 ();
 FILLCELL_X4 FILLER_87_63 ();
 FILLCELL_X2 FILLER_87_67 ();
 FILLCELL_X2 FILLER_87_137 ();
 FILLCELL_X1 FILLER_87_139 ();
 FILLCELL_X4 FILLER_87_154 ();
 FILLCELL_X2 FILLER_87_158 ();
 FILLCELL_X8 FILLER_87_167 ();
 FILLCELL_X2 FILLER_87_175 ();
 FILLCELL_X1 FILLER_87_177 ();
 FILLCELL_X1 FILLER_87_201 ();
 FILLCELL_X2 FILLER_87_224 ();
 FILLCELL_X1 FILLER_87_226 ();
 FILLCELL_X2 FILLER_87_254 ();
 FILLCELL_X1 FILLER_87_256 ();
 FILLCELL_X4 FILLER_87_281 ();
 FILLCELL_X2 FILLER_87_285 ();
 FILLCELL_X4 FILLER_87_304 ();
 FILLCELL_X2 FILLER_87_308 ();
 FILLCELL_X4 FILLER_87_317 ();
 FILLCELL_X2 FILLER_87_321 ();
 FILLCELL_X4 FILLER_87_330 ();
 FILLCELL_X1 FILLER_87_334 ();
 FILLCELL_X2 FILLER_87_349 ();
 FILLCELL_X1 FILLER_87_351 ();
 FILLCELL_X8 FILLER_87_356 ();
 FILLCELL_X4 FILLER_87_364 ();
 FILLCELL_X1 FILLER_87_368 ();
 FILLCELL_X8 FILLER_87_397 ();
 FILLCELL_X2 FILLER_87_405 ();
 FILLCELL_X16 FILLER_87_424 ();
 FILLCELL_X4 FILLER_87_440 ();
 FILLCELL_X2 FILLER_87_444 ();
 FILLCELL_X2 FILLER_87_477 ();
 FILLCELL_X4 FILLER_87_484 ();
 FILLCELL_X1 FILLER_87_488 ();
 FILLCELL_X16 FILLER_87_492 ();
 FILLCELL_X8 FILLER_87_508 ();
 FILLCELL_X1 FILLER_87_530 ();
 FILLCELL_X2 FILLER_87_548 ();
 FILLCELL_X1 FILLER_87_550 ();
 FILLCELL_X8 FILLER_87_559 ();
 FILLCELL_X2 FILLER_87_567 ();
 FILLCELL_X2 FILLER_87_590 ();
 FILLCELL_X1 FILLER_87_599 ();
 FILLCELL_X8 FILLER_87_621 ();
 FILLCELL_X4 FILLER_87_629 ();
 FILLCELL_X8 FILLER_87_643 ();
 FILLCELL_X4 FILLER_87_651 ();
 FILLCELL_X4 FILLER_87_659 ();
 FILLCELL_X4 FILLER_87_666 ();
 FILLCELL_X1 FILLER_87_670 ();
 FILLCELL_X2 FILLER_87_681 ();
 FILLCELL_X1 FILLER_87_683 ();
 FILLCELL_X4 FILLER_87_724 ();
 FILLCELL_X2 FILLER_87_738 ();
 FILLCELL_X8 FILLER_87_747 ();
 FILLCELL_X4 FILLER_87_755 ();
 FILLCELL_X2 FILLER_87_759 ();
 FILLCELL_X1 FILLER_87_761 ();
 FILLCELL_X4 FILLER_87_769 ();
 FILLCELL_X2 FILLER_87_773 ();
 FILLCELL_X16 FILLER_87_792 ();
 FILLCELL_X4 FILLER_87_808 ();
 FILLCELL_X2 FILLER_87_812 ();
 FILLCELL_X16 FILLER_88_1 ();
 FILLCELL_X1 FILLER_88_17 ();
 FILLCELL_X2 FILLER_88_38 ();
 FILLCELL_X1 FILLER_88_64 ();
 FILLCELL_X16 FILLER_88_79 ();
 FILLCELL_X4 FILLER_88_95 ();
 FILLCELL_X1 FILLER_88_99 ();
 FILLCELL_X1 FILLER_88_116 ();
 FILLCELL_X2 FILLER_88_139 ();
 FILLCELL_X1 FILLER_88_141 ();
 FILLCELL_X8 FILLER_88_145 ();
 FILLCELL_X2 FILLER_88_153 ();
 FILLCELL_X1 FILLER_88_155 ();
 FILLCELL_X8 FILLER_88_163 ();
 FILLCELL_X1 FILLER_88_171 ();
 FILLCELL_X16 FILLER_88_186 ();
 FILLCELL_X2 FILLER_88_202 ();
 FILLCELL_X4 FILLER_88_218 ();
 FILLCELL_X4 FILLER_88_246 ();
 FILLCELL_X16 FILLER_88_257 ();
 FILLCELL_X8 FILLER_88_280 ();
 FILLCELL_X2 FILLER_88_288 ();
 FILLCELL_X1 FILLER_88_290 ();
 FILLCELL_X2 FILLER_88_295 ();
 FILLCELL_X4 FILLER_88_300 ();
 FILLCELL_X2 FILLER_88_304 ();
 FILLCELL_X1 FILLER_88_306 ();
 FILLCELL_X8 FILLER_88_322 ();
 FILLCELL_X1 FILLER_88_330 ();
 FILLCELL_X2 FILLER_88_338 ();
 FILLCELL_X8 FILLER_88_364 ();
 FILLCELL_X4 FILLER_88_372 ();
 FILLCELL_X2 FILLER_88_376 ();
 FILLCELL_X1 FILLER_88_378 ();
 FILLCELL_X8 FILLER_88_400 ();
 FILLCELL_X4 FILLER_88_408 ();
 FILLCELL_X4 FILLER_88_416 ();
 FILLCELL_X4 FILLER_88_423 ();
 FILLCELL_X2 FILLER_88_427 ();
 FILLCELL_X1 FILLER_88_433 ();
 FILLCELL_X4 FILLER_88_437 ();
 FILLCELL_X1 FILLER_88_441 ();
 FILLCELL_X32 FILLER_88_452 ();
 FILLCELL_X2 FILLER_88_498 ();
 FILLCELL_X2 FILLER_88_538 ();
 FILLCELL_X4 FILLER_88_548 ();
 FILLCELL_X1 FILLER_88_552 ();
 FILLCELL_X2 FILLER_88_577 ();
 FILLCELL_X1 FILLER_88_579 ();
 FILLCELL_X4 FILLER_88_587 ();
 FILLCELL_X4 FILLER_88_607 ();
 FILLCELL_X2 FILLER_88_611 ();
 FILLCELL_X4 FILLER_88_615 ();
 FILLCELL_X8 FILLER_88_623 ();
 FILLCELL_X2 FILLER_88_632 ();
 FILLCELL_X8 FILLER_88_651 ();
 FILLCELL_X2 FILLER_88_659 ();
 FILLCELL_X1 FILLER_88_661 ();
 FILLCELL_X1 FILLER_88_666 ();
 FILLCELL_X1 FILLER_88_671 ();
 FILLCELL_X2 FILLER_88_724 ();
 FILLCELL_X2 FILLER_88_730 ();
 FILLCELL_X1 FILLER_88_732 ();
 FILLCELL_X4 FILLER_88_737 ();
 FILLCELL_X1 FILLER_88_741 ();
 FILLCELL_X2 FILLER_88_749 ();
 FILLCELL_X1 FILLER_88_753 ();
 FILLCELL_X4 FILLER_88_768 ();
 FILLCELL_X1 FILLER_88_779 ();
 FILLCELL_X4 FILLER_88_783 ();
 FILLCELL_X2 FILLER_88_787 ();
 FILLCELL_X1 FILLER_88_796 ();
 FILLCELL_X16 FILLER_89_1 ();
 FILLCELL_X8 FILLER_89_17 ();
 FILLCELL_X4 FILLER_89_25 ();
 FILLCELL_X2 FILLER_89_39 ();
 FILLCELL_X2 FILLER_89_45 ();
 FILLCELL_X1 FILLER_89_47 ();
 FILLCELL_X16 FILLER_89_51 ();
 FILLCELL_X4 FILLER_89_74 ();
 FILLCELL_X32 FILLER_89_85 ();
 FILLCELL_X8 FILLER_89_117 ();
 FILLCELL_X2 FILLER_89_125 ();
 FILLCELL_X1 FILLER_89_127 ();
 FILLCELL_X8 FILLER_89_131 ();
 FILLCELL_X2 FILLER_89_139 ();
 FILLCELL_X1 FILLER_89_141 ();
 FILLCELL_X2 FILLER_89_146 ();
 FILLCELL_X1 FILLER_89_148 ();
 FILLCELL_X8 FILLER_89_163 ();
 FILLCELL_X1 FILLER_89_171 ();
 FILLCELL_X4 FILLER_89_181 ();
 FILLCELL_X16 FILLER_89_209 ();
 FILLCELL_X1 FILLER_89_225 ();
 FILLCELL_X2 FILLER_89_246 ();
 FILLCELL_X1 FILLER_89_251 ();
 FILLCELL_X1 FILLER_89_259 ();
 FILLCELL_X2 FILLER_89_267 ();
 FILLCELL_X4 FILLER_89_279 ();
 FILLCELL_X2 FILLER_89_286 ();
 FILLCELL_X16 FILLER_89_293 ();
 FILLCELL_X8 FILLER_89_309 ();
 FILLCELL_X4 FILLER_89_317 ();
 FILLCELL_X2 FILLER_89_321 ();
 FILLCELL_X1 FILLER_89_323 ();
 FILLCELL_X8 FILLER_89_352 ();
 FILLCELL_X1 FILLER_89_360 ();
 FILLCELL_X2 FILLER_89_368 ();
 FILLCELL_X4 FILLER_89_384 ();
 FILLCELL_X8 FILLER_89_395 ();
 FILLCELL_X2 FILLER_89_403 ();
 FILLCELL_X4 FILLER_89_460 ();
 FILLCELL_X1 FILLER_89_464 ();
 FILLCELL_X4 FILLER_89_475 ();
 FILLCELL_X2 FILLER_89_479 ();
 FILLCELL_X8 FILLER_89_500 ();
 FILLCELL_X8 FILLER_89_531 ();
 FILLCELL_X4 FILLER_89_539 ();
 FILLCELL_X1 FILLER_89_553 ();
 FILLCELL_X1 FILLER_89_560 ();
 FILLCELL_X8 FILLER_89_568 ();
 FILLCELL_X4 FILLER_89_576 ();
 FILLCELL_X8 FILLER_89_587 ();
 FILLCELL_X2 FILLER_89_595 ();
 FILLCELL_X1 FILLER_89_597 ();
 FILLCELL_X4 FILLER_89_626 ();
 FILLCELL_X2 FILLER_89_630 ();
 FILLCELL_X2 FILLER_89_656 ();
 FILLCELL_X4 FILLER_89_682 ();
 FILLCELL_X2 FILLER_89_686 ();
 FILLCELL_X2 FILLER_89_692 ();
 FILLCELL_X2 FILLER_89_704 ();
 FILLCELL_X1 FILLER_89_718 ();
 FILLCELL_X1 FILLER_89_722 ();
 FILLCELL_X1 FILLER_89_727 ();
 FILLCELL_X2 FILLER_89_752 ();
 FILLCELL_X2 FILLER_89_764 ();
 FILLCELL_X16 FILLER_89_796 ();
 FILLCELL_X2 FILLER_89_812 ();
 FILLCELL_X8 FILLER_90_1 ();
 FILLCELL_X4 FILLER_90_9 ();
 FILLCELL_X1 FILLER_90_13 ();
 FILLCELL_X1 FILLER_90_35 ();
 FILLCELL_X2 FILLER_90_53 ();
 FILLCELL_X4 FILLER_90_76 ();
 FILLCELL_X1 FILLER_90_80 ();
 FILLCELL_X2 FILLER_90_95 ();
 FILLCELL_X1 FILLER_90_97 ();
 FILLCELL_X8 FILLER_90_119 ();
 FILLCELL_X2 FILLER_90_127 ();
 FILLCELL_X4 FILLER_90_174 ();
 FILLCELL_X2 FILLER_90_178 ();
 FILLCELL_X16 FILLER_90_194 ();
 FILLCELL_X1 FILLER_90_210 ();
 FILLCELL_X8 FILLER_90_214 ();
 FILLCELL_X4 FILLER_90_222 ();
 FILLCELL_X1 FILLER_90_250 ();
 FILLCELL_X1 FILLER_90_256 ();
 FILLCELL_X2 FILLER_90_274 ();
 FILLCELL_X4 FILLER_90_320 ();
 FILLCELL_X8 FILLER_90_337 ();
 FILLCELL_X2 FILLER_90_345 ();
 FILLCELL_X4 FILLER_90_354 ();
 FILLCELL_X1 FILLER_90_358 ();
 FILLCELL_X2 FILLER_90_376 ();
 FILLCELL_X2 FILLER_90_381 ();
 FILLCELL_X1 FILLER_90_383 ();
 FILLCELL_X16 FILLER_90_391 ();
 FILLCELL_X4 FILLER_90_407 ();
 FILLCELL_X2 FILLER_90_411 ();
 FILLCELL_X8 FILLER_90_416 ();
 FILLCELL_X4 FILLER_90_424 ();
 FILLCELL_X2 FILLER_90_428 ();
 FILLCELL_X8 FILLER_90_433 ();
 FILLCELL_X2 FILLER_90_441 ();
 FILLCELL_X8 FILLER_90_485 ();
 FILLCELL_X2 FILLER_90_493 ();
 FILLCELL_X2 FILLER_90_502 ();
 FILLCELL_X1 FILLER_90_504 ();
 FILLCELL_X16 FILLER_90_508 ();
 FILLCELL_X4 FILLER_90_524 ();
 FILLCELL_X16 FILLER_90_544 ();
 FILLCELL_X4 FILLER_90_560 ();
 FILLCELL_X2 FILLER_90_564 ();
 FILLCELL_X8 FILLER_90_573 ();
 FILLCELL_X2 FILLER_90_581 ();
 FILLCELL_X1 FILLER_90_583 ();
 FILLCELL_X8 FILLER_90_588 ();
 FILLCELL_X2 FILLER_90_596 ();
 FILLCELL_X8 FILLER_90_602 ();
 FILLCELL_X2 FILLER_90_610 ();
 FILLCELL_X4 FILLER_90_632 ();
 FILLCELL_X2 FILLER_90_636 ();
 FILLCELL_X1 FILLER_90_638 ();
 FILLCELL_X4 FILLER_90_646 ();
 FILLCELL_X2 FILLER_90_650 ();
 FILLCELL_X1 FILLER_90_652 ();
 FILLCELL_X16 FILLER_90_660 ();
 FILLCELL_X4 FILLER_90_676 ();
 FILLCELL_X4 FILLER_90_697 ();
 FILLCELL_X2 FILLER_90_701 ();
 FILLCELL_X16 FILLER_90_707 ();
 FILLCELL_X4 FILLER_90_723 ();
 FILLCELL_X1 FILLER_90_727 ();
 FILLCELL_X4 FILLER_90_731 ();
 FILLCELL_X1 FILLER_90_735 ();
 FILLCELL_X8 FILLER_90_739 ();
 FILLCELL_X8 FILLER_90_764 ();
 FILLCELL_X2 FILLER_90_772 ();
 FILLCELL_X1 FILLER_90_774 ();
 FILLCELL_X16 FILLER_90_796 ();
 FILLCELL_X2 FILLER_90_812 ();
 FILLCELL_X8 FILLER_91_1 ();
 FILLCELL_X1 FILLER_91_9 ();
 FILLCELL_X2 FILLER_91_34 ();
 FILLCELL_X1 FILLER_91_36 ();
 FILLCELL_X2 FILLER_91_40 ();
 FILLCELL_X1 FILLER_91_45 ();
 FILLCELL_X2 FILLER_91_64 ();
 FILLCELL_X1 FILLER_91_66 ();
 FILLCELL_X2 FILLER_91_71 ();
 FILLCELL_X4 FILLER_91_78 ();
 FILLCELL_X8 FILLER_91_89 ();
 FILLCELL_X2 FILLER_91_97 ();
 FILLCELL_X4 FILLER_91_110 ();
 FILLCELL_X2 FILLER_91_114 ();
 FILLCELL_X4 FILLER_91_146 ();
 FILLCELL_X1 FILLER_91_150 ();
 FILLCELL_X4 FILLER_91_154 ();
 FILLCELL_X1 FILLER_91_158 ();
 FILLCELL_X16 FILLER_91_162 ();
 FILLCELL_X2 FILLER_91_192 ();
 FILLCELL_X1 FILLER_91_194 ();
 FILLCELL_X1 FILLER_91_198 ();
 FILLCELL_X8 FILLER_91_202 ();
 FILLCELL_X4 FILLER_91_210 ();
 FILLCELL_X1 FILLER_91_214 ();
 FILLCELL_X1 FILLER_91_225 ();
 FILLCELL_X8 FILLER_91_238 ();
 FILLCELL_X4 FILLER_91_246 ();
 FILLCELL_X1 FILLER_91_250 ();
 FILLCELL_X8 FILLER_91_253 ();
 FILLCELL_X4 FILLER_91_261 ();
 FILLCELL_X1 FILLER_91_265 ();
 FILLCELL_X2 FILLER_91_279 ();
 FILLCELL_X1 FILLER_91_281 ();
 FILLCELL_X2 FILLER_91_285 ();
 FILLCELL_X2 FILLER_91_308 ();
 FILLCELL_X1 FILLER_91_310 ();
 FILLCELL_X8 FILLER_91_332 ();
 FILLCELL_X2 FILLER_91_340 ();
 FILLCELL_X2 FILLER_91_347 ();
 FILLCELL_X1 FILLER_91_357 ();
 FILLCELL_X2 FILLER_91_361 ();
 FILLCELL_X2 FILLER_91_416 ();
 FILLCELL_X16 FILLER_91_421 ();
 FILLCELL_X8 FILLER_91_437 ();
 FILLCELL_X2 FILLER_91_445 ();
 FILLCELL_X1 FILLER_91_447 ();
 FILLCELL_X16 FILLER_91_454 ();
 FILLCELL_X2 FILLER_91_470 ();
 FILLCELL_X8 FILLER_91_475 ();
 FILLCELL_X4 FILLER_91_483 ();
 FILLCELL_X2 FILLER_91_494 ();
 FILLCELL_X1 FILLER_91_496 ();
 FILLCELL_X4 FILLER_91_500 ();
 FILLCELL_X1 FILLER_91_504 ();
 FILLCELL_X1 FILLER_91_521 ();
 FILLCELL_X4 FILLER_91_557 ();
 FILLCELL_X1 FILLER_91_565 ();
 FILLCELL_X1 FILLER_91_575 ();
 FILLCELL_X4 FILLER_91_602 ();
 FILLCELL_X2 FILLER_91_606 ();
 FILLCELL_X4 FILLER_91_623 ();
 FILLCELL_X1 FILLER_91_627 ();
 FILLCELL_X8 FILLER_91_648 ();
 FILLCELL_X2 FILLER_91_656 ();
 FILLCELL_X1 FILLER_91_658 ();
 FILLCELL_X8 FILLER_91_669 ();
 FILLCELL_X4 FILLER_91_677 ();
 FILLCELL_X2 FILLER_91_681 ();
 FILLCELL_X1 FILLER_91_683 ();
 FILLCELL_X16 FILLER_91_688 ();
 FILLCELL_X4 FILLER_91_704 ();
 FILLCELL_X1 FILLER_91_708 ();
 FILLCELL_X8 FILLER_91_716 ();
 FILLCELL_X2 FILLER_91_724 ();
 FILLCELL_X8 FILLER_91_748 ();
 FILLCELL_X4 FILLER_91_769 ();
 FILLCELL_X1 FILLER_91_782 ();
 FILLCELL_X2 FILLER_91_793 ();
 FILLCELL_X16 FILLER_91_798 ();
 FILLCELL_X16 FILLER_92_1 ();
 FILLCELL_X8 FILLER_92_17 ();
 FILLCELL_X1 FILLER_92_25 ();
 FILLCELL_X8 FILLER_92_29 ();
 FILLCELL_X4 FILLER_92_37 ();
 FILLCELL_X1 FILLER_92_41 ();
 FILLCELL_X16 FILLER_92_59 ();
 FILLCELL_X4 FILLER_92_75 ();
 FILLCELL_X1 FILLER_92_79 ();
 FILLCELL_X4 FILLER_92_94 ();
 FILLCELL_X8 FILLER_92_126 ();
 FILLCELL_X4 FILLER_92_134 ();
 FILLCELL_X2 FILLER_92_138 ();
 FILLCELL_X1 FILLER_92_140 ();
 FILLCELL_X1 FILLER_92_153 ();
 FILLCELL_X1 FILLER_92_157 ();
 FILLCELL_X4 FILLER_92_174 ();
 FILLCELL_X1 FILLER_92_178 ();
 FILLCELL_X8 FILLER_92_200 ();
 FILLCELL_X2 FILLER_92_215 ();
 FILLCELL_X4 FILLER_92_224 ();
 FILLCELL_X2 FILLER_92_228 ();
 FILLCELL_X4 FILLER_92_237 ();
 FILLCELL_X1 FILLER_92_241 ();
 FILLCELL_X2 FILLER_92_266 ();
 FILLCELL_X32 FILLER_92_285 ();
 FILLCELL_X4 FILLER_92_317 ();
 FILLCELL_X1 FILLER_92_321 ();
 FILLCELL_X8 FILLER_92_329 ();
 FILLCELL_X1 FILLER_92_337 ();
 FILLCELL_X4 FILLER_92_362 ();
 FILLCELL_X1 FILLER_92_366 ();
 FILLCELL_X4 FILLER_92_372 ();
 FILLCELL_X1 FILLER_92_376 ();
 FILLCELL_X8 FILLER_92_397 ();
 FILLCELL_X2 FILLER_92_405 ();
 FILLCELL_X4 FILLER_92_424 ();
 FILLCELL_X2 FILLER_92_428 ();
 FILLCELL_X8 FILLER_92_457 ();
 FILLCELL_X1 FILLER_92_465 ();
 FILLCELL_X8 FILLER_92_494 ();
 FILLCELL_X4 FILLER_92_502 ();
 FILLCELL_X2 FILLER_92_506 ();
 FILLCELL_X16 FILLER_92_519 ();
 FILLCELL_X2 FILLER_92_535 ();
 FILLCELL_X1 FILLER_92_537 ();
 FILLCELL_X2 FILLER_92_551 ();
 FILLCELL_X4 FILLER_92_572 ();
 FILLCELL_X2 FILLER_92_576 ();
 FILLCELL_X1 FILLER_92_578 ();
 FILLCELL_X2 FILLER_92_614 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X8 FILLER_92_632 ();
 FILLCELL_X2 FILLER_92_640 ();
 FILLCELL_X1 FILLER_92_642 ();
 FILLCELL_X2 FILLER_92_678 ();
 FILLCELL_X1 FILLER_92_680 ();
 FILLCELL_X8 FILLER_92_702 ();
 FILLCELL_X4 FILLER_92_710 ();
 FILLCELL_X1 FILLER_92_714 ();
 FILLCELL_X4 FILLER_92_722 ();
 FILLCELL_X2 FILLER_92_726 ();
 FILLCELL_X1 FILLER_92_728 ();
 FILLCELL_X2 FILLER_92_732 ();
 FILLCELL_X1 FILLER_92_768 ();
 FILLCELL_X4 FILLER_92_786 ();
 FILLCELL_X1 FILLER_92_790 ();
 FILLCELL_X8 FILLER_92_801 ();
 FILLCELL_X4 FILLER_92_809 ();
 FILLCELL_X1 FILLER_92_813 ();
 FILLCELL_X16 FILLER_93_1 ();
 FILLCELL_X2 FILLER_93_17 ();
 FILLCELL_X1 FILLER_93_19 ();
 FILLCELL_X1 FILLER_93_27 ();
 FILLCELL_X1 FILLER_93_31 ();
 FILLCELL_X16 FILLER_93_42 ();
 FILLCELL_X2 FILLER_93_58 ();
 FILLCELL_X1 FILLER_93_60 ();
 FILLCELL_X2 FILLER_93_69 ();
 FILLCELL_X1 FILLER_93_71 ();
 FILLCELL_X4 FILLER_93_79 ();
 FILLCELL_X1 FILLER_93_83 ();
 FILLCELL_X32 FILLER_93_98 ();
 FILLCELL_X4 FILLER_93_130 ();
 FILLCELL_X2 FILLER_93_134 ();
 FILLCELL_X1 FILLER_93_136 ();
 FILLCELL_X8 FILLER_93_146 ();
 FILLCELL_X8 FILLER_93_171 ();
 FILLCELL_X1 FILLER_93_179 ();
 FILLCELL_X2 FILLER_93_194 ();
 FILLCELL_X4 FILLER_93_213 ();
 FILLCELL_X2 FILLER_93_224 ();
 FILLCELL_X4 FILLER_93_235 ();
 FILLCELL_X16 FILLER_93_246 ();
 FILLCELL_X4 FILLER_93_262 ();
 FILLCELL_X8 FILLER_93_273 ();
 FILLCELL_X2 FILLER_93_288 ();
 FILLCELL_X1 FILLER_93_290 ();
 FILLCELL_X4 FILLER_93_298 ();
 FILLCELL_X1 FILLER_93_302 ();
 FILLCELL_X2 FILLER_93_310 ();
 FILLCELL_X8 FILLER_93_319 ();
 FILLCELL_X2 FILLER_93_327 ();
 FILLCELL_X1 FILLER_93_329 ();
 FILLCELL_X16 FILLER_93_351 ();
 FILLCELL_X1 FILLER_93_367 ();
 FILLCELL_X32 FILLER_93_380 ();
 FILLCELL_X1 FILLER_93_412 ();
 FILLCELL_X4 FILLER_93_417 ();
 FILLCELL_X2 FILLER_93_421 ();
 FILLCELL_X1 FILLER_93_423 ();
 FILLCELL_X1 FILLER_93_451 ();
 FILLCELL_X8 FILLER_93_459 ();
 FILLCELL_X4 FILLER_93_467 ();
 FILLCELL_X1 FILLER_93_471 ();
 FILLCELL_X16 FILLER_93_475 ();
 FILLCELL_X4 FILLER_93_491 ();
 FILLCELL_X2 FILLER_93_495 ();
 FILLCELL_X1 FILLER_93_497 ();
 FILLCELL_X4 FILLER_93_507 ();
 FILLCELL_X2 FILLER_93_523 ();
 FILLCELL_X8 FILLER_93_529 ();
 FILLCELL_X4 FILLER_93_557 ();
 FILLCELL_X2 FILLER_93_561 ();
 FILLCELL_X4 FILLER_93_567 ();
 FILLCELL_X2 FILLER_93_571 ();
 FILLCELL_X1 FILLER_93_573 ();
 FILLCELL_X8 FILLER_93_581 ();
 FILLCELL_X4 FILLER_93_589 ();
 FILLCELL_X2 FILLER_93_593 ();
 FILLCELL_X8 FILLER_93_599 ();
 FILLCELL_X8 FILLER_93_611 ();
 FILLCELL_X8 FILLER_93_623 ();
 FILLCELL_X4 FILLER_93_631 ();
 FILLCELL_X1 FILLER_93_635 ();
 FILLCELL_X4 FILLER_93_638 ();
 FILLCELL_X1 FILLER_93_642 ();
 FILLCELL_X2 FILLER_93_650 ();
 FILLCELL_X1 FILLER_93_652 ();
 FILLCELL_X8 FILLER_93_667 ();
 FILLCELL_X4 FILLER_93_675 ();
 FILLCELL_X2 FILLER_93_679 ();
 FILLCELL_X4 FILLER_93_689 ();
 FILLCELL_X8 FILLER_93_700 ();
 FILLCELL_X2 FILLER_93_708 ();
 FILLCELL_X8 FILLER_93_734 ();
 FILLCELL_X2 FILLER_93_742 ();
 FILLCELL_X4 FILLER_93_750 ();
 FILLCELL_X2 FILLER_93_754 ();
 FILLCELL_X16 FILLER_93_762 ();
 FILLCELL_X2 FILLER_93_780 ();
 FILLCELL_X1 FILLER_93_795 ();
 FILLCELL_X1 FILLER_93_813 ();
 FILLCELL_X4 FILLER_94_1 ();
 FILLCELL_X2 FILLER_94_5 ();
 FILLCELL_X2 FILLER_94_24 ();
 FILLCELL_X2 FILLER_94_50 ();
 FILLCELL_X1 FILLER_94_52 ();
 FILLCELL_X2 FILLER_94_70 ();
 FILLCELL_X1 FILLER_94_72 ();
 FILLCELL_X8 FILLER_94_80 ();
 FILLCELL_X2 FILLER_94_88 ();
 FILLCELL_X1 FILLER_94_94 ();
 FILLCELL_X2 FILLER_94_99 ();
 FILLCELL_X2 FILLER_94_105 ();
 FILLCELL_X2 FILLER_94_111 ();
 FILLCELL_X1 FILLER_94_113 ();
 FILLCELL_X2 FILLER_94_157 ();
 FILLCELL_X8 FILLER_94_179 ();
 FILLCELL_X4 FILLER_94_187 ();
 FILLCELL_X1 FILLER_94_194 ();
 FILLCELL_X1 FILLER_94_198 ();
 FILLCELL_X1 FILLER_94_207 ();
 FILLCELL_X2 FILLER_94_215 ();
 FILLCELL_X2 FILLER_94_224 ();
 FILLCELL_X1 FILLER_94_226 ();
 FILLCELL_X4 FILLER_94_236 ();
 FILLCELL_X2 FILLER_94_250 ();
 FILLCELL_X16 FILLER_94_269 ();
 FILLCELL_X2 FILLER_94_285 ();
 FILLCELL_X1 FILLER_94_304 ();
 FILLCELL_X8 FILLER_94_309 ();
 FILLCELL_X2 FILLER_94_317 ();
 FILLCELL_X1 FILLER_94_319 ();
 FILLCELL_X2 FILLER_94_327 ();
 FILLCELL_X2 FILLER_94_336 ();
 FILLCELL_X1 FILLER_94_338 ();
 FILLCELL_X2 FILLER_94_356 ();
 FILLCELL_X1 FILLER_94_358 ();
 FILLCELL_X1 FILLER_94_362 ();
 FILLCELL_X4 FILLER_94_371 ();
 FILLCELL_X2 FILLER_94_375 ();
 FILLCELL_X1 FILLER_94_377 ();
 FILLCELL_X8 FILLER_94_384 ();
 FILLCELL_X4 FILLER_94_392 ();
 FILLCELL_X2 FILLER_94_396 ();
 FILLCELL_X1 FILLER_94_398 ();
 FILLCELL_X2 FILLER_94_406 ();
 FILLCELL_X1 FILLER_94_408 ();
 FILLCELL_X8 FILLER_94_429 ();
 FILLCELL_X4 FILLER_94_437 ();
 FILLCELL_X2 FILLER_94_441 ();
 FILLCELL_X1 FILLER_94_443 ();
 FILLCELL_X2 FILLER_94_450 ();
 FILLCELL_X1 FILLER_94_452 ();
 FILLCELL_X4 FILLER_94_470 ();
 FILLCELL_X2 FILLER_94_474 ();
 FILLCELL_X4 FILLER_94_490 ();
 FILLCELL_X1 FILLER_94_494 ();
 FILLCELL_X4 FILLER_94_498 ();
 FILLCELL_X2 FILLER_94_502 ();
 FILLCELL_X1 FILLER_94_510 ();
 FILLCELL_X8 FILLER_94_523 ();
 FILLCELL_X4 FILLER_94_531 ();
 FILLCELL_X2 FILLER_94_535 ();
 FILLCELL_X1 FILLER_94_537 ();
 FILLCELL_X1 FILLER_94_542 ();
 FILLCELL_X16 FILLER_94_582 ();
 FILLCELL_X4 FILLER_94_611 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X1 FILLER_94_632 ();
 FILLCELL_X4 FILLER_94_650 ();
 FILLCELL_X4 FILLER_94_662 ();
 FILLCELL_X2 FILLER_94_666 ();
 FILLCELL_X1 FILLER_94_668 ();
 FILLCELL_X1 FILLER_94_676 ();
 FILLCELL_X8 FILLER_94_710 ();
 FILLCELL_X4 FILLER_94_718 ();
 FILLCELL_X8 FILLER_94_729 ();
 FILLCELL_X4 FILLER_94_737 ();
 FILLCELL_X2 FILLER_94_741 ();
 FILLCELL_X8 FILLER_94_763 ();
 FILLCELL_X1 FILLER_94_771 ();
 FILLCELL_X4 FILLER_94_774 ();
 FILLCELL_X4 FILLER_94_788 ();
 FILLCELL_X1 FILLER_94_792 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X8 FILLER_95_33 ();
 FILLCELL_X1 FILLER_95_41 ();
 FILLCELL_X16 FILLER_95_57 ();
 FILLCELL_X1 FILLER_95_97 ();
 FILLCELL_X1 FILLER_95_115 ();
 FILLCELL_X4 FILLER_95_130 ();
 FILLCELL_X1 FILLER_95_134 ();
 FILLCELL_X16 FILLER_95_140 ();
 FILLCELL_X4 FILLER_95_156 ();
 FILLCELL_X2 FILLER_95_160 ();
 FILLCELL_X8 FILLER_95_167 ();
 FILLCELL_X2 FILLER_95_193 ();
 FILLCELL_X1 FILLER_95_199 ();
 FILLCELL_X32 FILLER_95_228 ();
 FILLCELL_X4 FILLER_95_260 ();
 FILLCELL_X1 FILLER_95_264 ();
 FILLCELL_X1 FILLER_95_279 ();
 FILLCELL_X2 FILLER_95_287 ();
 FILLCELL_X2 FILLER_95_296 ();
 FILLCELL_X2 FILLER_95_302 ();
 FILLCELL_X4 FILLER_95_322 ();
 FILLCELL_X4 FILLER_95_347 ();
 FILLCELL_X2 FILLER_95_351 ();
 FILLCELL_X16 FILLER_95_398 ();
 FILLCELL_X2 FILLER_95_414 ();
 FILLCELL_X16 FILLER_95_419 ();
 FILLCELL_X2 FILLER_95_435 ();
 FILLCELL_X2 FILLER_95_444 ();
 FILLCELL_X1 FILLER_95_446 ();
 FILLCELL_X2 FILLER_95_462 ();
 FILLCELL_X1 FILLER_95_474 ();
 FILLCELL_X16 FILLER_95_489 ();
 FILLCELL_X2 FILLER_95_505 ();
 FILLCELL_X1 FILLER_95_507 ();
 FILLCELL_X4 FILLER_95_528 ();
 FILLCELL_X8 FILLER_95_537 ();
 FILLCELL_X1 FILLER_95_545 ();
 FILLCELL_X4 FILLER_95_557 ();
 FILLCELL_X4 FILLER_95_578 ();
 FILLCELL_X2 FILLER_95_582 ();
 FILLCELL_X4 FILLER_95_588 ();
 FILLCELL_X2 FILLER_95_592 ();
 FILLCELL_X2 FILLER_95_610 ();
 FILLCELL_X1 FILLER_95_612 ();
 FILLCELL_X8 FILLER_95_638 ();
 FILLCELL_X4 FILLER_95_646 ();
 FILLCELL_X2 FILLER_95_650 ();
 FILLCELL_X16 FILLER_95_669 ();
 FILLCELL_X4 FILLER_95_685 ();
 FILLCELL_X2 FILLER_95_689 ();
 FILLCELL_X8 FILLER_95_695 ();
 FILLCELL_X2 FILLER_95_703 ();
 FILLCELL_X1 FILLER_95_705 ();
 FILLCELL_X4 FILLER_95_720 ();
 FILLCELL_X1 FILLER_95_724 ();
 FILLCELL_X1 FILLER_95_732 ();
 FILLCELL_X2 FILLER_95_740 ();
 FILLCELL_X1 FILLER_95_742 ();
 FILLCELL_X8 FILLER_95_746 ();
 FILLCELL_X2 FILLER_95_754 ();
 FILLCELL_X1 FILLER_95_756 ();
 FILLCELL_X4 FILLER_95_770 ();
 FILLCELL_X2 FILLER_95_774 ();
 FILLCELL_X1 FILLER_95_776 ();
 FILLCELL_X2 FILLER_95_781 ();
 FILLCELL_X4 FILLER_95_787 ();
 FILLCELL_X4 FILLER_95_808 ();
 FILLCELL_X2 FILLER_95_812 ();
 FILLCELL_X16 FILLER_96_1 ();
 FILLCELL_X8 FILLER_96_17 ();
 FILLCELL_X4 FILLER_96_25 ();
 FILLCELL_X2 FILLER_96_46 ();
 FILLCELL_X8 FILLER_96_65 ();
 FILLCELL_X4 FILLER_96_73 ();
 FILLCELL_X2 FILLER_96_77 ();
 FILLCELL_X1 FILLER_96_79 ();
 FILLCELL_X8 FILLER_96_94 ();
 FILLCELL_X2 FILLER_96_102 ();
 FILLCELL_X4 FILLER_96_112 ();
 FILLCELL_X2 FILLER_96_116 ();
 FILLCELL_X1 FILLER_96_118 ();
 FILLCELL_X4 FILLER_96_126 ();
 FILLCELL_X2 FILLER_96_130 ();
 FILLCELL_X1 FILLER_96_132 ();
 FILLCELL_X4 FILLER_96_154 ();
 FILLCELL_X1 FILLER_96_162 ();
 FILLCELL_X16 FILLER_96_167 ();
 FILLCELL_X2 FILLER_96_183 ();
 FILLCELL_X1 FILLER_96_185 ();
 FILLCELL_X16 FILLER_96_206 ();
 FILLCELL_X1 FILLER_96_222 ();
 FILLCELL_X4 FILLER_96_230 ();
 FILLCELL_X2 FILLER_96_234 ();
 FILLCELL_X1 FILLER_96_236 ();
 FILLCELL_X16 FILLER_96_240 ();
 FILLCELL_X2 FILLER_96_256 ();
 FILLCELL_X16 FILLER_96_279 ();
 FILLCELL_X4 FILLER_96_295 ();
 FILLCELL_X2 FILLER_96_303 ();
 FILLCELL_X4 FILLER_96_319 ();
 FILLCELL_X8 FILLER_96_330 ();
 FILLCELL_X4 FILLER_96_338 ();
 FILLCELL_X2 FILLER_96_342 ();
 FILLCELL_X16 FILLER_96_347 ();
 FILLCELL_X4 FILLER_96_363 ();
 FILLCELL_X1 FILLER_96_367 ();
 FILLCELL_X2 FILLER_96_379 ();
 FILLCELL_X4 FILLER_96_385 ();
 FILLCELL_X16 FILLER_96_396 ();
 FILLCELL_X1 FILLER_96_416 ();
 FILLCELL_X4 FILLER_96_423 ();
 FILLCELL_X1 FILLER_96_427 ();
 FILLCELL_X8 FILLER_96_479 ();
 FILLCELL_X4 FILLER_96_487 ();
 FILLCELL_X2 FILLER_96_491 ();
 FILLCELL_X1 FILLER_96_493 ();
 FILLCELL_X8 FILLER_96_504 ();
 FILLCELL_X4 FILLER_96_512 ();
 FILLCELL_X1 FILLER_96_516 ();
 FILLCELL_X2 FILLER_96_526 ();
 FILLCELL_X2 FILLER_96_532 ();
 FILLCELL_X4 FILLER_96_536 ();
 FILLCELL_X2 FILLER_96_540 ();
 FILLCELL_X4 FILLER_96_565 ();
 FILLCELL_X1 FILLER_96_569 ();
 FILLCELL_X8 FILLER_96_594 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X4 FILLER_96_632 ();
 FILLCELL_X16 FILLER_96_640 ();
 FILLCELL_X8 FILLER_96_656 ();
 FILLCELL_X2 FILLER_96_664 ();
 FILLCELL_X1 FILLER_96_666 ();
 FILLCELL_X4 FILLER_96_676 ();
 FILLCELL_X1 FILLER_96_680 ();
 FILLCELL_X4 FILLER_96_685 ();
 FILLCELL_X2 FILLER_96_689 ();
 FILLCELL_X2 FILLER_96_702 ();
 FILLCELL_X1 FILLER_96_704 ();
 FILLCELL_X4 FILLER_96_712 ();
 FILLCELL_X2 FILLER_96_716 ();
 FILLCELL_X1 FILLER_96_718 ();
 FILLCELL_X1 FILLER_96_743 ();
 FILLCELL_X2 FILLER_96_765 ();
 FILLCELL_X16 FILLER_96_789 ();
 FILLCELL_X8 FILLER_96_805 ();
 FILLCELL_X1 FILLER_96_813 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X2 FILLER_97_33 ();
 FILLCELL_X1 FILLER_97_35 ();
 FILLCELL_X2 FILLER_97_43 ();
 FILLCELL_X2 FILLER_97_48 ();
 FILLCELL_X1 FILLER_97_50 ();
 FILLCELL_X4 FILLER_97_75 ();
 FILLCELL_X2 FILLER_97_79 ();
 FILLCELL_X4 FILLER_97_85 ();
 FILLCELL_X2 FILLER_97_97 ();
 FILLCELL_X16 FILLER_97_116 ();
 FILLCELL_X8 FILLER_97_132 ();
 FILLCELL_X4 FILLER_97_149 ();
 FILLCELL_X1 FILLER_97_153 ();
 FILLCELL_X8 FILLER_97_171 ();
 FILLCELL_X4 FILLER_97_179 ();
 FILLCELL_X2 FILLER_97_183 ();
 FILLCELL_X1 FILLER_97_192 ();
 FILLCELL_X8 FILLER_97_210 ();
 FILLCELL_X4 FILLER_97_218 ();
 FILLCELL_X1 FILLER_97_222 ();
 FILLCELL_X1 FILLER_97_247 ();
 FILLCELL_X2 FILLER_97_269 ();
 FILLCELL_X1 FILLER_97_271 ();
 FILLCELL_X2 FILLER_97_276 ();
 FILLCELL_X4 FILLER_97_281 ();
 FILLCELL_X1 FILLER_97_285 ();
 FILLCELL_X1 FILLER_97_290 ();
 FILLCELL_X1 FILLER_97_294 ();
 FILLCELL_X1 FILLER_97_312 ();
 FILLCELL_X1 FILLER_97_320 ();
 FILLCELL_X2 FILLER_97_328 ();
 FILLCELL_X8 FILLER_97_337 ();
 FILLCELL_X4 FILLER_97_345 ();
 FILLCELL_X2 FILLER_97_349 ();
 FILLCELL_X1 FILLER_97_351 ();
 FILLCELL_X2 FILLER_97_359 ();
 FILLCELL_X4 FILLER_97_368 ();
 FILLCELL_X2 FILLER_97_372 ();
 FILLCELL_X8 FILLER_97_391 ();
 FILLCELL_X2 FILLER_97_399 ();
 FILLCELL_X1 FILLER_97_401 ();
 FILLCELL_X1 FILLER_97_423 ();
 FILLCELL_X8 FILLER_97_427 ();
 FILLCELL_X2 FILLER_97_435 ();
 FILLCELL_X1 FILLER_97_437 ();
 FILLCELL_X1 FILLER_97_441 ();
 FILLCELL_X1 FILLER_97_445 ();
 FILLCELL_X1 FILLER_97_449 ();
 FILLCELL_X2 FILLER_97_453 ();
 FILLCELL_X2 FILLER_97_459 ();
 FILLCELL_X8 FILLER_97_467 ();
 FILLCELL_X4 FILLER_97_475 ();
 FILLCELL_X16 FILLER_97_503 ();
 FILLCELL_X8 FILLER_97_526 ();
 FILLCELL_X1 FILLER_97_541 ();
 FILLCELL_X1 FILLER_97_551 ();
 FILLCELL_X8 FILLER_97_554 ();
 FILLCELL_X4 FILLER_97_562 ();
 FILLCELL_X2 FILLER_97_566 ();
 FILLCELL_X4 FILLER_97_576 ();
 FILLCELL_X2 FILLER_97_580 ();
 FILLCELL_X16 FILLER_97_607 ();
 FILLCELL_X4 FILLER_97_623 ();
 FILLCELL_X2 FILLER_97_627 ();
 FILLCELL_X1 FILLER_97_629 ();
 FILLCELL_X4 FILLER_97_655 ();
 FILLCELL_X1 FILLER_97_708 ();
 FILLCELL_X16 FILLER_97_741 ();
 FILLCELL_X8 FILLER_97_757 ();
 FILLCELL_X4 FILLER_97_765 ();
 FILLCELL_X4 FILLER_97_772 ();
 FILLCELL_X2 FILLER_97_776 ();
 FILLCELL_X16 FILLER_97_784 ();
 FILLCELL_X8 FILLER_97_800 ();
 FILLCELL_X4 FILLER_97_808 ();
 FILLCELL_X2 FILLER_97_812 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X8 FILLER_98_33 ();
 FILLCELL_X1 FILLER_98_41 ();
 FILLCELL_X16 FILLER_98_49 ();
 FILLCELL_X2 FILLER_98_65 ();
 FILLCELL_X1 FILLER_98_67 ();
 FILLCELL_X2 FILLER_98_76 ();
 FILLCELL_X4 FILLER_98_95 ();
 FILLCELL_X2 FILLER_98_99 ();
 FILLCELL_X4 FILLER_98_105 ();
 FILLCELL_X8 FILLER_98_117 ();
 FILLCELL_X2 FILLER_98_146 ();
 FILLCELL_X1 FILLER_98_148 ();
 FILLCELL_X2 FILLER_98_157 ();
 FILLCELL_X4 FILLER_98_167 ();
 FILLCELL_X2 FILLER_98_171 ();
 FILLCELL_X1 FILLER_98_190 ();
 FILLCELL_X4 FILLER_98_197 ();
 FILLCELL_X2 FILLER_98_211 ();
 FILLCELL_X8 FILLER_98_216 ();
 FILLCELL_X2 FILLER_98_224 ();
 FILLCELL_X1 FILLER_98_229 ();
 FILLCELL_X1 FILLER_98_234 ();
 FILLCELL_X1 FILLER_98_239 ();
 FILLCELL_X1 FILLER_98_243 ();
 FILLCELL_X1 FILLER_98_264 ();
 FILLCELL_X8 FILLER_98_299 ();
 FILLCELL_X4 FILLER_98_307 ();
 FILLCELL_X1 FILLER_98_318 ();
 FILLCELL_X16 FILLER_98_333 ();
 FILLCELL_X2 FILLER_98_349 ();
 FILLCELL_X4 FILLER_98_372 ();
 FILLCELL_X1 FILLER_98_376 ();
 FILLCELL_X32 FILLER_98_384 ();
 FILLCELL_X4 FILLER_98_416 ();
 FILLCELL_X1 FILLER_98_420 ();
 FILLCELL_X4 FILLER_98_444 ();
 FILLCELL_X16 FILLER_98_469 ();
 FILLCELL_X2 FILLER_98_485 ();
 FILLCELL_X1 FILLER_98_487 ();
 FILLCELL_X2 FILLER_98_502 ();
 FILLCELL_X1 FILLER_98_525 ();
 FILLCELL_X16 FILLER_98_545 ();
 FILLCELL_X1 FILLER_98_561 ();
 FILLCELL_X4 FILLER_98_579 ();
 FILLCELL_X8 FILLER_98_587 ();
 FILLCELL_X16 FILLER_98_599 ();
 FILLCELL_X8 FILLER_98_615 ();
 FILLCELL_X4 FILLER_98_623 ();
 FILLCELL_X1 FILLER_98_627 ();
 FILLCELL_X1 FILLER_98_636 ();
 FILLCELL_X2 FILLER_98_650 ();
 FILLCELL_X16 FILLER_98_678 ();
 FILLCELL_X2 FILLER_98_694 ();
 FILLCELL_X1 FILLER_98_696 ();
 FILLCELL_X4 FILLER_98_701 ();
 FILLCELL_X4 FILLER_98_709 ();
 FILLCELL_X2 FILLER_98_713 ();
 FILLCELL_X1 FILLER_98_715 ();
 FILLCELL_X4 FILLER_98_744 ();
 FILLCELL_X2 FILLER_98_748 ();
 FILLCELL_X1 FILLER_98_750 ();
 FILLCELL_X4 FILLER_98_767 ();
 FILLCELL_X2 FILLER_98_771 ();
 FILLCELL_X2 FILLER_98_776 ();
 FILLCELL_X1 FILLER_98_778 ();
 FILLCELL_X16 FILLER_98_786 ();
 FILLCELL_X8 FILLER_98_802 ();
 FILLCELL_X4 FILLER_98_810 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X4 FILLER_99_65 ();
 FILLCELL_X8 FILLER_99_86 ();
 FILLCELL_X2 FILLER_99_94 ();
 FILLCELL_X8 FILLER_99_122 ();
 FILLCELL_X8 FILLER_99_134 ();
 FILLCELL_X2 FILLER_99_142 ();
 FILLCELL_X1 FILLER_99_144 ();
 FILLCELL_X4 FILLER_99_149 ();
 FILLCELL_X2 FILLER_99_153 ();
 FILLCELL_X1 FILLER_99_155 ();
 FILLCELL_X4 FILLER_99_160 ();
 FILLCELL_X2 FILLER_99_164 ();
 FILLCELL_X8 FILLER_99_192 ();
 FILLCELL_X4 FILLER_99_200 ();
 FILLCELL_X2 FILLER_99_204 ();
 FILLCELL_X1 FILLER_99_206 ();
 FILLCELL_X1 FILLER_99_211 ();
 FILLCELL_X8 FILLER_99_215 ();
 FILLCELL_X2 FILLER_99_223 ();
 FILLCELL_X1 FILLER_99_225 ();
 FILLCELL_X8 FILLER_99_243 ();
 FILLCELL_X2 FILLER_99_251 ();
 FILLCELL_X1 FILLER_99_253 ();
 FILLCELL_X4 FILLER_99_267 ();
 FILLCELL_X2 FILLER_99_271 ();
 FILLCELL_X1 FILLER_99_273 ();
 FILLCELL_X8 FILLER_99_277 ();
 FILLCELL_X2 FILLER_99_285 ();
 FILLCELL_X8 FILLER_99_290 ();
 FILLCELL_X4 FILLER_99_298 ();
 FILLCELL_X1 FILLER_99_302 ();
 FILLCELL_X16 FILLER_99_341 ();
 FILLCELL_X2 FILLER_99_357 ();
 FILLCELL_X4 FILLER_99_373 ();
 FILLCELL_X1 FILLER_99_377 ();
 FILLCELL_X16 FILLER_99_392 ();
 FILLCELL_X8 FILLER_99_408 ();
 FILLCELL_X1 FILLER_99_416 ();
 FILLCELL_X8 FILLER_99_444 ();
 FILLCELL_X2 FILLER_99_452 ();
 FILLCELL_X4 FILLER_99_471 ();
 FILLCELL_X2 FILLER_99_475 ();
 FILLCELL_X4 FILLER_99_512 ();
 FILLCELL_X1 FILLER_99_520 ();
 FILLCELL_X4 FILLER_99_541 ();
 FILLCELL_X1 FILLER_99_545 ();
 FILLCELL_X8 FILLER_99_563 ();
 FILLCELL_X4 FILLER_99_571 ();
 FILLCELL_X2 FILLER_99_575 ();
 FILLCELL_X1 FILLER_99_577 ();
 FILLCELL_X2 FILLER_99_599 ();
 FILLCELL_X8 FILLER_99_609 ();
 FILLCELL_X4 FILLER_99_617 ();
 FILLCELL_X2 FILLER_99_621 ();
 FILLCELL_X1 FILLER_99_623 ();
 FILLCELL_X1 FILLER_99_662 ();
 FILLCELL_X2 FILLER_99_677 ();
 FILLCELL_X2 FILLER_99_683 ();
 FILLCELL_X8 FILLER_99_689 ();
 FILLCELL_X2 FILLER_99_697 ();
 FILLCELL_X8 FILLER_99_716 ();
 FILLCELL_X2 FILLER_99_724 ();
 FILLCELL_X1 FILLER_99_733 ();
 FILLCELL_X8 FILLER_99_737 ();
 FILLCELL_X1 FILLER_99_745 ();
 FILLCELL_X1 FILLER_99_763 ();
 FILLCELL_X2 FILLER_99_768 ();
 FILLCELL_X16 FILLER_99_797 ();
 FILLCELL_X1 FILLER_99_813 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X16 FILLER_100_65 ();
 FILLCELL_X8 FILLER_100_81 ();
 FILLCELL_X4 FILLER_100_89 ();
 FILLCELL_X2 FILLER_100_93 ();
 FILLCELL_X1 FILLER_100_95 ();
 FILLCELL_X16 FILLER_100_113 ();
 FILLCELL_X8 FILLER_100_129 ();
 FILLCELL_X2 FILLER_100_137 ();
 FILLCELL_X1 FILLER_100_139 ();
 FILLCELL_X1 FILLER_100_157 ();
 FILLCELL_X4 FILLER_100_175 ();
 FILLCELL_X2 FILLER_100_179 ();
 FILLCELL_X1 FILLER_100_181 ();
 FILLCELL_X4 FILLER_100_199 ();
 FILLCELL_X16 FILLER_100_220 ();
 FILLCELL_X8 FILLER_100_236 ();
 FILLCELL_X2 FILLER_100_244 ();
 FILLCELL_X1 FILLER_100_246 ();
 FILLCELL_X8 FILLER_100_264 ();
 FILLCELL_X4 FILLER_100_272 ();
 FILLCELL_X1 FILLER_100_276 ();
 FILLCELL_X8 FILLER_100_284 ();
 FILLCELL_X4 FILLER_100_292 ();
 FILLCELL_X2 FILLER_100_296 ();
 FILLCELL_X1 FILLER_100_302 ();
 FILLCELL_X2 FILLER_100_307 ();
 FILLCELL_X2 FILLER_100_314 ();
 FILLCELL_X4 FILLER_100_324 ();
 FILLCELL_X16 FILLER_100_332 ();
 FILLCELL_X2 FILLER_100_348 ();
 FILLCELL_X1 FILLER_100_350 ();
 FILLCELL_X8 FILLER_100_355 ();
 FILLCELL_X4 FILLER_100_363 ();
 FILLCELL_X4 FILLER_100_371 ();
 FILLCELL_X2 FILLER_100_375 ();
 FILLCELL_X1 FILLER_100_377 ();
 FILLCELL_X16 FILLER_100_386 ();
 FILLCELL_X4 FILLER_100_402 ();
 FILLCELL_X1 FILLER_100_406 ();
 FILLCELL_X2 FILLER_100_424 ();
 FILLCELL_X2 FILLER_100_438 ();
 FILLCELL_X16 FILLER_100_450 ();
 FILLCELL_X8 FILLER_100_466 ();
 FILLCELL_X2 FILLER_100_474 ();
 FILLCELL_X1 FILLER_100_476 ();
 FILLCELL_X16 FILLER_100_484 ();
 FILLCELL_X8 FILLER_100_500 ();
 FILLCELL_X4 FILLER_100_508 ();
 FILLCELL_X1 FILLER_100_512 ();
 FILLCELL_X16 FILLER_100_534 ();
 FILLCELL_X8 FILLER_100_550 ();
 FILLCELL_X2 FILLER_100_558 ();
 FILLCELL_X1 FILLER_100_560 ();
 FILLCELL_X1 FILLER_100_565 ();
 FILLCELL_X8 FILLER_100_570 ();
 FILLCELL_X1 FILLER_100_585 ();
 FILLCELL_X2 FILLER_100_599 ();
 FILLCELL_X1 FILLER_100_601 ();
 FILLCELL_X8 FILLER_100_619 ();
 FILLCELL_X4 FILLER_100_627 ();
 FILLCELL_X16 FILLER_100_632 ();
 FILLCELL_X8 FILLER_100_648 ();
 FILLCELL_X2 FILLER_100_656 ();
 FILLCELL_X2 FILLER_100_662 ();
 FILLCELL_X4 FILLER_100_668 ();
 FILLCELL_X2 FILLER_100_672 ();
 FILLCELL_X1 FILLER_100_691 ();
 FILLCELL_X8 FILLER_100_713 ();
 FILLCELL_X1 FILLER_100_721 ();
 FILLCELL_X8 FILLER_100_739 ();
 FILLCELL_X2 FILLER_100_747 ();
 FILLCELL_X1 FILLER_100_749 ();
 FILLCELL_X4 FILLER_100_767 ();
 FILLCELL_X16 FILLER_100_788 ();
 FILLCELL_X8 FILLER_100_804 ();
 FILLCELL_X2 FILLER_100_812 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X8 FILLER_101_257 ();
 FILLCELL_X4 FILLER_101_299 ();
 FILLCELL_X2 FILLER_101_303 ();
 FILLCELL_X8 FILLER_101_318 ();
 FILLCELL_X2 FILLER_101_326 ();
 FILLCELL_X1 FILLER_101_328 ();
 FILLCELL_X16 FILLER_101_363 ();
 FILLCELL_X16 FILLER_101_396 ();
 FILLCELL_X8 FILLER_101_412 ();
 FILLCELL_X4 FILLER_101_420 ();
 FILLCELL_X8 FILLER_101_454 ();
 FILLCELL_X1 FILLER_101_462 ();
 FILLCELL_X8 FILLER_101_483 ();
 FILLCELL_X1 FILLER_101_491 ();
 FILLCELL_X4 FILLER_101_499 ();
 FILLCELL_X8 FILLER_101_523 ();
 FILLCELL_X2 FILLER_101_531 ();
 FILLCELL_X8 FILLER_101_541 ();
 FILLCELL_X4 FILLER_101_549 ();
 FILLCELL_X1 FILLER_101_553 ();
 FILLCELL_X4 FILLER_101_592 ();
 FILLCELL_X2 FILLER_101_596 ();
 FILLCELL_X1 FILLER_101_602 ();
 FILLCELL_X32 FILLER_101_620 ();
 FILLCELL_X4 FILLER_101_652 ();
 FILLCELL_X1 FILLER_101_656 ();
 FILLCELL_X16 FILLER_101_674 ();
 FILLCELL_X2 FILLER_101_690 ();
 FILLCELL_X16 FILLER_101_708 ();
 FILLCELL_X8 FILLER_101_724 ();
 FILLCELL_X2 FILLER_101_732 ();
 FILLCELL_X1 FILLER_101_734 ();
 FILLCELL_X8 FILLER_101_738 ();
 FILLCELL_X1 FILLER_101_746 ();
 FILLCELL_X32 FILLER_101_750 ();
 FILLCELL_X32 FILLER_101_782 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X16 FILLER_102_225 ();
 FILLCELL_X8 FILLER_102_241 ();
 FILLCELL_X1 FILLER_102_249 ();
 FILLCELL_X1 FILLER_102_277 ();
 FILLCELL_X2 FILLER_102_281 ();
 FILLCELL_X1 FILLER_102_283 ();
 FILLCELL_X8 FILLER_102_287 ();
 FILLCELL_X4 FILLER_102_295 ();
 FILLCELL_X2 FILLER_102_329 ();
 FILLCELL_X1 FILLER_102_331 ();
 FILLCELL_X4 FILLER_102_339 ();
 FILLCELL_X2 FILLER_102_343 ();
 FILLCELL_X4 FILLER_102_348 ();
 FILLCELL_X4 FILLER_102_365 ();
 FILLCELL_X2 FILLER_102_375 ();
 FILLCELL_X1 FILLER_102_377 ();
 FILLCELL_X2 FILLER_102_381 ();
 FILLCELL_X16 FILLER_102_400 ();
 FILLCELL_X4 FILLER_102_416 ();
 FILLCELL_X1 FILLER_102_437 ();
 FILLCELL_X16 FILLER_102_459 ();
 FILLCELL_X1 FILLER_102_475 ();
 FILLCELL_X2 FILLER_102_486 ();
 FILLCELL_X8 FILLER_102_505 ();
 FILLCELL_X4 FILLER_102_513 ();
 FILLCELL_X2 FILLER_102_517 ();
 FILLCELL_X1 FILLER_102_519 ();
 FILLCELL_X4 FILLER_102_524 ();
 FILLCELL_X4 FILLER_102_545 ();
 FILLCELL_X2 FILLER_102_549 ();
 FILLCELL_X1 FILLER_102_551 ();
 FILLCELL_X16 FILLER_102_573 ();
 FILLCELL_X1 FILLER_102_589 ();
 FILLCELL_X32 FILLER_102_598 ();
 FILLCELL_X1 FILLER_102_630 ();
 FILLCELL_X8 FILLER_102_632 ();
 FILLCELL_X2 FILLER_102_640 ();
 FILLCELL_X8 FILLER_102_667 ();
 FILLCELL_X4 FILLER_102_675 ();
 FILLCELL_X2 FILLER_102_683 ();
 FILLCELL_X1 FILLER_102_685 ();
 FILLCELL_X4 FILLER_102_690 ();
 FILLCELL_X1 FILLER_102_694 ();
 FILLCELL_X16 FILLER_102_707 ();
 FILLCELL_X2 FILLER_102_733 ();
 FILLCELL_X1 FILLER_102_742 ();
 FILLCELL_X2 FILLER_102_750 ();
 FILLCELL_X1 FILLER_102_752 ();
 FILLCELL_X32 FILLER_102_761 ();
 FILLCELL_X16 FILLER_102_793 ();
 FILLCELL_X4 FILLER_102_809 ();
 FILLCELL_X1 FILLER_102_813 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X16 FILLER_103_257 ();
 FILLCELL_X2 FILLER_103_273 ();
 FILLCELL_X1 FILLER_103_275 ();
 FILLCELL_X8 FILLER_103_288 ();
 FILLCELL_X4 FILLER_103_296 ();
 FILLCELL_X4 FILLER_103_309 ();
 FILLCELL_X8 FILLER_103_333 ();
 FILLCELL_X1 FILLER_103_341 ();
 FILLCELL_X1 FILLER_103_349 ();
 FILLCELL_X2 FILLER_103_376 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X16 FILLER_103_449 ();
 FILLCELL_X4 FILLER_103_465 ();
 FILLCELL_X1 FILLER_103_469 ();
 FILLCELL_X8 FILLER_103_483 ();
 FILLCELL_X2 FILLER_103_494 ();
 FILLCELL_X8 FILLER_103_499 ();
 FILLCELL_X4 FILLER_103_507 ();
 FILLCELL_X2 FILLER_103_511 ();
 FILLCELL_X1 FILLER_103_513 ();
 FILLCELL_X4 FILLER_103_526 ();
 FILLCELL_X16 FILLER_103_542 ();
 FILLCELL_X4 FILLER_103_558 ();
 FILLCELL_X1 FILLER_103_566 ();
 FILLCELL_X4 FILLER_103_571 ();
 FILLCELL_X1 FILLER_103_575 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X2 FILLER_103_641 ();
 FILLCELL_X1 FILLER_103_643 ();
 FILLCELL_X4 FILLER_103_651 ();
 FILLCELL_X1 FILLER_103_655 ();
 FILLCELL_X2 FILLER_103_660 ();
 FILLCELL_X1 FILLER_103_662 ();
 FILLCELL_X1 FILLER_103_667 ();
 FILLCELL_X1 FILLER_103_672 ();
 FILLCELL_X1 FILLER_103_694 ();
 FILLCELL_X1 FILLER_103_712 ();
 FILLCELL_X32 FILLER_103_764 ();
 FILLCELL_X16 FILLER_103_796 ();
 FILLCELL_X2 FILLER_103_812 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X8 FILLER_104_257 ();
 FILLCELL_X2 FILLER_104_265 ();
 FILLCELL_X4 FILLER_104_312 ();
 FILLCELL_X2 FILLER_104_316 ();
 FILLCELL_X8 FILLER_104_325 ();
 FILLCELL_X4 FILLER_104_333 ();
 FILLCELL_X2 FILLER_104_337 ();
 FILLCELL_X4 FILLER_104_356 ();
 FILLCELL_X2 FILLER_104_360 ();
 FILLCELL_X1 FILLER_104_362 ();
 FILLCELL_X32 FILLER_104_380 ();
 FILLCELL_X32 FILLER_104_412 ();
 FILLCELL_X8 FILLER_104_444 ();
 FILLCELL_X4 FILLER_104_452 ();
 FILLCELL_X2 FILLER_104_456 ();
 FILLCELL_X1 FILLER_104_458 ();
 FILLCELL_X2 FILLER_104_476 ();
 FILLCELL_X1 FILLER_104_490 ();
 FILLCELL_X4 FILLER_104_505 ();
 FILLCELL_X2 FILLER_104_509 ();
 FILLCELL_X1 FILLER_104_528 ();
 FILLCELL_X1 FILLER_104_555 ();
 FILLCELL_X1 FILLER_104_598 ();
 FILLCELL_X8 FILLER_104_616 ();
 FILLCELL_X4 FILLER_104_624 ();
 FILLCELL_X2 FILLER_104_628 ();
 FILLCELL_X1 FILLER_104_630 ();
 FILLCELL_X16 FILLER_104_632 ();
 FILLCELL_X8 FILLER_104_682 ();
 FILLCELL_X2 FILLER_104_690 ();
 FILLCELL_X1 FILLER_104_692 ();
 FILLCELL_X32 FILLER_104_710 ();
 FILLCELL_X32 FILLER_104_742 ();
 FILLCELL_X32 FILLER_104_774 ();
 FILLCELL_X8 FILLER_104_806 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X2 FILLER_105_289 ();
 FILLCELL_X1 FILLER_105_291 ();
 FILLCELL_X4 FILLER_105_309 ();
 FILLCELL_X2 FILLER_105_313 ();
 FILLCELL_X32 FILLER_105_332 ();
 FILLCELL_X32 FILLER_105_364 ();
 FILLCELL_X32 FILLER_105_396 ();
 FILLCELL_X32 FILLER_105_428 ();
 FILLCELL_X2 FILLER_105_460 ();
 FILLCELL_X1 FILLER_105_462 ();
 FILLCELL_X4 FILLER_105_480 ();
 FILLCELL_X2 FILLER_105_484 ();
 FILLCELL_X1 FILLER_105_486 ();
 FILLCELL_X8 FILLER_105_504 ();
 FILLCELL_X1 FILLER_105_512 ();
 FILLCELL_X32 FILLER_105_547 ();
 FILLCELL_X2 FILLER_105_579 ();
 FILLCELL_X32 FILLER_105_598 ();
 FILLCELL_X32 FILLER_105_630 ();
 FILLCELL_X32 FILLER_105_662 ();
 FILLCELL_X32 FILLER_105_694 ();
 FILLCELL_X32 FILLER_105_726 ();
 FILLCELL_X32 FILLER_105_758 ();
 FILLCELL_X16 FILLER_105_790 ();
 FILLCELL_X8 FILLER_105_806 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X4 FILLER_106_481 ();
 FILLCELL_X1 FILLER_106_485 ();
 FILLCELL_X32 FILLER_106_503 ();
 FILLCELL_X32 FILLER_106_535 ();
 FILLCELL_X32 FILLER_106_567 ();
 FILLCELL_X32 FILLER_106_599 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X16 FILLER_106_792 ();
 FILLCELL_X4 FILLER_106_808 ();
 FILLCELL_X2 FILLER_106_812 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X16 FILLER_107_577 ();
 FILLCELL_X8 FILLER_107_593 ();
 FILLCELL_X2 FILLER_107_601 ();
 FILLCELL_X1 FILLER_107_603 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X8 FILLER_107_801 ();
 FILLCELL_X4 FILLER_107_809 ();
 FILLCELL_X1 FILLER_107_813 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X32 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_760 ();
 FILLCELL_X16 FILLER_108_792 ();
 FILLCELL_X4 FILLER_108_808 ();
 FILLCELL_X2 FILLER_108_812 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X16 FILLER_109_385 ();
 FILLCELL_X8 FILLER_109_401 ();
 FILLCELL_X32 FILLER_109_413 ();
 FILLCELL_X16 FILLER_109_445 ();
 FILLCELL_X8 FILLER_109_461 ();
 FILLCELL_X1 FILLER_109_472 ();
 FILLCELL_X8 FILLER_109_476 ();
 FILLCELL_X4 FILLER_109_484 ();
 FILLCELL_X2 FILLER_109_488 ();
 FILLCELL_X4 FILLER_109_493 ();
 FILLCELL_X2 FILLER_109_497 ();
 FILLCELL_X16 FILLER_109_502 ();
 FILLCELL_X4 FILLER_109_518 ();
 FILLCELL_X32 FILLER_109_528 ();
 FILLCELL_X16 FILLER_109_560 ();
 FILLCELL_X8 FILLER_109_576 ();
 FILLCELL_X2 FILLER_109_584 ();
 FILLCELL_X32 FILLER_109_590 ();
 FILLCELL_X8 FILLER_109_622 ();
 FILLCELL_X1 FILLER_109_630 ();
 FILLCELL_X32 FILLER_109_632 ();
 FILLCELL_X32 FILLER_109_664 ();
 FILLCELL_X32 FILLER_109_696 ();
 FILLCELL_X32 FILLER_109_728 ();
 FILLCELL_X32 FILLER_109_760 ();
 FILLCELL_X16 FILLER_109_792 ();
 FILLCELL_X4 FILLER_109_808 ();
 FILLCELL_X2 FILLER_109_812 ();
endmodule
