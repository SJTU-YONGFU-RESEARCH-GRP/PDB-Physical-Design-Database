module barrel_shifter (rotate,
    shift_direction,
    data_in,
    data_out,
    shift_amount);
 input rotate;
 input shift_direction;
 input [31:0] data_in;
 output [31:0] data_out;
 input [4:0] shift_amount;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire net56;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire net3;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire net67;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire net44;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire net1;
 wire net2;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net48;
 wire net51;
 wire net54;
 wire net57;
 wire net65;
 wire net66;
 wire net105;
 wire net68;
 wire net69;
 wire net70;

 BUF_X32 _0928_ (.A(shift_amount[0]),
    .Z(_0677_));
 INV_X32 _0929_ (.A(_0677_),
    .ZN(_0688_));
 BUF_X32 _0930_ (.A(_0688_),
    .Z(_0698_));
 BUF_X32 _0931_ (.A(_0698_),
    .Z(_0709_));
 BUF_X16 clone7 (.A(_0698_),
    .Z(net44));
 BUF_X4 _0933_ (.A(shift_amount[1]),
    .Z(_0729_));
 BUF_X8 _0934_ (.A(_0729_),
    .Z(_0739_));
 BUF_X4 clone3 (.A(_0041_),
    .Z(net3));
 INV_X4 _0936_ (.A(_0739_),
    .ZN(_0925_));
 CLKBUF_X3 _0937_ (.A(shift_direction),
    .Z(_0769_));
 BUF_X4 _0938_ (.A(_0769_),
    .Z(_0780_));
 CLKBUF_X3 _0939_ (.A(data_in[0]),
    .Z(_0790_));
 NAND2_X1 _0940_ (.A1(_0790_),
    .A2(net44),
    .ZN(_0800_));
 BUF_X4 _0941_ (.A(shift_amount[4]),
    .Z(_0811_));
 BUF_X4 _0942_ (.A(shift_amount[3]),
    .Z(_0821_));
 BUF_X4 _0943_ (.A(net7),
    .Z(_0832_));
 OR4_X2 _0944_ (.A1(_0811_),
    .A2(_0821_),
    .A3(_0832_),
    .A4(_0729_),
    .ZN(_0842_));
 OAI21_X1 _0945_ (.A(_0780_),
    .B1(_0800_),
    .B2(_0842_),
    .ZN(_0853_));
 BUF_X4 _0946_ (.A(_0677_),
    .Z(_0863_));
 OAI21_X2 _0947_ (.A(net6),
    .B1(_0842_),
    .B2(_0863_),
    .ZN(_0873_));
 BUF_X4 _0948_ (.A(_0873_),
    .Z(_0884_));
 INV_X4 _0949_ (.A(_0811_),
    .ZN(_0894_));
 BUF_X4 clone26 (.A(net69),
    .Z(net67));
 BUF_X8 _0951_ (.A(_0926_),
    .Z(_0914_));
 NOR2_X2 _0952_ (.A1(_0821_),
    .A2(_0832_),
    .ZN(_0000_));
 AOI21_X4 _0953_ (.A(_0894_),
    .B1(_0914_),
    .B2(_0000_),
    .ZN(_0010_));
 BUF_X4 _0954_ (.A(_0832_),
    .Z(_0021_));
 INV_X4 _0955_ (.A(_0914_),
    .ZN(_0031_));
 OR2_X4 _0956_ (.A1(_0811_),
    .A2(_0821_),
    .ZN(_0035_));
 NOR3_X4 _0957_ (.A1(_0021_),
    .A2(_0031_),
    .A3(_0035_),
    .ZN(_0036_));
 NOR3_X2 _0958_ (.A1(_0884_),
    .A2(_0010_),
    .A3(_0036_),
    .ZN(_0037_));
 BUF_X4 _0959_ (.A(_0037_),
    .Z(_0038_));
 BUF_X2 _0960_ (.A(data_in[28]),
    .Z(_0039_));
 BUF_X2 _0961_ (.A(data_in[30]),
    .Z(_0040_));
 BUF_X4 _0962_ (.A(_0927_),
    .Z(_0041_));
 MUX2_X1 _0963_ (.A(_0039_),
    .B(_0040_),
    .S(net69),
    .Z(_0042_));
 BUF_X2 _0964_ (.A(data_in[29]),
    .Z(_0043_));
 CLKBUF_X3 _0965_ (.A(data_in[31]),
    .Z(_0044_));
 BUF_X8 _0966_ (.A(_0041_),
    .Z(_0045_));
 MUX2_X2 _0967_ (.A(_0043_),
    .B(_0044_),
    .S(_0045_),
    .Z(_0046_));
 MUX2_X2 _0968_ (.A(_0042_),
    .B(_0046_),
    .S(_0863_),
    .Z(_0047_));
 BUF_X2 _0969_ (.A(data_in[25]),
    .Z(_0048_));
 BUF_X2 _0970_ (.A(data_in[27]),
    .Z(_0049_));
 BUF_X8 _0971_ (.A(_0041_),
    .Z(_0050_));
 MUX2_X1 _0972_ (.A(_0048_),
    .B(_0049_),
    .S(_0050_),
    .Z(_0051_));
 BUF_X2 _0973_ (.A(data_in[24]),
    .Z(_0052_));
 BUF_X2 _0974_ (.A(data_in[26]),
    .Z(_0053_));
 BUF_X8 _0975_ (.A(_0041_),
    .Z(_0054_));
 MUX2_X1 _0976_ (.A(_0052_),
    .B(_0053_),
    .S(_0054_),
    .Z(_0055_));
 BUF_X4 _0977_ (.A(_0688_),
    .Z(_0056_));
 MUX2_X1 _0978_ (.A(_0051_),
    .B(_0055_),
    .S(_0056_),
    .Z(_0057_));
 XOR2_X2 _0979_ (.A(_0832_),
    .B(_0926_),
    .Z(_0058_));
 BUF_X4 _0980_ (.A(_0058_),
    .Z(_0059_));
 MUX2_X1 _0981_ (.A(_0047_),
    .B(_0057_),
    .S(_0059_),
    .Z(_0060_));
 BUF_X2 _0982_ (.A(data_in[21]),
    .Z(_0061_));
 BUF_X2 _0983_ (.A(data_in[23]),
    .Z(_0062_));
 MUX2_X1 _0984_ (.A(_0061_),
    .B(_0062_),
    .S(_0050_),
    .Z(_0063_));
 BUF_X2 _0985_ (.A(data_in[20]),
    .Z(_0064_));
 BUF_X2 _0986_ (.A(data_in[22]),
    .Z(_0065_));
 MUX2_X1 _0987_ (.A(_0064_),
    .B(_0065_),
    .S(_0054_),
    .Z(_0066_));
 MUX2_X2 _0988_ (.A(_0063_),
    .B(_0066_),
    .S(_0056_),
    .Z(_0067_));
 BUF_X2 _0989_ (.A(data_in[17]),
    .Z(_0068_));
 BUF_X2 _0990_ (.A(data_in[19]),
    .Z(_0069_));
 MUX2_X1 _0991_ (.A(_0068_),
    .B(_0069_),
    .S(_0050_),
    .Z(_0070_));
 BUF_X2 _0992_ (.A(data_in[16]),
    .Z(_0071_));
 BUF_X2 _0993_ (.A(data_in[18]),
    .Z(_0072_));
 MUX2_X1 _0994_ (.A(_0071_),
    .B(_0072_),
    .S(_0054_),
    .Z(_0073_));
 MUX2_X1 _0995_ (.A(_0070_),
    .B(_0073_),
    .S(_0056_),
    .Z(_0074_));
 BUF_X4 _0996_ (.A(_0058_),
    .Z(_0075_));
 MUX2_X1 _0997_ (.A(_0067_),
    .B(_0074_),
    .S(_0075_),
    .Z(_0076_));
 INV_X4 _0998_ (.A(_0821_),
    .ZN(_0077_));
 NOR3_X4 _0999_ (.A1(net7),
    .A2(_0677_),
    .A3(_0729_),
    .ZN(_0078_));
 XNOR2_X2 _1000_ (.A(_0077_),
    .B(_0078_),
    .ZN(_0079_));
 BUF_X4 _1001_ (.A(_0079_),
    .Z(_0080_));
 MUX2_X1 _1002_ (.A(_0060_),
    .B(_0076_),
    .S(_0080_),
    .Z(_0081_));
 OR2_X1 _1003_ (.A1(_0821_),
    .A2(_0832_),
    .ZN(_0082_));
 OAI21_X4 _1004_ (.A(_0811_),
    .B1(_0031_),
    .B2(_0082_),
    .ZN(_0083_));
 INV_X2 _1005_ (.A(_0832_),
    .ZN(_0084_));
 NOR2_X4 _1006_ (.A1(_0811_),
    .A2(_0821_),
    .ZN(_0085_));
 NAND3_X4 _1007_ (.A1(_0084_),
    .A2(_0914_),
    .A3(_0085_),
    .ZN(_0086_));
 AOI21_X2 _1008_ (.A(_0873_),
    .B1(_0083_),
    .B2(_0086_),
    .ZN(_0087_));
 BUF_X4 _1009_ (.A(_0087_),
    .Z(_0088_));
 BUF_X4 _1010_ (.A(_0088_),
    .Z(_0089_));
 BUF_X2 _1011_ (.A(data_in[9]),
    .Z(_0090_));
 BUF_X2 _1012_ (.A(data_in[11]),
    .Z(_0091_));
 BUF_X8 _1013_ (.A(net69),
    .Z(_0092_));
 MUX2_X1 _1014_ (.A(_0090_),
    .B(_0091_),
    .S(net68),
    .Z(_0093_));
 BUF_X2 _1015_ (.A(data_in[8]),
    .Z(_0094_));
 BUF_X2 _1016_ (.A(data_in[10]),
    .Z(_0095_));
 MUX2_X1 _1017_ (.A(_0094_),
    .B(_0095_),
    .S(net3),
    .Z(_0096_));
 MUX2_X1 _1018_ (.A(_0093_),
    .B(_0096_),
    .S(net4),
    .Z(_0097_));
 BUF_X2 _1019_ (.A(data_in[3]),
    .Z(_0098_));
 BUF_X8 _1020_ (.A(_0050_),
    .Z(_0099_));
 MUX2_X1 _1021_ (.A(net5),
    .B(_0098_),
    .S(_0099_),
    .Z(_0100_));
 BUF_X2 _1022_ (.A(data_in[2]),
    .Z(_0101_));
 MUX2_X1 _1023_ (.A(_0790_),
    .B(_0101_),
    .S(_0099_),
    .Z(_0102_));
 BUF_X4 _1024_ (.A(_0056_),
    .Z(_0103_));
 MUX2_X1 _1025_ (.A(_0100_),
    .B(_0102_),
    .S(_0103_),
    .Z(_0104_));
 BUF_X4 _1026_ (.A(_0079_),
    .Z(_0105_));
 MUX2_X1 _1027_ (.A(_0097_),
    .B(_0104_),
    .S(_0105_),
    .Z(_0106_));
 BUF_X2 _1028_ (.A(data_in[13]),
    .Z(_0107_));
 BUF_X2 _1029_ (.A(data_in[15]),
    .Z(_0108_));
 MUX2_X1 _1030_ (.A(_0107_),
    .B(_0108_),
    .S(_0092_),
    .Z(_0109_));
 BUF_X2 _1031_ (.A(data_in[12]),
    .Z(_0110_));
 BUF_X2 _1032_ (.A(data_in[14]),
    .Z(_0111_));
 MUX2_X1 _1033_ (.A(_0110_),
    .B(_0111_),
    .S(net56),
    .Z(_0112_));
 MUX2_X1 _1034_ (.A(_0109_),
    .B(_0112_),
    .S(net4),
    .Z(_0113_));
 BUF_X2 _1035_ (.A(data_in[5]),
    .Z(_0114_));
 BUF_X2 _1036_ (.A(data_in[7]),
    .Z(_0115_));
 MUX2_X1 _1037_ (.A(_0114_),
    .B(_0115_),
    .S(net68),
    .Z(_0116_));
 BUF_X2 _1038_ (.A(data_in[4]),
    .Z(_0117_));
 BUF_X2 _1039_ (.A(data_in[6]),
    .Z(_0118_));
 MUX2_X1 _1040_ (.A(_0117_),
    .B(_0118_),
    .S(net3),
    .Z(_0119_));
 BUF_X4 _1041_ (.A(_0688_),
    .Z(_0120_));
 MUX2_X1 _1042_ (.A(_0116_),
    .B(_0119_),
    .S(_0120_),
    .Z(_0121_));
 MUX2_X1 _1043_ (.A(_0113_),
    .B(_0121_),
    .S(_0079_),
    .Z(_0122_));
 XNOR2_X2 _1044_ (.A(_0832_),
    .B(_0914_),
    .ZN(_0123_));
 BUF_X4 _1045_ (.A(_0123_),
    .Z(_0124_));
 BUF_X4 _1046_ (.A(_0124_),
    .Z(_0125_));
 MUX2_X1 _1047_ (.A(_0106_),
    .B(_0122_),
    .S(_0125_),
    .Z(_0126_));
 AOI221_X2 _1048_ (.A(_0853_),
    .B1(_0038_),
    .B2(_0081_),
    .C1(_0089_),
    .C2(_0126_),
    .ZN(_0127_));
 BUF_X4 _1049_ (.A(_0769_),
    .Z(_0128_));
 BUF_X4 _1050_ (.A(_0128_),
    .Z(_0129_));
 INV_X1 _1051_ (.A(_0790_),
    .ZN(_0130_));
 BUF_X4 _1052_ (.A(_0863_),
    .Z(_0131_));
 BUF_X4 _1053_ (.A(_0131_),
    .Z(_0132_));
 BUF_X4 _1054_ (.A(_0132_),
    .Z(_0133_));
 NOR2_X2 _1055_ (.A1(_0130_),
    .A2(_0133_),
    .ZN(_0134_));
 NAND2_X2 _1056_ (.A1(_0077_),
    .A2(_0078_),
    .ZN(_0135_));
 NOR2_X2 _1057_ (.A1(_0031_),
    .A2(_0135_),
    .ZN(_0136_));
 NAND2_X2 _1058_ (.A1(_0021_),
    .A2(_0031_),
    .ZN(_0137_));
 OR2_X1 _1059_ (.A1(_0863_),
    .A2(_0739_),
    .ZN(_0138_));
 NAND3_X2 _1060_ (.A1(_0084_),
    .A2(_0914_),
    .A3(_0138_),
    .ZN(_0139_));
 AOI21_X4 _1061_ (.A(_0077_),
    .B1(_0137_),
    .B2(_0139_),
    .ZN(_0140_));
 NOR2_X4 _1062_ (.A1(_0136_),
    .A2(_0140_),
    .ZN(_0141_));
 INV_X1 _1063_ (.A(net6),
    .ZN(_0142_));
 AOI21_X4 _1064_ (.A(_0142_),
    .B1(_0078_),
    .B2(_0085_),
    .ZN(_0143_));
 OAI21_X2 _1065_ (.A(_0143_),
    .B1(_0010_),
    .B2(_0036_),
    .ZN(_0144_));
 BUF_X4 _1066_ (.A(_0144_),
    .Z(_0145_));
 NOR3_X4 _1067_ (.A1(_0099_),
    .A2(_0141_),
    .A3(_0145_),
    .ZN(_0146_));
 AOI21_X1 _1068_ (.A(_0129_),
    .B1(_0134_),
    .B2(_0146_),
    .ZN(_0147_));
 CLKBUF_X3 _1069_ (.A(_0739_),
    .Z(_0148_));
 MUX2_X1 _1070_ (.A(_0048_),
    .B(_0049_),
    .S(_0148_),
    .Z(_0149_));
 CLKBUF_X3 _1071_ (.A(_0739_),
    .Z(_0150_));
 MUX2_X1 _1072_ (.A(_0052_),
    .B(_0053_),
    .S(_0150_),
    .Z(_0151_));
 BUF_X4 _1073_ (.A(_0056_),
    .Z(_0152_));
 MUX2_X1 _1074_ (.A(_0149_),
    .B(_0151_),
    .S(_0152_),
    .Z(_0153_));
 BUF_X4 _1075_ (.A(_0729_),
    .Z(_0154_));
 MUX2_X1 _1076_ (.A(_0043_),
    .B(_0044_),
    .S(_0154_),
    .Z(_0155_));
 MUX2_X1 _1077_ (.A(_0039_),
    .B(_0040_),
    .S(_0154_),
    .Z(_0156_));
 BUF_X4 _1078_ (.A(_0688_),
    .Z(_0157_));
 MUX2_X2 _1079_ (.A(_0155_),
    .B(_0156_),
    .S(_0157_),
    .Z(_0158_));
 MUX2_X2 _1080_ (.A(_0153_),
    .B(_0158_),
    .S(_0021_),
    .Z(_0159_));
 MUX2_X1 _1081_ (.A(_0061_),
    .B(_0062_),
    .S(_0150_),
    .Z(_0160_));
 BUF_X4 _1082_ (.A(_0739_),
    .Z(_0161_));
 MUX2_X1 _1083_ (.A(_0064_),
    .B(_0065_),
    .S(_0161_),
    .Z(_0162_));
 MUX2_X1 _1084_ (.A(_0160_),
    .B(_0162_),
    .S(_0103_),
    .Z(_0163_));
 MUX2_X1 _1085_ (.A(_0068_),
    .B(_0069_),
    .S(_0150_),
    .Z(_0164_));
 MUX2_X1 _1086_ (.A(_0071_),
    .B(_0072_),
    .S(_0154_),
    .Z(_0165_));
 MUX2_X1 _1087_ (.A(_0164_),
    .B(_0165_),
    .S(_0103_),
    .Z(_0166_));
 BUF_X4 _1088_ (.A(_0084_),
    .Z(_0167_));
 CLKBUF_X3 _1089_ (.A(_0167_),
    .Z(_0168_));
 MUX2_X1 _1090_ (.A(_0163_),
    .B(_0166_),
    .S(_0168_),
    .Z(_0169_));
 BUF_X4 _1091_ (.A(_0077_),
    .Z(_0170_));
 MUX2_X1 _1092_ (.A(_0159_),
    .B(_0169_),
    .S(_0170_),
    .Z(_0171_));
 CLKBUF_X3 _1093_ (.A(_0739_),
    .Z(_0172_));
 MUX2_X1 _1094_ (.A(_0107_),
    .B(_0108_),
    .S(_0172_),
    .Z(_0173_));
 MUX2_X1 _1095_ (.A(_0110_),
    .B(_0111_),
    .S(_0161_),
    .Z(_0174_));
 MUX2_X1 _1096_ (.A(_0173_),
    .B(_0174_),
    .S(net42),
    .Z(_0175_));
 MUX2_X1 _1097_ (.A(_0090_),
    .B(_0091_),
    .S(_0172_),
    .Z(_0176_));
 MUX2_X1 _1098_ (.A(_0094_),
    .B(_0095_),
    .S(_0172_),
    .Z(_0177_));
 MUX2_X1 _1099_ (.A(_0176_),
    .B(_0177_),
    .S(net42),
    .Z(_0178_));
 CLKBUF_X3 _1100_ (.A(_0167_),
    .Z(_0179_));
 MUX2_X1 _1101_ (.A(_0175_),
    .B(_0178_),
    .S(_0179_),
    .Z(_0180_));
 MUX2_X1 _1102_ (.A(_0114_),
    .B(_0115_),
    .S(_0739_),
    .Z(_0181_));
 MUX2_X1 _1103_ (.A(_0117_),
    .B(_0118_),
    .S(_0739_),
    .Z(_0182_));
 BUF_X4 _1104_ (.A(_0698_),
    .Z(_0183_));
 MUX2_X1 _1105_ (.A(_0181_),
    .B(_0182_),
    .S(_0183_),
    .Z(_0184_));
 MUX2_X1 _1106_ (.A(net5),
    .B(_0098_),
    .S(_0739_),
    .Z(_0185_));
 MUX2_X1 _1107_ (.A(_0790_),
    .B(_0101_),
    .S(_0739_),
    .Z(_0186_));
 MUX2_X1 _1108_ (.A(_0185_),
    .B(_0186_),
    .S(_0183_),
    .Z(_0187_));
 BUF_X4 _1109_ (.A(_0167_),
    .Z(_0188_));
 MUX2_X1 _1110_ (.A(_0184_),
    .B(_0187_),
    .S(_0188_),
    .Z(_0189_));
 BUF_X4 _1111_ (.A(_0077_),
    .Z(_0190_));
 MUX2_X1 _1112_ (.A(_0180_),
    .B(_0189_),
    .S(_0190_),
    .Z(_0191_));
 BUF_X4 _1113_ (.A(_0894_),
    .Z(_0192_));
 MUX2_X1 _1114_ (.A(_0171_),
    .B(_0191_),
    .S(_0192_),
    .Z(_0193_));
 INV_X1 _1115_ (.A(_0193_),
    .ZN(_0194_));
 AOI21_X2 _1116_ (.A(_0127_),
    .B1(_0147_),
    .B2(_0194_),
    .ZN(net8));
 INV_X2 _1117_ (.A(_0769_),
    .ZN(_0195_));
 BUF_X4 _1118_ (.A(_0195_),
    .Z(_0196_));
 BUF_X4 _1119_ (.A(_0811_),
    .Z(_0197_));
 BUF_X4 _1120_ (.A(_0077_),
    .Z(_0198_));
 BUF_X4 _1121_ (.A(_0198_),
    .Z(_0199_));
 MUX2_X1 _1122_ (.A(_0114_),
    .B(_0098_),
    .S(_0739_),
    .Z(_0200_));
 MUX2_X1 _1123_ (.A(_0118_),
    .B(_0117_),
    .S(_0150_),
    .Z(_0201_));
 BUF_X4 _1124_ (.A(_0056_),
    .Z(_0202_));
 MUX2_X1 _1125_ (.A(_0200_),
    .B(_0201_),
    .S(_0202_),
    .Z(_0203_));
 MUX2_X1 _1126_ (.A(_0090_),
    .B(_0115_),
    .S(_0154_),
    .Z(_0204_));
 MUX2_X1 _1127_ (.A(_0095_),
    .B(_0094_),
    .S(_0150_),
    .Z(_0205_));
 MUX2_X1 _1128_ (.A(_0204_),
    .B(_0205_),
    .S(_0202_),
    .Z(_0206_));
 CLKBUF_X3 _1129_ (.A(_0167_),
    .Z(_0207_));
 MUX2_X1 _1130_ (.A(_0203_),
    .B(_0206_),
    .S(_0207_),
    .Z(_0208_));
 MUX2_X2 _1131_ (.A(_0101_),
    .B(_0790_),
    .S(_0154_),
    .Z(_0209_));
 AND2_X2 _1132_ (.A1(net5),
    .A2(_0863_),
    .ZN(_0210_));
 AOI22_X4 _1133_ (.A1(_0183_),
    .A2(_0209_),
    .B1(_0210_),
    .B2(_0925_),
    .ZN(_0211_));
 INV_X1 _1134_ (.A(_0211_),
    .ZN(_0212_));
 BUF_X4 _1135_ (.A(_0021_),
    .Z(_0213_));
 NOR2_X1 _1136_ (.A1(_0077_),
    .A2(_0213_),
    .ZN(_0214_));
 AOI22_X2 _1137_ (.A1(_0199_),
    .A2(_0208_),
    .B1(_0212_),
    .B2(_0214_),
    .ZN(_0215_));
 NOR2_X2 _1138_ (.A1(_0197_),
    .A2(_0215_),
    .ZN(_0216_));
 CLKBUF_X3 _1139_ (.A(_0059_),
    .Z(_0217_));
 BUF_X4 _1140_ (.A(_0217_),
    .Z(_0218_));
 BUF_X4 _1141_ (.A(_0080_),
    .Z(_0219_));
 MUX2_X1 _1142_ (.A(_0062_),
    .B(_0048_),
    .S(_0054_),
    .Z(_0220_));
 MUX2_X1 _1143_ (.A(_0065_),
    .B(_0052_),
    .S(_0092_),
    .Z(_0221_));
 MUX2_X1 _1144_ (.A(_0220_),
    .B(_0221_),
    .S(net4),
    .Z(_0222_));
 NOR2_X1 _1145_ (.A1(_0219_),
    .A2(_0222_),
    .ZN(_0223_));
 BUF_X4 _1146_ (.A(_0821_),
    .Z(_0224_));
 XNOR2_X2 _1147_ (.A(_0224_),
    .B(_0078_),
    .ZN(_0225_));
 BUF_X4 _1148_ (.A(_0225_),
    .Z(_0226_));
 BUF_X4 _1149_ (.A(_0226_),
    .Z(_0227_));
 MUX2_X1 _1150_ (.A(_0108_),
    .B(_0068_),
    .S(_0045_),
    .Z(_0228_));
 MUX2_X1 _1151_ (.A(_0111_),
    .B(_0071_),
    .S(net67),
    .Z(_0229_));
 MUX2_X1 _1152_ (.A(_0228_),
    .B(_0229_),
    .S(_0056_),
    .Z(_0230_));
 NOR2_X1 _1153_ (.A1(_0227_),
    .A2(_0230_),
    .ZN(_0231_));
 NOR4_X2 _1154_ (.A1(_0145_),
    .A2(_0218_),
    .A3(_0223_),
    .A4(_0231_),
    .ZN(_0232_));
 NAND2_X2 _1155_ (.A1(_0083_),
    .A2(_0086_),
    .ZN(_0233_));
 BUF_X4 _1156_ (.A(_0233_),
    .Z(_0234_));
 MUX2_X1 _1157_ (.A(_0069_),
    .B(_0061_),
    .S(_0054_),
    .Z(_0235_));
 MUX2_X1 _1158_ (.A(_0072_),
    .B(_0064_),
    .S(net67),
    .Z(_0236_));
 MUX2_X1 _1159_ (.A(_0235_),
    .B(_0236_),
    .S(net4),
    .Z(_0237_));
 MUX2_X1 _1160_ (.A(_0091_),
    .B(_0107_),
    .S(_0045_),
    .Z(_0238_));
 BUF_X4 clone17 (.A(_0041_),
    .Z(net56));
 MUX2_X1 _1162_ (.A(_0095_),
    .B(_0110_),
    .S(net54),
    .Z(_0240_));
 MUX2_X1 _1163_ (.A(_0238_),
    .B(_0240_),
    .S(_0120_),
    .Z(_0241_));
 MUX2_X1 _1164_ (.A(_0237_),
    .B(_0241_),
    .S(_0079_),
    .Z(_0242_));
 NAND3_X1 _1165_ (.A1(_0234_),
    .A2(_0218_),
    .A3(_0242_),
    .ZN(_0243_));
 INV_X4 _1166_ (.A(net54),
    .ZN(_0244_));
 MUX2_X2 _1167_ (.A(_0040_),
    .B(_0044_),
    .S(_0863_),
    .Z(_0245_));
 AND2_X1 _1168_ (.A1(_0244_),
    .A2(_0245_),
    .ZN(_0246_));
 MUX2_X1 _1169_ (.A(_0049_),
    .B(_0043_),
    .S(net1),
    .Z(_0247_));
 MUX2_X1 _1170_ (.A(_0053_),
    .B(_0039_),
    .S(net67),
    .Z(_0248_));
 MUX2_X1 _1171_ (.A(_0247_),
    .B(_0248_),
    .S(_0698_),
    .Z(_0249_));
 MUX2_X1 _1172_ (.A(_0246_),
    .B(_0249_),
    .S(_0075_),
    .Z(_0250_));
 NOR3_X4 _1173_ (.A1(_0010_),
    .A2(_0036_),
    .A3(_0225_),
    .ZN(_0251_));
 NAND2_X1 _1174_ (.A1(_0250_),
    .A2(_0251_),
    .ZN(_0252_));
 AOI21_X1 _1175_ (.A(_0884_),
    .B1(_0243_),
    .B2(_0252_),
    .ZN(_0253_));
 NOR4_X2 _1176_ (.A1(_0253_),
    .A2(_0216_),
    .A3(_0232_),
    .A4(_0196_),
    .ZN(_0254_));
 BUF_X4 _1177_ (.A(_0088_),
    .Z(_0255_));
 BUF_X4 _1178_ (.A(_0105_),
    .Z(_0256_));
 MUX2_X1 _1179_ (.A(_0095_),
    .B(_0094_),
    .S(_0050_),
    .Z(_0257_));
 MUX2_X1 _1180_ (.A(_0118_),
    .B(_0117_),
    .S(net67),
    .Z(_0258_));
 MUX2_X1 _1181_ (.A(_0257_),
    .B(_0258_),
    .S(_0123_),
    .Z(_0259_));
 MUX2_X1 _1182_ (.A(_0114_),
    .B(_0098_),
    .S(net1),
    .Z(_0260_));
 MUX2_X1 _1183_ (.A(_0090_),
    .B(_0115_),
    .S(net1),
    .Z(_0261_));
 MUX2_X1 _1184_ (.A(_0260_),
    .B(_0261_),
    .S(net105),
    .Z(_0262_));
 MUX2_X1 _1185_ (.A(_0259_),
    .B(_0262_),
    .S(_0132_),
    .Z(_0263_));
 NAND2_X1 _1186_ (.A1(_0256_),
    .A2(_0263_),
    .ZN(_0264_));
 OR3_X2 _1187_ (.A1(_0832_),
    .A2(_0677_),
    .A3(_0729_),
    .ZN(_0265_));
 NAND2_X1 _1188_ (.A1(_0224_),
    .A2(_0265_),
    .ZN(_0266_));
 NAND3_X2 _1189_ (.A1(_0135_),
    .A2(_0266_),
    .A3(_0075_),
    .ZN(_0267_));
 MUX2_X1 _1190_ (.A(_0101_),
    .B(_0790_),
    .S(net56),
    .Z(_0268_));
 AOI22_X2 _1191_ (.A1(_0244_),
    .A2(_0210_),
    .B1(_0268_),
    .B2(_0056_),
    .ZN(_0269_));
 OAI21_X2 _1192_ (.A(_0264_),
    .B1(_0267_),
    .B2(_0269_),
    .ZN(_0270_));
 AOI21_X1 _1193_ (.A(_0129_),
    .B1(_0255_),
    .B2(_0270_),
    .ZN(_0271_));
 MUX2_X1 _1194_ (.A(_0053_),
    .B(_0039_),
    .S(_0161_),
    .Z(_0272_));
 MUX2_X2 _1195_ (.A(_0049_),
    .B(_0043_),
    .S(_0154_),
    .Z(_0273_));
 BUF_X4 _1196_ (.A(_0863_),
    .Z(_0274_));
 MUX2_X2 _1197_ (.A(_0272_),
    .B(_0273_),
    .S(_0274_),
    .Z(_0275_));
 NOR2_X2 _1198_ (.A1(_0167_),
    .A2(_0739_),
    .ZN(_0276_));
 AOI22_X4 _1199_ (.A1(_0188_),
    .A2(_0275_),
    .B1(_0276_),
    .B2(_0245_),
    .ZN(_0277_));
 NAND2_X2 _1200_ (.A1(_0811_),
    .A2(_0198_),
    .ZN(_0278_));
 NOR2_X1 _1201_ (.A1(_0277_),
    .A2(_0278_),
    .ZN(_0279_));
 MUX2_X1 _1202_ (.A(_0062_),
    .B(_0048_),
    .S(_0161_),
    .Z(_0280_));
 MUX2_X1 _1203_ (.A(_0065_),
    .B(_0052_),
    .S(_0150_),
    .Z(_0281_));
 MUX2_X1 _1204_ (.A(_0280_),
    .B(_0281_),
    .S(_0157_),
    .Z(_0282_));
 MUX2_X1 _1205_ (.A(_0069_),
    .B(_0061_),
    .S(_0161_),
    .Z(_0283_));
 MUX2_X1 _1206_ (.A(_0072_),
    .B(_0064_),
    .S(_0150_),
    .Z(_0284_));
 MUX2_X1 _1207_ (.A(_0283_),
    .B(_0284_),
    .S(_0157_),
    .Z(_0285_));
 MUX2_X1 _1208_ (.A(_0282_),
    .B(_0285_),
    .S(_0168_),
    .Z(_0286_));
 MUX2_X1 _1209_ (.A(_0108_),
    .B(_0068_),
    .S(_0154_),
    .Z(_0287_));
 MUX2_X1 _1210_ (.A(_0111_),
    .B(_0071_),
    .S(_0150_),
    .Z(_0288_));
 MUX2_X1 _1211_ (.A(_0287_),
    .B(_0288_),
    .S(_0157_),
    .Z(_0289_));
 MUX2_X1 _1212_ (.A(_0091_),
    .B(_0107_),
    .S(_0161_),
    .Z(_0290_));
 MUX2_X1 _1213_ (.A(_0095_),
    .B(_0110_),
    .S(_0172_),
    .Z(_0291_));
 MUX2_X1 _1214_ (.A(_0290_),
    .B(_0291_),
    .S(net42),
    .Z(_0292_));
 MUX2_X1 _1215_ (.A(_0289_),
    .B(_0292_),
    .S(_0188_),
    .Z(_0293_));
 BUF_X4 _1216_ (.A(_0190_),
    .Z(_0294_));
 MUX2_X1 _1217_ (.A(_0286_),
    .B(_0293_),
    .S(_0294_),
    .Z(_0295_));
 AOI21_X2 _1218_ (.A(_0279_),
    .B1(_0295_),
    .B2(_0192_),
    .ZN(_0296_));
 AOI21_X2 _1219_ (.A(_0254_),
    .B1(_0271_),
    .B2(_0296_),
    .ZN(net9));
 MUX2_X1 _1220_ (.A(_0115_),
    .B(_0114_),
    .S(_0148_),
    .Z(_0297_));
 MUX2_X1 _1221_ (.A(_0201_),
    .B(_0297_),
    .S(_0152_),
    .Z(_0298_));
 MUX2_X1 _1222_ (.A(_0091_),
    .B(_0090_),
    .S(_0148_),
    .Z(_0299_));
 MUX2_X1 _1223_ (.A(_0205_),
    .B(_0299_),
    .S(_0103_),
    .Z(_0300_));
 MUX2_X1 _1224_ (.A(_0298_),
    .B(_0300_),
    .S(_0179_),
    .Z(_0301_));
 MUX2_X1 _1225_ (.A(_0098_),
    .B(net5),
    .S(_0739_),
    .Z(_0302_));
 MUX2_X2 _1226_ (.A(_0209_),
    .B(_0302_),
    .S(_0120_),
    .Z(_0303_));
 AOI22_X1 _1227_ (.A1(_0199_),
    .A2(_0301_),
    .B1(_0303_),
    .B2(_0214_),
    .ZN(_0304_));
 OR2_X1 _1228_ (.A1(_0197_),
    .A2(_0304_),
    .ZN(_0305_));
 BUF_X4 _1229_ (.A(_0195_),
    .Z(_0306_));
 AOI211_X2 _1230_ (.A(_0884_),
    .B(_0105_),
    .C1(_0086_),
    .C2(_0083_),
    .ZN(_0307_));
 MUX2_X1 _1231_ (.A(_0055_),
    .B(_0220_),
    .S(net2),
    .Z(_0308_));
 MUX2_X1 _1232_ (.A(_0066_),
    .B(_0235_),
    .S(net2),
    .Z(_0309_));
 MUX2_X1 _1233_ (.A(_0308_),
    .B(_0309_),
    .S(_0059_),
    .Z(_0310_));
 AOI21_X1 _1234_ (.A(_0306_),
    .B1(_0307_),
    .B2(_0310_),
    .ZN(_0311_));
 NOR2_X2 _1235_ (.A1(_0884_),
    .A2(_0227_),
    .ZN(_0312_));
 INV_X1 _1236_ (.A(_0044_),
    .ZN(_0313_));
 NOR3_X2 _1237_ (.A1(_0131_),
    .A2(_0313_),
    .A3(_0099_),
    .ZN(_0314_));
 MUX2_X1 _1238_ (.A(_0042_),
    .B(_0247_),
    .S(_0688_),
    .Z(_0315_));
 MUX2_X1 _1239_ (.A(_0314_),
    .B(_0315_),
    .S(_0059_),
    .Z(_0316_));
 MUX2_X1 _1240_ (.A(_0073_),
    .B(_0228_),
    .S(net2),
    .Z(_0317_));
 MUX2_X1 _1241_ (.A(_0112_),
    .B(_0238_),
    .S(net2),
    .Z(_0318_));
 MUX2_X1 _1242_ (.A(_0317_),
    .B(_0318_),
    .S(_0059_),
    .Z(_0319_));
 MUX2_X1 _1243_ (.A(_0316_),
    .B(_0319_),
    .S(_0234_),
    .Z(_0320_));
 NAND2_X1 _1244_ (.A1(_0312_),
    .A2(_0320_),
    .ZN(_0321_));
 AND3_X1 _1245_ (.A1(_0305_),
    .A2(_0311_),
    .A3(_0321_),
    .ZN(_0322_));
 MUX2_X1 _1246_ (.A(_0151_),
    .B(_0280_),
    .S(_0202_),
    .Z(_0323_));
 MUX2_X1 _1247_ (.A(_0162_),
    .B(_0283_),
    .S(_0157_),
    .Z(_0324_));
 MUX2_X1 _1248_ (.A(_0323_),
    .B(_0324_),
    .S(_0207_),
    .Z(_0325_));
 MUX2_X1 _1249_ (.A(_0165_),
    .B(_0287_),
    .S(_0120_),
    .Z(_0326_));
 MUX2_X1 _1250_ (.A(_0174_),
    .B(_0290_),
    .S(_0120_),
    .Z(_0327_));
 MUX2_X1 _1251_ (.A(_0326_),
    .B(_0327_),
    .S(_0167_),
    .Z(_0328_));
 MUX2_X1 _1252_ (.A(_0325_),
    .B(_0328_),
    .S(_0199_),
    .Z(_0329_));
 NAND3_X1 _1253_ (.A1(_0207_),
    .A2(_0133_),
    .A3(_0156_),
    .ZN(_0330_));
 AOI22_X4 _1254_ (.A1(_0167_),
    .A2(_0273_),
    .B1(_0276_),
    .B2(_0044_),
    .ZN(_0331_));
 OAI21_X4 _1255_ (.A(_0330_),
    .B1(_0331_),
    .B2(_0133_),
    .ZN(_0332_));
 NOR2_X4 _1256_ (.A1(_0894_),
    .A2(_0224_),
    .ZN(_0333_));
 AOI22_X2 _1257_ (.A1(_0192_),
    .A2(_0329_),
    .B1(_0332_),
    .B2(_0333_),
    .ZN(_0334_));
 BUF_X4 _1258_ (.A(_0769_),
    .Z(_0335_));
 BUF_X4 _1259_ (.A(_0335_),
    .Z(_0336_));
 MUX2_X1 _1260_ (.A(_0098_),
    .B(net5),
    .S(net67),
    .Z(_0337_));
 MUX2_X2 _1261_ (.A(_0268_),
    .B(_0337_),
    .S(_0698_),
    .Z(_0338_));
 NAND3_X1 _1262_ (.A1(_0227_),
    .A2(_0218_),
    .A3(net65),
    .ZN(_0339_));
 MUX2_X1 _1263_ (.A(_0115_),
    .B(_0114_),
    .S(_0092_),
    .Z(_0340_));
 MUX2_X1 _1264_ (.A(_0258_),
    .B(_0340_),
    .S(_0120_),
    .Z(_0341_));
 OR2_X1 _1265_ (.A1(_0217_),
    .A2(_0341_),
    .ZN(_0342_));
 MUX2_X1 _1266_ (.A(_0091_),
    .B(_0090_),
    .S(_0092_),
    .Z(_0343_));
 MUX2_X1 _1267_ (.A(_0257_),
    .B(_0343_),
    .S(_0157_),
    .Z(_0344_));
 OAI21_X1 _1268_ (.A(_0342_),
    .B1(_0344_),
    .B2(_0124_),
    .ZN(_0345_));
 OAI21_X1 _1269_ (.A(_0339_),
    .B1(_0345_),
    .B2(_0227_),
    .ZN(_0346_));
 AOI21_X1 _1270_ (.A(_0336_),
    .B1(_0255_),
    .B2(_0346_),
    .ZN(_0347_));
 AOI21_X2 _1271_ (.A(_0322_),
    .B1(_0334_),
    .B2(_0347_),
    .ZN(net10));
 NOR2_X2 _1272_ (.A1(_0010_),
    .A2(_0036_),
    .ZN(_0348_));
 BUF_X4 _1273_ (.A(_0348_),
    .Z(_0349_));
 NOR2_X2 _1274_ (.A1(_0349_),
    .A2(_0080_),
    .ZN(_0350_));
 OR2_X1 _1275_ (.A1(_0217_),
    .A2(_0057_),
    .ZN(_0351_));
 BUF_X4 _1276_ (.A(_0124_),
    .Z(_0352_));
 OAI21_X1 _1277_ (.A(_0351_),
    .B1(_0067_),
    .B2(_0352_),
    .ZN(_0353_));
 AOI21_X1 _1278_ (.A(_0884_),
    .B1(_0350_),
    .B2(_0353_),
    .ZN(_0354_));
 AND4_X1 _1279_ (.A1(_0083_),
    .A2(_0086_),
    .A3(_0079_),
    .A4(_0047_),
    .ZN(_0355_));
 AOI21_X1 _1280_ (.A(_0355_),
    .B1(_0113_),
    .B2(_0233_),
    .ZN(_0356_));
 AOI21_X1 _1281_ (.A(_0226_),
    .B1(_0124_),
    .B2(_0074_),
    .ZN(_0357_));
 OAI22_X2 _1282_ (.A1(_0125_),
    .A2(_0356_),
    .B1(_0357_),
    .B2(_0349_),
    .ZN(_0358_));
 NOR2_X2 _1283_ (.A1(_0863_),
    .A2(_0739_),
    .ZN(_0359_));
 NAND3_X1 _1284_ (.A1(_0213_),
    .A2(_0790_),
    .A3(_0359_),
    .ZN(_0360_));
 NAND3_X1 _1285_ (.A1(_0168_),
    .A2(_0133_),
    .A3(_0302_),
    .ZN(_0361_));
 MUX2_X1 _1286_ (.A(_0117_),
    .B(_0101_),
    .S(_0739_),
    .Z(_0362_));
 NAND3_X1 _1287_ (.A1(_0168_),
    .A2(net44),
    .A3(_0362_),
    .ZN(_0363_));
 NAND3_X1 _1288_ (.A1(_0360_),
    .A2(_0361_),
    .A3(_0363_),
    .ZN(_0364_));
 MUX2_X1 _1289_ (.A(_0094_),
    .B(_0118_),
    .S(_0154_),
    .Z(_0365_));
 MUX2_X1 _1290_ (.A(_0297_),
    .B(_0365_),
    .S(_0202_),
    .Z(_0366_));
 MUX2_X1 _1291_ (.A(_0110_),
    .B(_0095_),
    .S(_0154_),
    .Z(_0367_));
 MUX2_X1 _1292_ (.A(_0299_),
    .B(_0367_),
    .S(_0152_),
    .Z(_0368_));
 MUX2_X1 _1293_ (.A(_0366_),
    .B(_0368_),
    .S(_0168_),
    .Z(_0369_));
 MUX2_X1 _1294_ (.A(_0364_),
    .B(_0369_),
    .S(_0198_),
    .Z(_0370_));
 BUF_X4 _1295_ (.A(_0894_),
    .Z(_0371_));
 AOI221_X2 _1296_ (.A(_0306_),
    .B1(_0354_),
    .B2(_0358_),
    .C1(_0370_),
    .C2(_0371_),
    .ZN(_0372_));
 MUX2_X1 _1297_ (.A(_0153_),
    .B(_0163_),
    .S(_0179_),
    .Z(_0373_));
 CLKBUF_X3 _1298_ (.A(_0188_),
    .Z(_0374_));
 MUX2_X1 _1299_ (.A(_0166_),
    .B(_0175_),
    .S(_0374_),
    .Z(_0375_));
 MUX2_X1 _1300_ (.A(_0373_),
    .B(_0375_),
    .S(_0294_),
    .Z(_0376_));
 NAND2_X1 _1301_ (.A1(_0192_),
    .A2(_0376_),
    .ZN(_0377_));
 MUX2_X1 _1302_ (.A(_0340_),
    .B(_0343_),
    .S(net105),
    .Z(_0378_));
 MUX2_X1 _1303_ (.A(_0094_),
    .B(_0118_),
    .S(net1),
    .Z(_0379_));
 MUX2_X1 _1304_ (.A(_0110_),
    .B(_0095_),
    .S(net56),
    .Z(_0380_));
 MUX2_X1 _1305_ (.A(_0379_),
    .B(_0380_),
    .S(net105),
    .Z(_0381_));
 MUX2_X1 _1306_ (.A(_0378_),
    .B(_0381_),
    .S(_0183_),
    .Z(_0382_));
 NAND2_X1 _1307_ (.A1(_0256_),
    .A2(_0382_),
    .ZN(_0383_));
 NOR3_X1 _1308_ (.A1(_0130_),
    .A2(_0132_),
    .A3(_0099_),
    .ZN(_0384_));
 NOR2_X2 _1309_ (.A1(_0021_),
    .A2(_0739_),
    .ZN(_0385_));
 XNOR2_X1 _1310_ (.A(_0224_),
    .B(_0385_),
    .ZN(_0386_));
 NAND2_X1 _1311_ (.A1(_0384_),
    .A2(_0386_),
    .ZN(_0387_));
 MUX2_X1 _1312_ (.A(_0117_),
    .B(_0101_),
    .S(net1),
    .Z(_0388_));
 MUX2_X1 _1313_ (.A(_0337_),
    .B(_0388_),
    .S(_0183_),
    .Z(_0389_));
 NAND2_X1 _1314_ (.A1(_0217_),
    .A2(_0389_),
    .ZN(_0390_));
 OAI221_X2 _1315_ (.A(_0383_),
    .B1(_0387_),
    .B2(_0217_),
    .C1(_0256_),
    .C2(_0390_),
    .ZN(_0391_));
 NOR2_X2 _1316_ (.A1(_0213_),
    .A2(_0278_),
    .ZN(_0392_));
 AOI221_X2 _1317_ (.A(_0128_),
    .B1(_0391_),
    .B2(_0089_),
    .C1(_0392_),
    .C2(_0158_),
    .ZN(_0393_));
 AOI21_X2 _1318_ (.A(_0372_),
    .B1(_0377_),
    .B2(_0393_),
    .ZN(net11));
 MUX2_X2 _1319_ (.A(net5),
    .B(_0790_),
    .S(_0863_),
    .Z(_0394_));
 AND2_X2 _1320_ (.A1(_0244_),
    .A2(_0394_),
    .ZN(_0395_));
 MUX2_X1 _1321_ (.A(_0260_),
    .B(_0388_),
    .S(_0131_),
    .Z(_0396_));
 MUX2_X1 _1322_ (.A(_0395_),
    .B(_0396_),
    .S(_0059_),
    .Z(_0397_));
 MUX2_X1 _1323_ (.A(_0261_),
    .B(_0379_),
    .S(_0131_),
    .Z(_0398_));
 MUX2_X1 _1324_ (.A(_0107_),
    .B(_0091_),
    .S(net56),
    .Z(_0399_));
 MUX2_X1 _1325_ (.A(_0380_),
    .B(_0399_),
    .S(_0698_),
    .Z(_0400_));
 MUX2_X1 _1326_ (.A(_0398_),
    .B(_0400_),
    .S(_0075_),
    .Z(_0401_));
 MUX2_X2 _1327_ (.A(_0397_),
    .B(_0401_),
    .S(_0080_),
    .Z(_0402_));
 MUX2_X1 _1328_ (.A(_0160_),
    .B(_0281_),
    .S(_0274_),
    .Z(_0403_));
 MUX2_X1 _1329_ (.A(_0149_),
    .B(_0272_),
    .S(_0274_),
    .Z(_0404_));
 MUX2_X1 _1330_ (.A(_0403_),
    .B(_0404_),
    .S(_0213_),
    .Z(_0405_));
 NOR2_X1 _1331_ (.A1(_0197_),
    .A2(_0199_),
    .ZN(_0406_));
 AOI221_X2 _1332_ (.A(_0128_),
    .B1(_0402_),
    .B2(_0089_),
    .C1(_0405_),
    .C2(_0406_),
    .ZN(_0407_));
 MUX2_X1 _1333_ (.A(_0164_),
    .B(_0284_),
    .S(_0274_),
    .Z(_0408_));
 MUX2_X1 _1334_ (.A(_0173_),
    .B(_0288_),
    .S(_0132_),
    .Z(_0409_));
 MUX2_X1 _1335_ (.A(_0408_),
    .B(_0409_),
    .S(_0179_),
    .Z(_0410_));
 NAND2_X1 _1336_ (.A1(net44),
    .A2(_0155_),
    .ZN(_0411_));
 NAND3_X1 _1337_ (.A1(_0133_),
    .A2(_0925_),
    .A3(_0040_),
    .ZN(_0412_));
 AOI21_X1 _1338_ (.A(_0213_),
    .B1(_0411_),
    .B2(_0412_),
    .ZN(_0413_));
 MUX2_X1 _1339_ (.A(_0410_),
    .B(_0413_),
    .S(_0197_),
    .Z(_0414_));
 NAND2_X1 _1340_ (.A1(_0294_),
    .A2(_0414_),
    .ZN(_0415_));
 MUX2_X2 _1341_ (.A(_0109_),
    .B(_0229_),
    .S(_0274_),
    .Z(_0416_));
 AND2_X1 _1342_ (.A1(_0863_),
    .A2(_0040_),
    .ZN(_0417_));
 AOI22_X4 _1343_ (.A1(_0157_),
    .A2(net41),
    .B1(_0417_),
    .B2(_0244_),
    .ZN(_0418_));
 INV_X1 _1344_ (.A(_0418_),
    .ZN(_0419_));
 AOI22_X4 _1345_ (.A1(_0234_),
    .A2(_0416_),
    .B1(_0419_),
    .B2(_0251_),
    .ZN(_0420_));
 MUX2_X2 _1346_ (.A(_0070_),
    .B(_0236_),
    .S(_0274_),
    .Z(_0421_));
 AOI21_X2 _1347_ (.A(_0227_),
    .B1(_0125_),
    .B2(_0421_),
    .ZN(_0422_));
 OAI22_X4 _1348_ (.A1(_0125_),
    .A2(_0420_),
    .B1(_0422_),
    .B2(_0349_),
    .ZN(_0423_));
 MUX2_X1 _1349_ (.A(_0063_),
    .B(_0221_),
    .S(_0131_),
    .Z(_0424_));
 MUX2_X2 _1350_ (.A(_0051_),
    .B(_0248_),
    .S(_0131_),
    .Z(_0425_));
 MUX2_X1 _1351_ (.A(_0424_),
    .B(_0425_),
    .S(_0123_),
    .Z(_0426_));
 INV_X1 _1352_ (.A(_0426_),
    .ZN(_0427_));
 AOI21_X2 _1353_ (.A(_0884_),
    .B1(_0350_),
    .B2(_0427_),
    .ZN(_0428_));
 MUX2_X1 _1354_ (.A(_0200_),
    .B(_0362_),
    .S(_0131_),
    .Z(_0429_));
 AND2_X1 _1355_ (.A1(_0925_),
    .A2(_0394_),
    .ZN(_0430_));
 MUX2_X1 _1356_ (.A(_0429_),
    .B(_0430_),
    .S(_0021_),
    .Z(_0431_));
 MUX2_X1 _1357_ (.A(_0204_),
    .B(_0365_),
    .S(_0131_),
    .Z(_0432_));
 MUX2_X1 _1358_ (.A(_0107_),
    .B(_0091_),
    .S(_0154_),
    .Z(_0433_));
 MUX2_X1 _1359_ (.A(_0367_),
    .B(_0433_),
    .S(_0120_),
    .Z(_0434_));
 MUX2_X1 _1360_ (.A(_0432_),
    .B(_0434_),
    .S(_0167_),
    .Z(_0435_));
 MUX2_X1 _1361_ (.A(_0431_),
    .B(_0435_),
    .S(_0198_),
    .Z(_0436_));
 AOI22_X4 _1362_ (.A1(_0423_),
    .A2(_0428_),
    .B1(_0436_),
    .B2(_0192_),
    .ZN(_0437_));
 AOI22_X4 _1363_ (.A1(_0407_),
    .A2(_0415_),
    .B1(_0437_),
    .B2(_0129_),
    .ZN(net12));
 MUX2_X1 _1364_ (.A(_0111_),
    .B(_0110_),
    .S(net3),
    .Z(_0438_));
 MUX2_X1 _1365_ (.A(_0399_),
    .B(_0438_),
    .S(_0056_),
    .Z(_0439_));
 NOR2_X1 _1366_ (.A1(_0084_),
    .A2(_0914_),
    .ZN(_0440_));
 NOR3_X2 _1367_ (.A1(_0021_),
    .A2(_0031_),
    .A3(_0359_),
    .ZN(_0441_));
 OAI21_X4 _1368_ (.A(_0224_),
    .B1(_0440_),
    .B2(_0441_),
    .ZN(_0442_));
 NOR2_X2 _1369_ (.A1(_0821_),
    .A2(_0265_),
    .ZN(_0443_));
 NAND2_X2 _1370_ (.A1(_0914_),
    .A2(_0443_),
    .ZN(_0444_));
 AOI21_X2 _1371_ (.A(_0439_),
    .B1(_0442_),
    .B2(_0444_),
    .ZN(_0445_));
 MUX2_X1 _1372_ (.A(_0257_),
    .B(_0261_),
    .S(_0131_),
    .Z(_0446_));
 NAND2_X1 _1373_ (.A1(_0832_),
    .A2(_0914_),
    .ZN(_0447_));
 OR2_X1 _1374_ (.A1(_0832_),
    .A2(_0914_),
    .ZN(_0448_));
 OAI21_X2 _1375_ (.A(_0447_),
    .B1(_0448_),
    .B2(_0359_),
    .ZN(_0449_));
 AOI22_X4 _1376_ (.A1(_0031_),
    .A2(_0443_),
    .B1(_0224_),
    .B2(_0449_),
    .ZN(_0450_));
 OAI21_X2 _1377_ (.A(_0087_),
    .B1(_0446_),
    .B2(_0450_),
    .ZN(_0451_));
 NOR2_X2 _1378_ (.A1(_0059_),
    .A2(_0269_),
    .ZN(_0452_));
 MUX2_X1 _1379_ (.A(_0258_),
    .B(_0260_),
    .S(_0131_),
    .Z(_0453_));
 AOI21_X4 _1380_ (.A(_0452_),
    .B1(_0453_),
    .B2(_0059_),
    .ZN(_0454_));
 AOI211_X2 _1381_ (.A(_0451_),
    .B(_0445_),
    .C1(_0226_),
    .C2(_0454_),
    .ZN(_0455_));
 AND2_X1 _1382_ (.A1(_0385_),
    .A2(_0333_),
    .ZN(_0456_));
 AOI21_X1 _1383_ (.A(_0769_),
    .B1(_0245_),
    .B2(_0456_),
    .ZN(_0457_));
 INV_X1 _1384_ (.A(_0457_),
    .ZN(_0458_));
 MUX2_X1 _1385_ (.A(_0282_),
    .B(_0275_),
    .S(_0021_),
    .Z(_0459_));
 MUX2_X1 _1386_ (.A(_0285_),
    .B(_0289_),
    .S(_0207_),
    .Z(_0460_));
 MUX2_X1 _1387_ (.A(_0459_),
    .B(_0460_),
    .S(_0198_),
    .Z(_0461_));
 NOR3_X1 _1388_ (.A1(_0455_),
    .A2(_0458_),
    .A3(_0461_),
    .ZN(_0462_));
 MUX2_X1 _1389_ (.A(_0237_),
    .B(_0230_),
    .S(_0075_),
    .Z(_0463_));
 NOR3_X4 _1390_ (.A1(_0463_),
    .A2(_0226_),
    .A3(_0349_),
    .ZN(_0464_));
 OAI21_X4 _1391_ (.A(_0780_),
    .B1(_0884_),
    .B2(_0464_),
    .ZN(_0465_));
 NAND4_X1 _1392_ (.A1(_0224_),
    .A2(_0167_),
    .A3(_0914_),
    .A4(_0138_),
    .ZN(_0466_));
 OAI221_X2 _1393_ (.A(_0466_),
    .B1(_0137_),
    .B2(_0077_),
    .C1(_0894_),
    .C2(_0138_),
    .ZN(_0467_));
 AOI21_X1 _1394_ (.A(_0233_),
    .B1(_0246_),
    .B2(_0467_),
    .ZN(_0468_));
 MUX2_X1 _1395_ (.A(_0249_),
    .B(_0222_),
    .S(_0075_),
    .Z(_0469_));
 INV_X1 _1396_ (.A(_0469_),
    .ZN(_0470_));
 AOI21_X2 _1397_ (.A(_0468_),
    .B1(_0470_),
    .B2(_0350_),
    .ZN(_0471_));
 OAI221_X2 _1398_ (.A(_0465_),
    .B1(_0455_),
    .B2(_0458_),
    .C1(_0471_),
    .C2(_0195_),
    .ZN(_0472_));
 BUF_X4 _1399_ (.A(_0197_),
    .Z(_0473_));
 OAI21_X1 _1400_ (.A(_0465_),
    .B1(_0471_),
    .B2(_0306_),
    .ZN(_0474_));
 CLKBUF_X3 _1401_ (.A(_0224_),
    .Z(_0475_));
 NAND2_X1 _1402_ (.A1(_0213_),
    .A2(_0211_),
    .ZN(_0476_));
 OR2_X1 _1403_ (.A1(_0213_),
    .A2(_0203_),
    .ZN(_0477_));
 NAND3_X1 _1404_ (.A1(_0475_),
    .A2(_0476_),
    .A3(_0477_),
    .ZN(_0478_));
 MUX2_X1 _1405_ (.A(_0111_),
    .B(_0110_),
    .S(_0148_),
    .Z(_0479_));
 MUX2_X1 _1406_ (.A(_0433_),
    .B(_0479_),
    .S(_0202_),
    .Z(_0480_));
 MUX2_X1 _1407_ (.A(_0206_),
    .B(_0480_),
    .S(_0168_),
    .Z(_0481_));
 NAND2_X1 _1408_ (.A1(_0190_),
    .A2(_0481_),
    .ZN(_0482_));
 AND2_X1 _1409_ (.A1(_0478_),
    .A2(_0482_),
    .ZN(_0483_));
 AOI221_X2 _1410_ (.A(_0462_),
    .B1(_0473_),
    .B2(_0472_),
    .C1(_0474_),
    .C2(_0483_),
    .ZN(net13));
 MUX2_X1 _1411_ (.A(_0308_),
    .B(_0315_),
    .S(_0123_),
    .Z(_0484_));
 NOR3_X2 _1412_ (.A1(_0349_),
    .A2(_0256_),
    .A3(_0484_),
    .ZN(_0485_));
 AOI21_X2 _1413_ (.A(_0234_),
    .B1(_0314_),
    .B2(_0467_),
    .ZN(_0486_));
 MUX2_X1 _1414_ (.A(_0309_),
    .B(_0317_),
    .S(_0075_),
    .Z(_0487_));
 NOR3_X2 _1415_ (.A1(_0349_),
    .A2(_0227_),
    .A3(_0487_),
    .ZN(_0488_));
 NOR4_X4 _1416_ (.A1(_0884_),
    .A2(_0485_),
    .A3(_0486_),
    .A4(_0488_),
    .ZN(_0489_));
 MUX2_X2 _1417_ (.A(_0298_),
    .B(_0303_),
    .S(_0021_),
    .Z(_0490_));
 MUX2_X1 _1418_ (.A(_0108_),
    .B(_0107_),
    .S(_0148_),
    .Z(_0491_));
 MUX2_X1 _1419_ (.A(_0479_),
    .B(_0491_),
    .S(_0103_),
    .Z(_0492_));
 MUX2_X1 _1420_ (.A(_0300_),
    .B(_0492_),
    .S(_0168_),
    .Z(_0493_));
 MUX2_X1 _1421_ (.A(_0490_),
    .B(_0493_),
    .S(_0170_),
    .Z(_0494_));
 MUX2_X2 _1422_ (.A(_0341_),
    .B(_0338_),
    .S(_0124_),
    .Z(_0495_));
 NOR2_X2 _1423_ (.A1(_0256_),
    .A2(_0495_),
    .ZN(_0496_));
 MUX2_X1 _1424_ (.A(_0108_),
    .B(_0107_),
    .S(_0092_),
    .Z(_0497_));
 MUX2_X2 _1425_ (.A(_0438_),
    .B(_0497_),
    .S(_0120_),
    .Z(_0498_));
 AOI21_X2 _1426_ (.A(_0498_),
    .B1(_0442_),
    .B2(_0444_),
    .ZN(_0499_));
 NOR2_X2 _1427_ (.A1(_0344_),
    .A2(_0450_),
    .ZN(_0500_));
 NOR4_X2 _1428_ (.A1(_0145_),
    .A2(_0496_),
    .A3(_0499_),
    .A4(_0500_),
    .ZN(_0501_));
 NOR2_X2 _1429_ (.A1(_0133_),
    .A2(_0313_),
    .ZN(_0502_));
 AOI21_X1 _1430_ (.A(_0780_),
    .B1(_0502_),
    .B2(_0456_),
    .ZN(_0503_));
 INV_X1 _1431_ (.A(_0503_),
    .ZN(_0504_));
 MUX2_X1 _1432_ (.A(_0156_),
    .B(_0273_),
    .S(_0103_),
    .Z(_0505_));
 MUX2_X1 _1433_ (.A(_0323_),
    .B(_0505_),
    .S(_0021_),
    .Z(_0506_));
 MUX2_X1 _1434_ (.A(_0324_),
    .B(_0326_),
    .S(_0167_),
    .Z(_0507_));
 MUX2_X1 _1435_ (.A(_0506_),
    .B(_0507_),
    .S(_0190_),
    .Z(_0508_));
 OAI33_X1 _1436_ (.A1(_0489_),
    .A2(_0196_),
    .A3(_0494_),
    .B1(_0501_),
    .B2(_0504_),
    .B3(_0508_),
    .ZN(_0509_));
 OAI22_X2 _1437_ (.A1(_0196_),
    .A2(_0489_),
    .B1(_0501_),
    .B2(_0504_),
    .ZN(_0510_));
 BUF_X4 _1438_ (.A(_0197_),
    .Z(_0511_));
 AOI21_X2 _1439_ (.A(_0509_),
    .B1(_0510_),
    .B2(_0511_),
    .ZN(net14));
 MUX2_X1 _1440_ (.A(_0388_),
    .B(_0379_),
    .S(net105),
    .Z(_0512_));
 NAND3_X1 _1441_ (.A1(net44),
    .A2(_0135_),
    .A3(_0266_),
    .ZN(_0513_));
 MUX2_X1 _1442_ (.A(_0340_),
    .B(_0337_),
    .S(_0123_),
    .Z(_0514_));
 NAND2_X1 _1443_ (.A1(_0198_),
    .A2(_0133_),
    .ZN(_0515_));
 OAI22_X2 _1444_ (.A1(_0512_),
    .A2(_0513_),
    .B1(_0514_),
    .B2(_0515_),
    .ZN(_0516_));
 MUX2_X1 _1445_ (.A(_0071_),
    .B(_0111_),
    .S(net3),
    .Z(_0517_));
 MUX2_X1 _1446_ (.A(_0497_),
    .B(_0517_),
    .S(net4),
    .Z(_0518_));
 AOI21_X1 _1447_ (.A(_0518_),
    .B1(_0442_),
    .B2(_0444_),
    .ZN(_0519_));
 MUX2_X1 _1448_ (.A(_0343_),
    .B(_0380_),
    .S(_0157_),
    .Z(_0520_));
 OAI21_X1 _1449_ (.A(_0088_),
    .B1(_0450_),
    .B2(_0520_),
    .ZN(_0521_));
 NOR3_X2 _1450_ (.A1(_0516_),
    .A2(_0519_),
    .A3(_0521_),
    .ZN(_0522_));
 NAND2_X1 _1451_ (.A1(_0244_),
    .A2(_0134_),
    .ZN(_0523_));
 OAI21_X1 _1452_ (.A(_0038_),
    .B1(_0140_),
    .B2(_0136_),
    .ZN(_0524_));
 OAI21_X2 _1453_ (.A(_0306_),
    .B1(_0523_),
    .B2(_0524_),
    .ZN(_0525_));
 AND2_X4 _1454_ (.A1(_0089_),
    .A2(_0081_),
    .ZN(_0526_));
 INV_X1 _1455_ (.A(_0456_),
    .ZN(_0527_));
 OAI21_X1 _1456_ (.A(_0335_),
    .B1(_0800_),
    .B2(_0527_),
    .ZN(_0528_));
 MUX2_X1 _1457_ (.A(_0302_),
    .B(_0362_),
    .S(_0183_),
    .Z(_0529_));
 MUX2_X1 _1458_ (.A(_0529_),
    .B(_0366_),
    .S(_0179_),
    .Z(_0530_));
 MUX2_X1 _1459_ (.A(_0071_),
    .B(_0111_),
    .S(_0161_),
    .Z(_0531_));
 MUX2_X1 _1460_ (.A(_0491_),
    .B(_0531_),
    .S(_0152_),
    .Z(_0532_));
 MUX2_X1 _1461_ (.A(_0368_),
    .B(_0532_),
    .S(_0179_),
    .Z(_0533_));
 MUX2_X1 _1462_ (.A(_0530_),
    .B(_0533_),
    .S(_0190_),
    .Z(_0534_));
 OAI33_X1 _1463_ (.A1(_0171_),
    .A2(_0522_),
    .A3(_0525_),
    .B1(_0526_),
    .B2(_0528_),
    .B3(_0534_),
    .ZN(_0535_));
 OAI22_X2 _1464_ (.A1(_0522_),
    .A2(_0525_),
    .B1(_0526_),
    .B2(_0528_),
    .ZN(_0536_));
 AOI21_X2 _1465_ (.A(_0535_),
    .B1(_0536_),
    .B2(_0511_),
    .ZN(net15));
 NAND4_X1 _1466_ (.A1(_0135_),
    .A2(_0266_),
    .A3(_0124_),
    .A4(_0418_),
    .ZN(_0537_));
 OAI221_X2 _1467_ (.A(_0537_),
    .B1(_0450_),
    .B2(_0424_),
    .C1(_0267_),
    .C2(_0425_),
    .ZN(_0538_));
 AOI21_X2 _1468_ (.A(_0421_),
    .B1(_0442_),
    .B2(_0444_),
    .ZN(_0539_));
 NOR3_X4 _1469_ (.A1(_0145_),
    .A2(_0538_),
    .A3(_0539_),
    .ZN(_0540_));
 NAND2_X1 _1470_ (.A1(_0394_),
    .A2(_0456_),
    .ZN(_0541_));
 NAND2_X1 _1471_ (.A1(_0780_),
    .A2(_0541_),
    .ZN(_0542_));
 MUX2_X1 _1472_ (.A(_0429_),
    .B(_0432_),
    .S(_0207_),
    .Z(_0543_));
 MUX2_X1 _1473_ (.A(_0068_),
    .B(_0108_),
    .S(_0161_),
    .Z(_0544_));
 MUX2_X1 _1474_ (.A(_0531_),
    .B(_0544_),
    .S(_0157_),
    .Z(_0545_));
 MUX2_X1 _1475_ (.A(_0434_),
    .B(_0545_),
    .S(_0207_),
    .Z(_0546_));
 MUX2_X1 _1476_ (.A(_0543_),
    .B(_0546_),
    .S(_0198_),
    .Z(_0547_));
 NOR3_X1 _1477_ (.A1(_0540_),
    .A2(_0542_),
    .A3(_0547_),
    .ZN(_0548_));
 MUX2_X1 _1478_ (.A(_0380_),
    .B(_0517_),
    .S(net105),
    .Z(_0549_));
 MUX2_X1 _1479_ (.A(_0068_),
    .B(_0108_),
    .S(net56),
    .Z(_0550_));
 MUX2_X1 _1480_ (.A(_0399_),
    .B(_0550_),
    .S(net105),
    .Z(_0551_));
 MUX2_X2 _1481_ (.A(_0549_),
    .B(_0551_),
    .S(_0103_),
    .Z(_0552_));
 NOR3_X4 _1482_ (.A1(_0348_),
    .A2(_0226_),
    .A3(_0552_),
    .ZN(_0553_));
 MUX2_X2 _1483_ (.A(_0262_),
    .B(_0512_),
    .S(_0274_),
    .Z(_0554_));
 NOR3_X2 _1484_ (.A1(_0348_),
    .A2(_0080_),
    .A3(_0554_),
    .ZN(_0555_));
 AOI21_X2 _1485_ (.A(_0233_),
    .B1(_0395_),
    .B2(_0467_),
    .ZN(_0556_));
 NOR4_X4 _1486_ (.A1(_0555_),
    .A2(_0553_),
    .A3(_0884_),
    .A4(_0556_),
    .ZN(_0557_));
 OAI22_X2 _1487_ (.A1(_0557_),
    .A2(_0128_),
    .B1(_0540_),
    .B2(_0542_),
    .ZN(_0558_));
 NOR2_X1 _1488_ (.A1(_0128_),
    .A2(_0557_),
    .ZN(_0559_));
 MUX2_X1 _1489_ (.A(_0403_),
    .B(_0408_),
    .S(_0207_),
    .Z(_0560_));
 AND2_X1 _1490_ (.A1(_0170_),
    .A2(_0560_),
    .ZN(_0561_));
 NAND2_X1 _1491_ (.A1(_0411_),
    .A2(_0412_),
    .ZN(_0562_));
 MUX2_X1 _1492_ (.A(_0562_),
    .B(_0404_),
    .S(_0188_),
    .Z(_0563_));
 AOI21_X2 _1493_ (.A(_0561_),
    .B1(_0563_),
    .B2(_0475_),
    .ZN(_0564_));
 AOI221_X2 _1494_ (.A(_0548_),
    .B1(_0473_),
    .B2(_0558_),
    .C1(_0559_),
    .C2(_0564_),
    .ZN(net16));
 NAND2_X1 _1495_ (.A1(_0374_),
    .A2(_0333_),
    .ZN(_0565_));
 OAI21_X1 _1496_ (.A(_0780_),
    .B1(_0211_),
    .B2(_0565_),
    .ZN(_0566_));
 MUX2_X1 _1497_ (.A(_0237_),
    .B(_0222_),
    .S(_0123_),
    .Z(_0567_));
 MUX2_X2 _1498_ (.A(_0250_),
    .B(_0567_),
    .S(_0080_),
    .Z(_0568_));
 MUX2_X1 _1499_ (.A(_0072_),
    .B(_0071_),
    .S(_0148_),
    .Z(_0569_));
 MUX2_X1 _1500_ (.A(_0544_),
    .B(_0569_),
    .S(_0202_),
    .Z(_0570_));
 MUX2_X1 _1501_ (.A(_0480_),
    .B(_0570_),
    .S(_0207_),
    .Z(_0571_));
 MUX2_X1 _1502_ (.A(_0208_),
    .B(_0571_),
    .S(_0198_),
    .Z(_0572_));
 AOI221_X2 _1503_ (.A(_0566_),
    .B1(_0568_),
    .B2(_0088_),
    .C1(_0371_),
    .C2(_0572_),
    .ZN(_0573_));
 MUX2_X1 _1504_ (.A(_0072_),
    .B(_0071_),
    .S(net68),
    .Z(_0574_));
 MUX2_X1 _1505_ (.A(_0438_),
    .B(_0574_),
    .S(_0059_),
    .Z(_0575_));
 MUX2_X1 _1506_ (.A(_0551_),
    .B(_0575_),
    .S(net44),
    .Z(_0576_));
 MUX2_X1 _1507_ (.A(_0263_),
    .B(_0576_),
    .S(_0219_),
    .Z(_0577_));
 NAND2_X1 _1508_ (.A1(_0255_),
    .A2(_0577_),
    .ZN(_0578_));
 NAND2_X1 _1509_ (.A1(_0244_),
    .A2(_0210_),
    .ZN(_0579_));
 INV_X1 _1510_ (.A(_0268_),
    .ZN(_0580_));
 OAI21_X2 _1511_ (.A(_0579_),
    .B1(_0580_),
    .B2(_0133_),
    .ZN(_0581_));
 NAND2_X2 _1512_ (.A1(_0143_),
    .A2(_0349_),
    .ZN(_0582_));
 NOR2_X1 _1513_ (.A1(_0141_),
    .A2(_0582_),
    .ZN(_0583_));
 NAND2_X1 _1514_ (.A1(_0190_),
    .A2(_0286_),
    .ZN(_0584_));
 OAI21_X2 _1515_ (.A(_0584_),
    .B1(_0277_),
    .B2(_0199_),
    .ZN(_0585_));
 AOI221_X2 _1516_ (.A(_0128_),
    .B1(_0581_),
    .B2(_0583_),
    .C1(_0585_),
    .C2(_0371_),
    .ZN(_0586_));
 AOI21_X2 _1517_ (.A(_0573_),
    .B1(_0578_),
    .B2(_0586_),
    .ZN(net17));
 MUX2_X1 _1518_ (.A(_0069_),
    .B(_0068_),
    .S(net68),
    .Z(_0587_));
 MUX2_X2 _1519_ (.A(_0574_),
    .B(_0587_),
    .S(_0120_),
    .Z(_0588_));
 AOI22_X2 _1520_ (.A1(_0251_),
    .A2(net65),
    .B1(_0588_),
    .B2(_0233_),
    .ZN(_0589_));
 AOI21_X1 _1521_ (.A(_0226_),
    .B1(_0352_),
    .B2(_0498_),
    .ZN(_0590_));
 OAI22_X2 _1522_ (.A1(_0125_),
    .A2(_0589_),
    .B1(_0590_),
    .B2(_0349_),
    .ZN(_0591_));
 AOI21_X1 _1523_ (.A(_0884_),
    .B1(_0345_),
    .B2(_0350_),
    .ZN(_0592_));
 MUX2_X1 _1524_ (.A(_0325_),
    .B(_0332_),
    .S(_0224_),
    .Z(_0593_));
 AOI221_X2 _1525_ (.A(_0335_),
    .B1(_0591_),
    .B2(_0592_),
    .C1(_0593_),
    .C2(_0371_),
    .ZN(_0594_));
 MUX2_X1 _1526_ (.A(_0069_),
    .B(_0068_),
    .S(_0148_),
    .Z(_0595_));
 MUX2_X1 _1527_ (.A(_0569_),
    .B(_0595_),
    .S(_0709_),
    .Z(_0596_));
 MUX2_X1 _1528_ (.A(_0492_),
    .B(_0596_),
    .S(_0188_),
    .Z(_0597_));
 MUX2_X1 _1529_ (.A(_0301_),
    .B(_0597_),
    .S(_0294_),
    .Z(_0598_));
 NAND2_X1 _1530_ (.A1(_0192_),
    .A2(_0598_),
    .ZN(_0599_));
 MUX2_X1 _1531_ (.A(_0310_),
    .B(_0316_),
    .S(_0226_),
    .Z(_0600_));
 AOI221_X2 _1532_ (.A(_0306_),
    .B1(_0303_),
    .B2(_0392_),
    .C1(net48),
    .C2(_0089_),
    .ZN(_0601_));
 AOI21_X2 _1533_ (.A(_0594_),
    .B1(_0601_),
    .B2(_0599_),
    .ZN(net18));
 OR3_X1 _1534_ (.A1(_0582_),
    .A2(_0538_),
    .A3(_0539_),
    .ZN(_0602_));
 AND2_X1 _1535_ (.A1(_0385_),
    .A2(_0085_),
    .ZN(_0603_));
 MUX2_X1 _1536_ (.A(_0101_),
    .B(_0117_),
    .S(net54),
    .Z(_0604_));
 MUX2_X1 _1537_ (.A(_0100_),
    .B(_0604_),
    .S(_0132_),
    .Z(_0605_));
 MUX2_X1 _1538_ (.A(_0093_),
    .B(_0240_),
    .S(_0274_),
    .Z(_0606_));
 MUX2_X1 _1539_ (.A(_0605_),
    .B(_0606_),
    .S(_0226_),
    .Z(_0607_));
 MUX2_X1 _1540_ (.A(_0118_),
    .B(_0094_),
    .S(net54),
    .Z(_0608_));
 MUX2_X1 _1541_ (.A(_0116_),
    .B(_0608_),
    .S(_0132_),
    .Z(_0609_));
 MUX2_X1 _1542_ (.A(_0416_),
    .B(_0609_),
    .S(_0105_),
    .Z(_0610_));
 MUX2_X1 _1543_ (.A(_0607_),
    .B(_0610_),
    .S(_0125_),
    .Z(_0611_));
 AOI221_X2 _1544_ (.A(_0306_),
    .B1(_0603_),
    .B2(_0394_),
    .C1(_0611_),
    .C2(_0089_),
    .ZN(_0612_));
 MUX2_X1 _1545_ (.A(_0118_),
    .B(_0094_),
    .S(_0172_),
    .Z(_0613_));
 MUX2_X1 _1546_ (.A(_0181_),
    .B(_0613_),
    .S(_0132_),
    .Z(_0614_));
 NOR2_X1 _1547_ (.A1(_0188_),
    .A2(_0614_),
    .ZN(_0615_));
 MUX2_X1 _1548_ (.A(_0101_),
    .B(_0117_),
    .S(_0739_),
    .Z(_0616_));
 MUX2_X1 _1549_ (.A(_0185_),
    .B(_0616_),
    .S(_0132_),
    .Z(_0617_));
 NOR2_X1 _1550_ (.A1(_0213_),
    .A2(_0617_),
    .ZN(_0618_));
 NOR3_X1 _1551_ (.A1(_0475_),
    .A2(_0615_),
    .A3(_0618_),
    .ZN(_0619_));
 MUX2_X1 _1552_ (.A(_0176_),
    .B(_0291_),
    .S(_0132_),
    .Z(_0620_));
 MUX2_X1 _1553_ (.A(_0409_),
    .B(_0620_),
    .S(_0179_),
    .Z(_0621_));
 AOI21_X1 _1554_ (.A(_0619_),
    .B1(_0621_),
    .B2(_0475_),
    .ZN(_0622_));
 MUX2_X1 _1555_ (.A(_0564_),
    .B(_0622_),
    .S(_0192_),
    .Z(_0623_));
 AOI21_X2 _1556_ (.A(_0336_),
    .B1(_0146_),
    .B2(_0394_),
    .ZN(_0624_));
 AOI22_X4 _1557_ (.A1(_0602_),
    .A2(_0612_),
    .B1(_0623_),
    .B2(_0624_),
    .ZN(net19));
 AOI21_X2 _1558_ (.A(_0780_),
    .B1(_0307_),
    .B2(_0382_),
    .ZN(_0625_));
 AND2_X1 _1559_ (.A1(_0352_),
    .A2(_0518_),
    .ZN(_0626_));
 MUX2_X1 _1560_ (.A(_0064_),
    .B(_0072_),
    .S(net68),
    .Z(_0627_));
 MUX2_X1 _1561_ (.A(_0587_),
    .B(_0627_),
    .S(_0120_),
    .Z(_0628_));
 AOI21_X2 _1562_ (.A(_0626_),
    .B1(_0628_),
    .B2(_0218_),
    .ZN(_0629_));
 NAND2_X2 _1563_ (.A1(_0088_),
    .A2(_0256_),
    .ZN(_0630_));
 NAND2_X1 _1564_ (.A1(_0125_),
    .A2(_0384_),
    .ZN(_0631_));
 AND2_X1 _1565_ (.A1(_0390_),
    .A2(_0631_),
    .ZN(_0632_));
 NAND2_X1 _1566_ (.A1(_0256_),
    .A2(_0037_),
    .ZN(_0633_));
 OAI221_X2 _1567_ (.A(_0625_),
    .B1(_0629_),
    .B2(_0630_),
    .C1(_0632_),
    .C2(_0633_),
    .ZN(_0634_));
 AND2_X1 _1568_ (.A1(_0190_),
    .A2(_0373_),
    .ZN(_0635_));
 AND2_X1 _1569_ (.A1(_0158_),
    .A2(_0214_),
    .ZN(_0636_));
 AND3_X1 _1570_ (.A1(_0135_),
    .A2(_0266_),
    .A3(_0217_),
    .ZN(_0637_));
 NAND2_X1 _1571_ (.A1(_0047_),
    .A2(_0637_),
    .ZN(_0638_));
 OAI21_X1 _1572_ (.A(_0067_),
    .B1(_0140_),
    .B2(_0136_),
    .ZN(_0639_));
 AOI21_X1 _1573_ (.A(_0145_),
    .B1(_0638_),
    .B2(_0639_),
    .ZN(_0640_));
 AND3_X1 _1574_ (.A1(_0360_),
    .A2(_0361_),
    .A3(_0363_),
    .ZN(_0641_));
 OR2_X1 _1575_ (.A1(_0145_),
    .A2(_0450_),
    .ZN(_0642_));
 INV_X1 _1576_ (.A(_0057_),
    .ZN(_0643_));
 OAI221_X2 _1577_ (.A(_0780_),
    .B1(_0278_),
    .B2(_0641_),
    .C1(_0642_),
    .C2(_0643_),
    .ZN(_0644_));
 MUX2_X1 _1578_ (.A(_0064_),
    .B(_0072_),
    .S(_0161_),
    .Z(_0645_));
 MUX2_X1 _1579_ (.A(_0595_),
    .B(_0645_),
    .S(_0152_),
    .Z(_0646_));
 MUX2_X1 _1580_ (.A(_0532_),
    .B(_0646_),
    .S(_0168_),
    .Z(_0647_));
 MUX2_X1 _1581_ (.A(_0369_),
    .B(_0647_),
    .S(_0190_),
    .Z(_0648_));
 OAI33_X1 _1582_ (.A1(_0634_),
    .A2(_0635_),
    .A3(_0636_),
    .B1(_0640_),
    .B2(_0644_),
    .B3(_0648_),
    .ZN(_0649_));
 OAI21_X1 _1583_ (.A(_0634_),
    .B1(_0640_),
    .B2(_0644_),
    .ZN(_0650_));
 AOI21_X2 _1584_ (.A(_0649_),
    .B1(_0650_),
    .B2(_0511_),
    .ZN(net20));
 NOR3_X1 _1585_ (.A1(_0080_),
    .A2(_0124_),
    .A3(_0418_),
    .ZN(_0651_));
 AOI21_X2 _1586_ (.A(_0651_),
    .B1(_0080_),
    .B2(_0426_),
    .ZN(_0652_));
 OAI21_X2 _1587_ (.A(_0780_),
    .B1(_0145_),
    .B2(_0652_),
    .ZN(_0653_));
 MUX2_X1 _1588_ (.A(_0061_),
    .B(_0069_),
    .S(_0161_),
    .Z(_0654_));
 MUX2_X1 _1589_ (.A(_0645_),
    .B(_0654_),
    .S(_0157_),
    .Z(_0655_));
 MUX2_X1 _1590_ (.A(_0545_),
    .B(_0655_),
    .S(_0207_),
    .Z(_0656_));
 MUX2_X1 _1591_ (.A(_0435_),
    .B(_0656_),
    .S(_0198_),
    .Z(_0657_));
 AOI221_X2 _1592_ (.A(_0653_),
    .B1(_0431_),
    .B2(_0333_),
    .C1(_0371_),
    .C2(_0657_),
    .ZN(_0658_));
 MUX2_X1 _1593_ (.A(_0061_),
    .B(_0069_),
    .S(net54),
    .Z(_0659_));
 MUX2_X1 _1594_ (.A(_0627_),
    .B(_0659_),
    .S(_0103_),
    .Z(_0660_));
 MUX2_X1 _1595_ (.A(_0517_),
    .B(_0550_),
    .S(net42),
    .Z(_0661_));
 MUX2_X1 _1596_ (.A(_0660_),
    .B(_0661_),
    .S(_0124_),
    .Z(_0662_));
 MUX2_X1 _1597_ (.A(_0397_),
    .B(_0662_),
    .S(_0234_),
    .Z(_0663_));
 AOI221_X2 _1598_ (.A(_0128_),
    .B1(_0307_),
    .B2(_0401_),
    .C1(_0663_),
    .C2(_0312_),
    .ZN(_0664_));
 MUX2_X1 _1599_ (.A(_0405_),
    .B(_0413_),
    .S(_0475_),
    .Z(_0665_));
 NAND2_X1 _1600_ (.A1(_0192_),
    .A2(_0665_),
    .ZN(_0666_));
 AOI21_X2 _1601_ (.A(_0658_),
    .B1(_0664_),
    .B2(_0666_),
    .ZN(net21));
 NAND3_X1 _1602_ (.A1(_0333_),
    .A2(_0476_),
    .A3(_0477_),
    .ZN(_0667_));
 AND3_X1 _1603_ (.A1(_0226_),
    .A2(_0075_),
    .A3(_0246_),
    .ZN(_0668_));
 AOI21_X2 _1604_ (.A(_0668_),
    .B1(_0469_),
    .B2(_0080_),
    .ZN(_0669_));
 OAI21_X1 _1605_ (.A(_0667_),
    .B1(_0669_),
    .B2(_0145_),
    .ZN(_0670_));
 NAND2_X1 _1606_ (.A1(_0129_),
    .A2(_0670_),
    .ZN(_0671_));
 NOR3_X1 _1607_ (.A1(_0234_),
    .A2(_0227_),
    .A3(_0454_),
    .ZN(_0672_));
 MUX2_X1 _1608_ (.A(_0065_),
    .B(_0064_),
    .S(net54),
    .Z(_0673_));
 MUX2_X1 _1609_ (.A(_0659_),
    .B(_0673_),
    .S(_0152_),
    .Z(_0674_));
 MUX2_X1 _1610_ (.A(_0550_),
    .B(_0574_),
    .S(_0183_),
    .Z(_0675_));
 MUX2_X1 _1611_ (.A(_0674_),
    .B(_0675_),
    .S(_0352_),
    .Z(_0676_));
 NAND2_X1 _1612_ (.A1(_0219_),
    .A2(_0676_),
    .ZN(_0678_));
 MUX2_X1 _1613_ (.A(_0439_),
    .B(_0446_),
    .S(_0352_),
    .Z(_0679_));
 NAND2_X1 _1614_ (.A1(_0227_),
    .A2(_0679_),
    .ZN(_0680_));
 AOI21_X1 _1615_ (.A(_0349_),
    .B1(_0678_),
    .B2(_0680_),
    .ZN(_0681_));
 OAI21_X2 _1616_ (.A(_0143_),
    .B1(_0672_),
    .B2(_0681_),
    .ZN(_0682_));
 AND2_X1 _1617_ (.A1(_0224_),
    .A2(_0385_),
    .ZN(_0683_));
 AOI22_X2 _1618_ (.A1(_0170_),
    .A2(_0459_),
    .B1(_0683_),
    .B2(_0245_),
    .ZN(_0684_));
 NOR2_X1 _1619_ (.A1(_0128_),
    .A2(_0684_),
    .ZN(_0685_));
 MUX2_X1 _1620_ (.A(_0065_),
    .B(_0064_),
    .S(_0148_),
    .Z(_0686_));
 MUX2_X1 _1621_ (.A(_0654_),
    .B(_0686_),
    .S(_0152_),
    .Z(_0687_));
 MUX2_X1 _1622_ (.A(_0570_),
    .B(_0687_),
    .S(_0168_),
    .Z(_0689_));
 MUX2_X1 _1623_ (.A(_0481_),
    .B(_0689_),
    .S(_0199_),
    .Z(_0690_));
 AOI21_X2 _1624_ (.A(_0685_),
    .B1(_0690_),
    .B2(_0336_),
    .ZN(_0691_));
 OAI221_X2 _1625_ (.A(_0671_),
    .B1(_0682_),
    .B2(_0129_),
    .C1(_0511_),
    .C2(_0691_),
    .ZN(net22));
 NOR3_X1 _1626_ (.A1(_0077_),
    .A2(_0313_),
    .A3(_0265_),
    .ZN(_0692_));
 AOI21_X2 _1627_ (.A(_0692_),
    .B1(_0506_),
    .B2(_0170_),
    .ZN(_0693_));
 NOR2_X1 _1628_ (.A1(_0336_),
    .A2(_0693_),
    .ZN(_0694_));
 MUX2_X1 _1629_ (.A(_0062_),
    .B(_0061_),
    .S(_0172_),
    .Z(_0695_));
 MUX2_X1 _1630_ (.A(_0686_),
    .B(_0695_),
    .S(_0709_),
    .Z(_0696_));
 MUX2_X1 _1631_ (.A(_0596_),
    .B(_0696_),
    .S(_0179_),
    .Z(_0697_));
 MUX2_X1 _1632_ (.A(_0493_),
    .B(_0697_),
    .S(_0199_),
    .Z(_0699_));
 AOI21_X2 _1633_ (.A(_0694_),
    .B1(_0699_),
    .B2(_0129_),
    .ZN(_0700_));
 MUX2_X1 _1634_ (.A(_0062_),
    .B(_0061_),
    .S(net54),
    .Z(_0701_));
 MUX2_X1 _1635_ (.A(_0673_),
    .B(_0701_),
    .S(_0202_),
    .Z(_0702_));
 MUX2_X1 _1636_ (.A(_0498_),
    .B(_0702_),
    .S(_0105_),
    .Z(_0703_));
 MUX2_X1 _1637_ (.A(_0344_),
    .B(_0588_),
    .S(_0105_),
    .Z(_0704_));
 MUX2_X1 _1638_ (.A(_0703_),
    .B(_0704_),
    .S(_0352_),
    .Z(_0705_));
 AND2_X1 _1639_ (.A1(_0219_),
    .A2(_0495_),
    .ZN(_0706_));
 MUX2_X1 _1640_ (.A(_0705_),
    .B(_0706_),
    .S(_0349_),
    .Z(_0707_));
 AOI21_X4 _1641_ (.A(_0336_),
    .B1(_0143_),
    .B2(_0707_),
    .ZN(_0708_));
 AND2_X1 _1642_ (.A1(_0217_),
    .A2(_0314_),
    .ZN(_0710_));
 MUX2_X1 _1643_ (.A(_0484_),
    .B(_0710_),
    .S(_0227_),
    .Z(_0711_));
 AOI221_X2 _1644_ (.A(_0195_),
    .B1(_0333_),
    .B2(_0490_),
    .C1(net51),
    .C2(_0089_),
    .ZN(_0712_));
 OAI22_X4 _1645_ (.A1(_0511_),
    .A2(_0700_),
    .B1(_0708_),
    .B2(_0712_),
    .ZN(net23));
 AND3_X1 _1646_ (.A1(_0475_),
    .A2(_0134_),
    .A3(_0385_),
    .ZN(_0713_));
 AOI21_X2 _1647_ (.A(_0713_),
    .B1(_0530_),
    .B2(_0294_),
    .ZN(_0714_));
 NAND2_X1 _1648_ (.A1(_0473_),
    .A2(_0714_),
    .ZN(_0715_));
 MUX2_X1 _1649_ (.A(_0052_),
    .B(_0065_),
    .S(_0150_),
    .Z(_0716_));
 MUX2_X1 _1650_ (.A(_0695_),
    .B(_0716_),
    .S(_0709_),
    .Z(_0717_));
 MUX2_X1 _1651_ (.A(_0646_),
    .B(_0717_),
    .S(_0374_),
    .Z(_0718_));
 MUX2_X1 _1652_ (.A(_0533_),
    .B(_0718_),
    .S(_0294_),
    .Z(_0719_));
 OAI21_X2 _1653_ (.A(_0715_),
    .B1(_0719_),
    .B2(_0511_),
    .ZN(_0720_));
 NOR2_X4 _1654_ (.A1(_0144_),
    .A2(_0226_),
    .ZN(_0721_));
 AOI21_X2 _1655_ (.A(_0196_),
    .B1(net40),
    .B2(_0721_),
    .ZN(_0722_));
 NOR2_X2 _1656_ (.A1(_0352_),
    .A2(_0387_),
    .ZN(_0723_));
 MUX2_X1 _1657_ (.A(_0512_),
    .B(_0514_),
    .S(_0133_),
    .Z(_0724_));
 AND2_X1 _1658_ (.A1(_0219_),
    .A2(_0724_),
    .ZN(_0725_));
 OAI21_X2 _1659_ (.A(_0038_),
    .B1(_0723_),
    .B2(_0725_),
    .ZN(_0726_));
 MUX2_X1 _1660_ (.A(_0052_),
    .B(_0065_),
    .S(net54),
    .Z(_0727_));
 MUX2_X1 _1661_ (.A(_0701_),
    .B(_0727_),
    .S(_0202_),
    .Z(_0728_));
 MUX2_X1 _1662_ (.A(_0518_),
    .B(_0728_),
    .S(_0079_),
    .Z(_0730_));
 MUX2_X1 _1663_ (.A(_0520_),
    .B(_0628_),
    .S(_0105_),
    .Z(_0731_));
 MUX2_X1 _1664_ (.A(_0730_),
    .B(_0731_),
    .S(_0352_),
    .Z(_0732_));
 AOI221_X2 _1665_ (.A(_0335_),
    .B1(_0159_),
    .B2(_0085_),
    .C1(_0732_),
    .C2(_0089_),
    .ZN(_0733_));
 AOI22_X4 _1666_ (.A1(_0720_),
    .A2(_0722_),
    .B1(_0726_),
    .B2(_0733_),
    .ZN(net24));
 AOI22_X2 _1667_ (.A1(_0190_),
    .A2(_0543_),
    .B1(_0683_),
    .B2(_0394_),
    .ZN(_0734_));
 NAND2_X1 _1668_ (.A1(_0473_),
    .A2(_0734_),
    .ZN(_0735_));
 MUX2_X1 _1669_ (.A(_0048_),
    .B(_0062_),
    .S(_0150_),
    .Z(_0736_));
 MUX2_X1 _1670_ (.A(_0716_),
    .B(_0736_),
    .S(_0202_),
    .Z(_0737_));
 MUX2_X1 _1671_ (.A(_0655_),
    .B(_0737_),
    .S(_0374_),
    .Z(_0738_));
 MUX2_X1 _1672_ (.A(_0546_),
    .B(_0738_),
    .S(_0294_),
    .Z(_0740_));
 OAI21_X1 _1673_ (.A(_0735_),
    .B1(_0740_),
    .B2(_0511_),
    .ZN(_0741_));
 NAND2_X1 _1674_ (.A1(_0124_),
    .A2(_0418_),
    .ZN(_0742_));
 OAI21_X2 _1675_ (.A(_0742_),
    .B1(_0425_),
    .B2(_0124_),
    .ZN(_0743_));
 OAI21_X1 _1676_ (.A(_0336_),
    .B1(_0743_),
    .B2(_0630_),
    .ZN(_0744_));
 INV_X1 _1677_ (.A(_0744_),
    .ZN(_0745_));
 AOI21_X1 _1678_ (.A(_0336_),
    .B1(_0085_),
    .B2(_0563_),
    .ZN(_0746_));
 AOI22_X2 _1679_ (.A1(_0637_),
    .A2(_0395_),
    .B1(_0554_),
    .B2(_0219_),
    .ZN(_0747_));
 NOR2_X1 _1680_ (.A1(_0582_),
    .A2(_0747_),
    .ZN(_0748_));
 MUX2_X1 _1681_ (.A(_0048_),
    .B(_0062_),
    .S(_0099_),
    .Z(_0749_));
 MUX2_X1 _1682_ (.A(_0727_),
    .B(_0749_),
    .S(_0709_),
    .Z(_0751_));
 MUX2_X1 _1683_ (.A(_0660_),
    .B(_0751_),
    .S(_0217_),
    .Z(_0752_));
 MUX2_X1 _1684_ (.A(_0552_),
    .B(_0752_),
    .S(_0219_),
    .Z(_0753_));
 AOI21_X2 _1685_ (.A(_0748_),
    .B1(_0753_),
    .B2(_0255_),
    .ZN(_0754_));
 AOI22_X2 _1686_ (.A1(_0741_),
    .A2(_0745_),
    .B1(_0746_),
    .B2(_0754_),
    .ZN(net25));
 OAI21_X1 _1687_ (.A(_0195_),
    .B1(_0035_),
    .B2(_0277_),
    .ZN(_0755_));
 MUX2_X1 _1688_ (.A(_0053_),
    .B(_0052_),
    .S(net54),
    .Z(_0756_));
 MUX2_X1 _1689_ (.A(_0749_),
    .B(_0756_),
    .S(_0152_),
    .Z(_0757_));
 MUX2_X1 _1690_ (.A(_0674_),
    .B(_0757_),
    .S(_0075_),
    .Z(_0758_));
 MUX2_X1 _1691_ (.A(_0576_),
    .B(_0758_),
    .S(_0256_),
    .Z(_0759_));
 AOI221_X2 _1692_ (.A(_0755_),
    .B1(_0270_),
    .B2(_0038_),
    .C1(_0759_),
    .C2(_0089_),
    .ZN(_0760_));
 AOI21_X1 _1693_ (.A(_0196_),
    .B1(_0250_),
    .B2(_0721_),
    .ZN(_0761_));
 NAND2_X1 _1694_ (.A1(_0473_),
    .A2(_0215_),
    .ZN(_0762_));
 MUX2_X1 _1695_ (.A(_0053_),
    .B(_0052_),
    .S(_0172_),
    .Z(_0763_));
 MUX2_X1 _1696_ (.A(_0736_),
    .B(_0763_),
    .S(_0103_),
    .Z(_0764_));
 MUX2_X1 _1697_ (.A(_0687_),
    .B(_0764_),
    .S(_0374_),
    .Z(_0765_));
 MUX2_X1 _1698_ (.A(_0571_),
    .B(_0765_),
    .S(_0294_),
    .Z(_0766_));
 OAI21_X2 _1699_ (.A(_0762_),
    .B1(_0766_),
    .B2(_0511_),
    .ZN(_0767_));
 AOI21_X2 _1700_ (.A(_0760_),
    .B1(_0761_),
    .B2(_0767_),
    .ZN(net26));
 NAND2_X1 _1701_ (.A1(_0473_),
    .A2(_0304_),
    .ZN(_0768_));
 MUX2_X1 _1702_ (.A(_0049_),
    .B(_0048_),
    .S(_0172_),
    .Z(_0770_));
 MUX2_X1 _1703_ (.A(_0763_),
    .B(_0770_),
    .S(_0183_),
    .Z(_0771_));
 MUX2_X1 _1704_ (.A(_0696_),
    .B(_0771_),
    .S(_0374_),
    .Z(_0772_));
 MUX2_X1 _1705_ (.A(_0597_),
    .B(_0772_),
    .S(_0199_),
    .Z(_0773_));
 OAI21_X2 _1706_ (.A(_0768_),
    .B1(_0773_),
    .B2(_0473_),
    .ZN(_0774_));
 AOI21_X2 _1707_ (.A(_0196_),
    .B1(_0316_),
    .B2(_0721_),
    .ZN(_0775_));
 AOI221_X2 _1708_ (.A(_0335_),
    .B1(_0085_),
    .B2(_0332_),
    .C1(_0346_),
    .C2(_0038_),
    .ZN(_0776_));
 MUX2_X1 _1709_ (.A(_0049_),
    .B(_0048_),
    .S(net54),
    .Z(_0777_));
 MUX2_X1 _1710_ (.A(_0756_),
    .B(_0777_),
    .S(_0202_),
    .Z(_0778_));
 MUX2_X1 _1711_ (.A(_0588_),
    .B(_0778_),
    .S(_0105_),
    .Z(_0779_));
 MUX2_X1 _1712_ (.A(_0703_),
    .B(_0779_),
    .S(_0218_),
    .Z(_0781_));
 NAND2_X2 _1713_ (.A1(_0255_),
    .A2(_0781_),
    .ZN(_0782_));
 AOI22_X4 _1714_ (.A1(_0774_),
    .A2(_0775_),
    .B1(_0776_),
    .B2(_0782_),
    .ZN(net27));
 NOR2_X2 _1715_ (.A1(_0213_),
    .A2(_0035_),
    .ZN(_0783_));
 AOI221_X2 _1716_ (.A(_0335_),
    .B1(_0391_),
    .B2(_0038_),
    .C1(_0783_),
    .C2(_0158_),
    .ZN(_0784_));
 MUX2_X1 _1717_ (.A(_0039_),
    .B(_0053_),
    .S(_0099_),
    .Z(_0785_));
 MUX2_X1 _1718_ (.A(_0777_),
    .B(_0785_),
    .S(net44),
    .Z(_0786_));
 MUX2_X1 _1719_ (.A(_0628_),
    .B(_0786_),
    .S(_0256_),
    .Z(_0787_));
 MUX2_X1 _1720_ (.A(_0730_),
    .B(_0787_),
    .S(_0218_),
    .Z(_0788_));
 NAND2_X1 _1721_ (.A1(_0255_),
    .A2(_0788_),
    .ZN(_0789_));
 MUX2_X1 _1722_ (.A(_0039_),
    .B(_0053_),
    .S(_0148_),
    .Z(_0791_));
 MUX2_X1 _1723_ (.A(_0770_),
    .B(_0791_),
    .S(_0709_),
    .Z(_0792_));
 MUX2_X1 _1724_ (.A(_0717_),
    .B(_0792_),
    .S(_0179_),
    .Z(_0793_));
 MUX2_X1 _1725_ (.A(_0647_),
    .B(_0793_),
    .S(_0170_),
    .Z(_0794_));
 MUX2_X1 _1726_ (.A(_0370_),
    .B(_0794_),
    .S(_0371_),
    .Z(_0795_));
 INV_X1 _1727_ (.A(_0795_),
    .ZN(_0796_));
 NOR2_X2 _1728_ (.A1(_0141_),
    .A2(_0145_),
    .ZN(_0797_));
 AOI21_X2 _1729_ (.A(_0196_),
    .B1(_0797_),
    .B2(_0047_),
    .ZN(_0798_));
 AOI22_X4 _1730_ (.A1(_0784_),
    .A2(_0789_),
    .B1(_0796_),
    .B2(_0798_),
    .ZN(net28));
 MUX2_X1 _1731_ (.A(_0043_),
    .B(_0049_),
    .S(_0148_),
    .Z(_0799_));
 MUX2_X1 _1732_ (.A(_0791_),
    .B(_0799_),
    .S(_0152_),
    .Z(_0801_));
 MUX2_X1 _1733_ (.A(_0737_),
    .B(_0801_),
    .S(_0207_),
    .Z(_0802_));
 MUX2_X1 _1734_ (.A(_0656_),
    .B(_0802_),
    .S(_0198_),
    .Z(_0803_));
 MUX2_X1 _1735_ (.A(_0436_),
    .B(_0803_),
    .S(_0371_),
    .Z(_0804_));
 NOR3_X1 _1736_ (.A1(_0125_),
    .A2(_0418_),
    .A3(_0630_),
    .ZN(_0805_));
 NOR3_X2 _1737_ (.A1(_0196_),
    .A2(_0804_),
    .A3(_0805_),
    .ZN(_0806_));
 MUX2_X1 _1738_ (.A(_0043_),
    .B(_0049_),
    .S(_0099_),
    .Z(_0807_));
 MUX2_X1 _1739_ (.A(_0785_),
    .B(_0807_),
    .S(net44),
    .Z(_0808_));
 MUX2_X1 _1740_ (.A(_0751_),
    .B(_0808_),
    .S(_0217_),
    .Z(_0809_));
 MUX2_X1 _1741_ (.A(_0662_),
    .B(_0809_),
    .S(_0219_),
    .Z(_0810_));
 AOI22_X4 _1742_ (.A1(_0038_),
    .A2(net57),
    .B1(_0810_),
    .B2(_0255_),
    .ZN(_0812_));
 AOI21_X2 _1743_ (.A(_0336_),
    .B1(_0783_),
    .B2(_0562_),
    .ZN(_0813_));
 AOI21_X4 _1744_ (.A(_0806_),
    .B1(_0812_),
    .B2(_0813_),
    .ZN(net29));
 NAND2_X1 _1745_ (.A1(_0374_),
    .A2(_0085_),
    .ZN(_0814_));
 OAI21_X1 _1746_ (.A(_0780_),
    .B1(_0211_),
    .B2(_0814_),
    .ZN(_0815_));
 MUX2_X1 _1747_ (.A(_0098_),
    .B(_0114_),
    .S(net3),
    .Z(_0816_));
 MUX2_X1 _1748_ (.A(_0604_),
    .B(_0816_),
    .S(_0274_),
    .Z(_0817_));
 MUX2_X1 _1749_ (.A(_0241_),
    .B(_0817_),
    .S(_0079_),
    .Z(_0818_));
 MUX2_X1 _1750_ (.A(_0115_),
    .B(_0090_),
    .S(_0045_),
    .Z(_0819_));
 MUX2_X1 _1751_ (.A(_0608_),
    .B(_0819_),
    .S(_0274_),
    .Z(_0820_));
 MUX2_X1 _1752_ (.A(_0230_),
    .B(_0820_),
    .S(_0079_),
    .Z(_0822_));
 MUX2_X1 _1753_ (.A(_0818_),
    .B(_0822_),
    .S(_0352_),
    .Z(_0823_));
 AOI221_X2 _1754_ (.A(_0815_),
    .B1(_0823_),
    .B2(_0088_),
    .C1(_0038_),
    .C2(_0568_),
    .ZN(_0824_));
 NAND2_X1 _1755_ (.A1(_0475_),
    .A2(_0293_),
    .ZN(_0825_));
 MUX2_X1 _1756_ (.A(_0115_),
    .B(_0090_),
    .S(_0172_),
    .Z(_0826_));
 MUX2_X1 _1757_ (.A(_0613_),
    .B(_0826_),
    .S(_0132_),
    .Z(_0827_));
 MUX2_X1 _1758_ (.A(_0098_),
    .B(_0114_),
    .S(_0739_),
    .Z(_0828_));
 MUX2_X1 _1759_ (.A(_0616_),
    .B(_0828_),
    .S(_0133_),
    .Z(_0829_));
 MUX2_X1 _1760_ (.A(_0827_),
    .B(_0829_),
    .S(_0374_),
    .Z(_0830_));
 NAND2_X1 _1761_ (.A1(_0294_),
    .A2(_0830_),
    .ZN(_0831_));
 AOI21_X1 _1762_ (.A(_0197_),
    .B1(_0825_),
    .B2(_0831_),
    .ZN(_0833_));
 AOI21_X1 _1763_ (.A(_0833_),
    .B1(_0585_),
    .B2(_0511_),
    .ZN(_0834_));
 AOI21_X1 _1764_ (.A(_0336_),
    .B1(_0797_),
    .B2(_0581_),
    .ZN(_0835_));
 AOI21_X2 _1765_ (.A(_0824_),
    .B1(_0834_),
    .B2(_0835_),
    .ZN(net30));
 NAND3_X1 _1766_ (.A1(_0197_),
    .A2(_0478_),
    .A3(_0482_),
    .ZN(_0836_));
 NAND2_X1 _1767_ (.A1(_0475_),
    .A2(_0689_),
    .ZN(_0837_));
 MUX2_X1 _1768_ (.A(_0040_),
    .B(_0039_),
    .S(_0172_),
    .Z(_0838_));
 MUX2_X1 _1769_ (.A(_0799_),
    .B(_0838_),
    .S(net42),
    .Z(_0839_));
 MUX2_X1 _1770_ (.A(_0764_),
    .B(_0839_),
    .S(_0168_),
    .Z(_0840_));
 NAND2_X1 _1771_ (.A1(_0190_),
    .A2(_0840_),
    .ZN(_0841_));
 NAND3_X1 _1772_ (.A1(_0894_),
    .A2(_0837_),
    .A3(_0841_),
    .ZN(_0843_));
 AOI221_X2 _1773_ (.A(_0306_),
    .B1(_0146_),
    .B2(_0245_),
    .C1(_0836_),
    .C2(_0843_),
    .ZN(_0844_));
 MUX2_X1 _1774_ (.A(_0040_),
    .B(_0039_),
    .S(_0099_),
    .Z(_0845_));
 MUX2_X1 _1775_ (.A(_0807_),
    .B(_0845_),
    .S(_0709_),
    .Z(_0846_));
 MUX2_X1 _1776_ (.A(_0757_),
    .B(_0846_),
    .S(_0218_),
    .Z(_0847_));
 MUX2_X1 _1777_ (.A(_0676_),
    .B(_0847_),
    .S(_0219_),
    .Z(_0848_));
 NOR2_X1 _1778_ (.A1(_0446_),
    .A2(_0450_),
    .ZN(_0849_));
 NOR2_X1 _1779_ (.A1(_0582_),
    .A2(_0849_),
    .ZN(_0850_));
 AOI21_X1 _1780_ (.A(_0445_),
    .B1(_0454_),
    .B2(_0227_),
    .ZN(_0851_));
 AOI22_X4 _1781_ (.A1(_0848_),
    .A2(_0255_),
    .B1(_0850_),
    .B2(_0851_),
    .ZN(_0852_));
 AOI21_X1 _1782_ (.A(_0336_),
    .B1(_0603_),
    .B2(_0245_),
    .ZN(_0854_));
 AOI21_X4 _1783_ (.A(_0844_),
    .B1(_0852_),
    .B2(_0854_),
    .ZN(net31));
 MUX2_X1 _1784_ (.A(_0044_),
    .B(_0043_),
    .S(_0739_),
    .Z(_0855_));
 MUX2_X1 _1785_ (.A(_0838_),
    .B(_0855_),
    .S(_0183_),
    .Z(_0856_));
 MUX2_X1 _1786_ (.A(_0771_),
    .B(_0856_),
    .S(_0188_),
    .Z(_0857_));
 MUX2_X1 _1787_ (.A(_0697_),
    .B(_0857_),
    .S(_0170_),
    .Z(_0858_));
 MUX2_X1 _1788_ (.A(_0494_),
    .B(_0858_),
    .S(_0371_),
    .Z(_0859_));
 INV_X1 _1789_ (.A(_0859_),
    .ZN(_0860_));
 AOI21_X2 _1790_ (.A(_0196_),
    .B1(_0146_),
    .B2(_0502_),
    .ZN(_0861_));
 OR4_X2 _1791_ (.A1(_0582_),
    .A2(_0496_),
    .A3(_0499_),
    .A4(_0500_),
    .ZN(_0862_));
 MUX2_X1 _1792_ (.A(_0044_),
    .B(_0043_),
    .S(_0099_),
    .Z(_0864_));
 MUX2_X1 _1793_ (.A(_0845_),
    .B(_0864_),
    .S(_0152_),
    .Z(_0865_));
 MUX2_X1 _1794_ (.A(_0702_),
    .B(_0865_),
    .S(_0105_),
    .Z(_0866_));
 MUX2_X1 _1795_ (.A(_0779_),
    .B(_0866_),
    .S(_0218_),
    .Z(_0867_));
 AOI221_X2 _1796_ (.A(_0335_),
    .B1(_0603_),
    .B2(_0502_),
    .C1(_0089_),
    .C2(_0867_),
    .ZN(_0868_));
 AOI22_X4 _1797_ (.A1(_0860_),
    .A2(_0861_),
    .B1(_0868_),
    .B2(_0862_),
    .ZN(net32));
 MUX2_X1 _1798_ (.A(_0096_),
    .B(_0819_),
    .S(net2),
    .Z(_0869_));
 MUX2_X1 _1799_ (.A(_0119_),
    .B(_0816_),
    .S(_0056_),
    .Z(_0870_));
 MUX2_X1 _1800_ (.A(_0869_),
    .B(_0870_),
    .S(_0059_),
    .Z(_0871_));
 MUX2_X1 _1801_ (.A(_0319_),
    .B(_0871_),
    .S(_0105_),
    .Z(_0872_));
 MUX2_X1 _1802_ (.A(_0600_),
    .B(_0872_),
    .S(_0234_),
    .Z(_0874_));
 AOI221_X2 _1803_ (.A(_0306_),
    .B1(_0303_),
    .B2(_0783_),
    .C1(_0143_),
    .C2(_0874_),
    .ZN(_0875_));
 AOI21_X1 _1804_ (.A(_0129_),
    .B1(_0797_),
    .B2(net66),
    .ZN(_0876_));
 MUX2_X1 _1805_ (.A(_0177_),
    .B(_0826_),
    .S(_0103_),
    .Z(_0877_));
 NOR2_X1 _1806_ (.A1(_0374_),
    .A2(_0877_),
    .ZN(_0878_));
 MUX2_X1 _1807_ (.A(_0182_),
    .B(_0828_),
    .S(_0183_),
    .Z(_0879_));
 NOR2_X1 _1808_ (.A1(_0213_),
    .A2(_0879_),
    .ZN(_0880_));
 NOR3_X2 _1809_ (.A1(_0035_),
    .A2(_0878_),
    .A3(_0880_),
    .ZN(_0881_));
 MUX2_X1 _1810_ (.A(_0328_),
    .B(_0332_),
    .S(_0811_),
    .Z(_0882_));
 AOI221_X2 _1811_ (.A(_0881_),
    .B1(_0882_),
    .B2(_0475_),
    .C1(_0333_),
    .C2(_0325_),
    .ZN(_0883_));
 AOI21_X2 _1812_ (.A(_0875_),
    .B1(_0876_),
    .B2(_0883_),
    .ZN(net33));
 OAI21_X1 _1813_ (.A(_0780_),
    .B1(_0035_),
    .B2(_0641_),
    .ZN(_0885_));
 MUX2_X1 _1814_ (.A(_0074_),
    .B(_0097_),
    .S(_0079_),
    .Z(_0886_));
 MUX2_X1 _1815_ (.A(_0122_),
    .B(_0886_),
    .S(_0352_),
    .Z(_0887_));
 OR2_X1 _1816_ (.A1(_0643_),
    .A2(_0450_),
    .ZN(_0888_));
 NAND3_X1 _1817_ (.A1(_0638_),
    .A2(_0639_),
    .A3(_0888_),
    .ZN(_0889_));
 AOI221_X2 _1818_ (.A(_0885_),
    .B1(_0887_),
    .B2(_0088_),
    .C1(_0038_),
    .C2(_0889_),
    .ZN(_0890_));
 NOR2_X1 _1819_ (.A1(_0632_),
    .A2(_0630_),
    .ZN(_0891_));
 NOR2_X1 _1820_ (.A1(_0129_),
    .A2(_0891_),
    .ZN(_0892_));
 OR3_X1 _1821_ (.A1(_0371_),
    .A2(_0635_),
    .A3(_0636_),
    .ZN(_0893_));
 MUX2_X1 _1822_ (.A(_0178_),
    .B(_0184_),
    .S(_0374_),
    .Z(_0895_));
 MUX2_X1 _1823_ (.A(_0375_),
    .B(_0895_),
    .S(_0294_),
    .Z(_0896_));
 OAI21_X2 _1824_ (.A(_0893_),
    .B1(_0896_),
    .B2(_0511_),
    .ZN(_0897_));
 AOI21_X4 _1825_ (.A(_0890_),
    .B1(_0892_),
    .B2(_0897_),
    .ZN(net34));
 AOI21_X1 _1826_ (.A(_0306_),
    .B1(_0085_),
    .B2(_0431_),
    .ZN(_0898_));
 OAI21_X1 _1827_ (.A(_0898_),
    .B1(_0652_),
    .B2(_0582_),
    .ZN(_0899_));
 MUX2_X1 _1828_ (.A(_0421_),
    .B(_0606_),
    .S(_0079_),
    .Z(_0900_));
 MUX2_X1 _1829_ (.A(_0610_),
    .B(_0900_),
    .S(_0125_),
    .Z(_0901_));
 AOI21_X2 _1830_ (.A(_0899_),
    .B1(_0901_),
    .B2(_0255_),
    .ZN(_0902_));
 AOI21_X2 _1831_ (.A(_0129_),
    .B1(_0397_),
    .B2(_0721_),
    .ZN(_0903_));
 MUX2_X1 _1832_ (.A(_0620_),
    .B(_0614_),
    .S(_0188_),
    .Z(_0905_));
 MUX2_X1 _1833_ (.A(_0410_),
    .B(_0905_),
    .S(_0170_),
    .Z(_0906_));
 MUX2_X1 _1834_ (.A(_0665_),
    .B(_0906_),
    .S(_0192_),
    .Z(_0907_));
 INV_X1 _1835_ (.A(_0907_),
    .ZN(_0908_));
 AOI21_X4 _1836_ (.A(_0902_),
    .B1(_0903_),
    .B2(_0908_),
    .ZN(net35));
 OAI21_X1 _1837_ (.A(_0195_),
    .B1(_0454_),
    .B2(_0630_),
    .ZN(_0909_));
 NAND2_X1 _1838_ (.A1(_0475_),
    .A2(_0460_),
    .ZN(_0910_));
 MUX2_X1 _1839_ (.A(_0292_),
    .B(_0827_),
    .S(_0188_),
    .Z(_0911_));
 NAND2_X1 _1840_ (.A1(_0199_),
    .A2(_0911_),
    .ZN(_0912_));
 NAND3_X1 _1841_ (.A1(_0371_),
    .A2(_0910_),
    .A3(_0912_),
    .ZN(_0913_));
 NAND2_X1 _1842_ (.A1(_0197_),
    .A2(_0684_),
    .ZN(_0915_));
 AOI21_X2 _1843_ (.A(_0909_),
    .B1(_0913_),
    .B2(_0915_),
    .ZN(_0916_));
 NAND3_X1 _1844_ (.A1(_0085_),
    .A2(_0476_),
    .A3(_0477_),
    .ZN(_0917_));
 AND2_X1 _1845_ (.A1(_0335_),
    .A2(_0917_),
    .ZN(_0918_));
 NOR2_X1 _1846_ (.A1(_0234_),
    .A2(_0669_),
    .ZN(_0919_));
 MUX2_X1 _1847_ (.A(_0242_),
    .B(_0822_),
    .S(_0217_),
    .Z(_0920_));
 AOI21_X2 _1848_ (.A(_0919_),
    .B1(_0920_),
    .B2(_0234_),
    .ZN(_0921_));
 NOR2_X1 _1849_ (.A1(_0196_),
    .A2(_0143_),
    .ZN(_0922_));
 AOI221_X2 _1850_ (.A(_0916_),
    .B1(_0918_),
    .B2(_0921_),
    .C1(_0922_),
    .C2(_0917_),
    .ZN(net36));
 NAND2_X1 _1851_ (.A1(_0197_),
    .A2(_0693_),
    .ZN(_0923_));
 MUX2_X1 _1852_ (.A(_0327_),
    .B(_0877_),
    .S(_0179_),
    .Z(_0001_));
 NOR2_X1 _1853_ (.A1(_0035_),
    .A2(_0001_),
    .ZN(_0002_));
 NOR3_X1 _1854_ (.A1(_0811_),
    .A2(_0170_),
    .A3(_0507_),
    .ZN(_0003_));
 NOR2_X2 _1855_ (.A1(_0002_),
    .A2(_0003_),
    .ZN(_0004_));
 AOI221_X2 _1856_ (.A(_0335_),
    .B1(_0495_),
    .B2(_0721_),
    .C1(_0923_),
    .C2(_0004_),
    .ZN(_0005_));
 MUX2_X1 _1857_ (.A(_0318_),
    .B(_0869_),
    .S(_0075_),
    .Z(_0006_));
 MUX2_X1 _1858_ (.A(_0487_),
    .B(_0006_),
    .S(_0256_),
    .Z(_0007_));
 MUX2_X1 _1859_ (.A(_0711_),
    .B(_0007_),
    .S(_0234_),
    .Z(_0008_));
 AOI22_X2 _1860_ (.A1(_0085_),
    .A2(_0490_),
    .B1(_0008_),
    .B2(_0143_),
    .ZN(_0009_));
 AOI21_X2 _1861_ (.A(_0005_),
    .B1(_0009_),
    .B2(_0129_),
    .ZN(net37));
 NAND3_X1 _1862_ (.A1(_0219_),
    .A2(_0060_),
    .A3(_0038_),
    .ZN(_0011_));
 AND2_X1 _1863_ (.A1(_0128_),
    .A2(_0011_),
    .ZN(_0012_));
 MUX2_X1 _1864_ (.A(_0067_),
    .B(_0113_),
    .S(_0080_),
    .Z(_0013_));
 OAI221_X1 _1865_ (.A(_0255_),
    .B1(_0218_),
    .B2(_0013_),
    .C1(_0097_),
    .C2(_0141_),
    .ZN(_0014_));
 NOR2_X1 _1866_ (.A1(_0074_),
    .A2(_0267_),
    .ZN(_0015_));
 OAI221_X1 _1867_ (.A(_0012_),
    .B1(_0014_),
    .B2(_0015_),
    .C1(_0473_),
    .C2(_0714_),
    .ZN(_0016_));
 NAND2_X1 _1868_ (.A1(_0159_),
    .A2(_0333_),
    .ZN(_0017_));
 AOI221_X2 _1869_ (.A(_0769_),
    .B1(_0088_),
    .B2(_0723_),
    .C1(_0724_),
    .C2(_0721_),
    .ZN(_0018_));
 MUX2_X1 _1870_ (.A(_0169_),
    .B(_0180_),
    .S(_0199_),
    .Z(_0019_));
 INV_X1 _1871_ (.A(_0019_),
    .ZN(_0020_));
 OAI211_X2 _1872_ (.A(_0017_),
    .B(_0018_),
    .C1(_0020_),
    .C2(_0473_),
    .ZN(_0022_));
 AND2_X2 _1873_ (.A1(_0016_),
    .A2(_0022_),
    .ZN(net38));
 MUX2_X1 _1874_ (.A(_0416_),
    .B(_0424_),
    .S(_0225_),
    .Z(_0023_));
 NAND3_X1 _1875_ (.A1(_0088_),
    .A2(_0125_),
    .A3(_0023_),
    .ZN(_0024_));
 OAI21_X1 _1876_ (.A(_0024_),
    .B1(_0633_),
    .B2(_0743_),
    .ZN(_0025_));
 AND3_X2 _1877_ (.A1(_0088_),
    .A2(_0218_),
    .A3(_0900_),
    .ZN(_0026_));
 NAND2_X1 _1878_ (.A1(_0335_),
    .A2(_0734_),
    .ZN(_0027_));
 OR3_X1 _1879_ (.A1(_0025_),
    .A2(_0026_),
    .A3(_0027_),
    .ZN(_0028_));
 AOI21_X1 _1880_ (.A(_0128_),
    .B1(_0333_),
    .B2(_0563_),
    .ZN(_0029_));
 MUX2_X1 _1881_ (.A(_0560_),
    .B(_0621_),
    .S(_0170_),
    .Z(_0030_));
 INV_X1 _1882_ (.A(_0030_),
    .ZN(_0032_));
 OAI221_X1 _1883_ (.A(_0029_),
    .B1(_0032_),
    .B2(_0473_),
    .C1(_0145_),
    .C2(_0747_),
    .ZN(_0033_));
 OR4_X2 _1884_ (.A1(_0192_),
    .A2(_0306_),
    .A3(_0025_),
    .A4(_0026_),
    .ZN(_0034_));
 AND3_X4 _1885_ (.A1(_0034_),
    .A2(_0033_),
    .A3(_0028_),
    .ZN(net39));
 HA_X1 _1886_ (.A(_0709_),
    .B(_0925_),
    .CO(_0926_),
    .S(_0927_));
 BUF_X2 clone1 (.A(_0927_),
    .Z(net1));
 INV_X2 clone2 (.A(_0677_),
    .ZN(net2));
 BUF_X4 clone4 (.A(_0688_),
    .Z(net4));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_239 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_240 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_241 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_242 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_243 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_244 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_245 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_246 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_247 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_248 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_249 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_250 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_251 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_252 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_253 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_254 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_255 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_256 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_257 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_258 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_259 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_260 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_261 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_262 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_263 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_264 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_267 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_268 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_269 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_270 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_271 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_272 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_273 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_274 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_275 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_276 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_277 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_278 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_279 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_280 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_281 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_282 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_283 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_284 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_285 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_286 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_287 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_288 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_289 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_290 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_291 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_292 ();
 CLKBUF_X3 input1 (.A(data_in[1]),
    .Z(net5));
 CLKBUF_X2 input2 (.A(rotate),
    .Z(net6));
 BUF_X2 input3 (.A(shift_amount[2]),
    .Z(net7));
 BUF_X1 output4 (.A(net8),
    .Z(data_out[0]));
 BUF_X1 output5 (.A(net9),
    .Z(data_out[10]));
 BUF_X1 output6 (.A(net10),
    .Z(data_out[11]));
 BUF_X1 output7 (.A(net11),
    .Z(data_out[12]));
 BUF_X2 output8 (.A(net12),
    .Z(data_out[13]));
 BUF_X1 output9 (.A(net13),
    .Z(data_out[14]));
 BUF_X1 output10 (.A(net14),
    .Z(data_out[15]));
 BUF_X1 output11 (.A(net15),
    .Z(data_out[16]));
 BUF_X1 output12 (.A(net16),
    .Z(data_out[17]));
 BUF_X1 output13 (.A(net17),
    .Z(data_out[18]));
 BUF_X1 output14 (.A(net18),
    .Z(data_out[19]));
 BUF_X1 output15 (.A(net19),
    .Z(data_out[1]));
 BUF_X1 output16 (.A(net20),
    .Z(data_out[20]));
 BUF_X1 output17 (.A(net21),
    .Z(data_out[21]));
 BUF_X1 output18 (.A(net22),
    .Z(data_out[22]));
 BUF_X2 output19 (.A(net23),
    .Z(data_out[23]));
 BUF_X1 output20 (.A(net24),
    .Z(data_out[24]));
 BUF_X1 output21 (.A(net25),
    .Z(data_out[25]));
 BUF_X1 output22 (.A(net26),
    .Z(data_out[26]));
 BUF_X1 output23 (.A(net27),
    .Z(data_out[27]));
 BUF_X1 output24 (.A(net28),
    .Z(data_out[28]));
 BUF_X1 output25 (.A(net29),
    .Z(data_out[29]));
 BUF_X1 output26 (.A(net30),
    .Z(data_out[2]));
 BUF_X1 output27 (.A(net31),
    .Z(data_out[30]));
 BUF_X2 output28 (.A(net32),
    .Z(data_out[31]));
 BUF_X1 output29 (.A(net33),
    .Z(data_out[3]));
 BUF_X1 output30 (.A(net34),
    .Z(data_out[4]));
 BUF_X1 output31 (.A(net35),
    .Z(data_out[5]));
 BUF_X1 output32 (.A(net36),
    .Z(data_out[6]));
 BUF_X1 output33 (.A(net37),
    .Z(data_out[7]));
 BUF_X1 output34 (.A(net38),
    .Z(data_out[8]));
 BUF_X1 output35 (.A(net39),
    .Z(data_out[9]));
 BUF_X1 rebuffer1 (.A(_0060_),
    .Z(net40));
 BUF_X1 rebuffer2 (.A(_0046_),
    .Z(net41));
 BUF_X16 clone5 (.A(_0698_),
    .Z(net42));
 BUF_X2 rebuffer11 (.A(_0600_),
    .Z(net48));
 BUF_X1 rebuffer14 (.A(_0711_),
    .Z(net51));
 BUF_X8 rebuffer17 (.A(_0045_),
    .Z(net54));
 BUF_X2 rebuffer20 (.A(_0402_),
    .Z(net57));
 BUF_X1 rebuffer28 (.A(_0338_),
    .Z(net65));
 BUF_X1 rebuffer29 (.A(net65),
    .Z(net66));
 BUF_X4 rebuffer68 (.A(_0058_),
    .Z(net105));
 BUF_X4 clone27 (.A(net69),
    .Z(net68));
 BUF_X4 clone28 (.A(net70),
    .Z(net69));
 BUF_X1 rebuffer30 (.A(_0927_),
    .Z(net70));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X8 FILLER_0_257 ();
 FILLCELL_X4 FILLER_0_265 ();
 FILLCELL_X4 FILLER_0_277 ();
 FILLCELL_X1 FILLER_0_281 ();
 FILLCELL_X1 FILLER_0_302 ();
 FILLCELL_X1 FILLER_0_319 ();
 FILLCELL_X4 FILLER_0_328 ();
 FILLCELL_X2 FILLER_0_336 ();
 FILLCELL_X1 FILLER_0_342 ();
 FILLCELL_X4 FILLER_0_355 ();
 FILLCELL_X32 FILLER_0_364 ();
 FILLCELL_X32 FILLER_0_396 ();
 FILLCELL_X32 FILLER_0_428 ();
 FILLCELL_X32 FILLER_0_460 ();
 FILLCELL_X32 FILLER_0_492 ();
 FILLCELL_X32 FILLER_0_524 ();
 FILLCELL_X32 FILLER_0_556 ();
 FILLCELL_X32 FILLER_0_588 ();
 FILLCELL_X8 FILLER_0_620 ();
 FILLCELL_X2 FILLER_0_628 ();
 FILLCELL_X1 FILLER_0_630 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X32 FILLER_0_792 ();
 FILLCELL_X32 FILLER_0_824 ();
 FILLCELL_X4 FILLER_0_856 ();
 FILLCELL_X2 FILLER_0_860 ();
 FILLCELL_X1 FILLER_0_862 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X16 FILLER_1_289 ();
 FILLCELL_X8 FILLER_1_305 ();
 FILLCELL_X4 FILLER_1_313 ();
 FILLCELL_X1 FILLER_1_317 ();
 FILLCELL_X16 FILLER_1_322 ();
 FILLCELL_X1 FILLER_1_338 ();
 FILLCELL_X32 FILLER_1_348 ();
 FILLCELL_X32 FILLER_1_380 ();
 FILLCELL_X32 FILLER_1_412 ();
 FILLCELL_X32 FILLER_1_444 ();
 FILLCELL_X32 FILLER_1_476 ();
 FILLCELL_X32 FILLER_1_508 ();
 FILLCELL_X32 FILLER_1_540 ();
 FILLCELL_X32 FILLER_1_572 ();
 FILLCELL_X32 FILLER_1_604 ();
 FILLCELL_X32 FILLER_1_636 ();
 FILLCELL_X32 FILLER_1_668 ();
 FILLCELL_X32 FILLER_1_700 ();
 FILLCELL_X32 FILLER_1_732 ();
 FILLCELL_X32 FILLER_1_764 ();
 FILLCELL_X32 FILLER_1_796 ();
 FILLCELL_X32 FILLER_1_828 ();
 FILLCELL_X2 FILLER_1_860 ();
 FILLCELL_X1 FILLER_1_862 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X8 FILLER_2_289 ();
 FILLCELL_X2 FILLER_2_297 ();
 FILLCELL_X1 FILLER_2_299 ();
 FILLCELL_X16 FILLER_2_304 ();
 FILLCELL_X8 FILLER_2_324 ();
 FILLCELL_X4 FILLER_2_332 ();
 FILLCELL_X2 FILLER_2_336 ();
 FILLCELL_X1 FILLER_2_338 ();
 FILLCELL_X32 FILLER_2_343 ();
 FILLCELL_X32 FILLER_2_375 ();
 FILLCELL_X32 FILLER_2_407 ();
 FILLCELL_X32 FILLER_2_439 ();
 FILLCELL_X32 FILLER_2_471 ();
 FILLCELL_X32 FILLER_2_503 ();
 FILLCELL_X32 FILLER_2_535 ();
 FILLCELL_X32 FILLER_2_567 ();
 FILLCELL_X32 FILLER_2_599 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X32 FILLER_2_824 ();
 FILLCELL_X4 FILLER_2_856 ();
 FILLCELL_X2 FILLER_2_860 ();
 FILLCELL_X1 FILLER_2_862 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X8 FILLER_3_321 ();
 FILLCELL_X2 FILLER_3_333 ();
 FILLCELL_X1 FILLER_3_335 ();
 FILLCELL_X32 FILLER_3_340 ();
 FILLCELL_X32 FILLER_3_372 ();
 FILLCELL_X32 FILLER_3_404 ();
 FILLCELL_X32 FILLER_3_436 ();
 FILLCELL_X32 FILLER_3_468 ();
 FILLCELL_X32 FILLER_3_500 ();
 FILLCELL_X32 FILLER_3_532 ();
 FILLCELL_X32 FILLER_3_564 ();
 FILLCELL_X32 FILLER_3_596 ();
 FILLCELL_X32 FILLER_3_628 ();
 FILLCELL_X32 FILLER_3_660 ();
 FILLCELL_X32 FILLER_3_692 ();
 FILLCELL_X32 FILLER_3_724 ();
 FILLCELL_X32 FILLER_3_756 ();
 FILLCELL_X32 FILLER_3_788 ();
 FILLCELL_X32 FILLER_3_820 ();
 FILLCELL_X8 FILLER_3_852 ();
 FILLCELL_X2 FILLER_3_860 ();
 FILLCELL_X1 FILLER_3_862 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X4 FILLER_4_856 ();
 FILLCELL_X2 FILLER_4_860 ();
 FILLCELL_X1 FILLER_4_862 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X32 FILLER_5_801 ();
 FILLCELL_X16 FILLER_5_833 ();
 FILLCELL_X8 FILLER_5_849 ();
 FILLCELL_X4 FILLER_5_857 ();
 FILLCELL_X2 FILLER_5_861 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X32 FILLER_6_824 ();
 FILLCELL_X4 FILLER_6_856 ();
 FILLCELL_X2 FILLER_6_860 ();
 FILLCELL_X1 FILLER_6_862 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X8 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_301 ();
 FILLCELL_X32 FILLER_7_333 ();
 FILLCELL_X32 FILLER_7_365 ();
 FILLCELL_X32 FILLER_7_397 ();
 FILLCELL_X32 FILLER_7_429 ();
 FILLCELL_X32 FILLER_7_461 ();
 FILLCELL_X32 FILLER_7_493 ();
 FILLCELL_X32 FILLER_7_525 ();
 FILLCELL_X32 FILLER_7_557 ();
 FILLCELL_X32 FILLER_7_589 ();
 FILLCELL_X32 FILLER_7_621 ();
 FILLCELL_X32 FILLER_7_653 ();
 FILLCELL_X32 FILLER_7_685 ();
 FILLCELL_X32 FILLER_7_717 ();
 FILLCELL_X32 FILLER_7_749 ();
 FILLCELL_X32 FILLER_7_781 ();
 FILLCELL_X32 FILLER_7_813 ();
 FILLCELL_X16 FILLER_7_845 ();
 FILLCELL_X2 FILLER_7_861 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X32 FILLER_8_824 ();
 FILLCELL_X4 FILLER_8_856 ();
 FILLCELL_X2 FILLER_8_860 ();
 FILLCELL_X1 FILLER_8_862 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X32 FILLER_9_801 ();
 FILLCELL_X16 FILLER_9_833 ();
 FILLCELL_X8 FILLER_9_849 ();
 FILLCELL_X4 FILLER_9_857 ();
 FILLCELL_X2 FILLER_9_861 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X32 FILLER_10_824 ();
 FILLCELL_X4 FILLER_10_856 ();
 FILLCELL_X2 FILLER_10_860 ();
 FILLCELL_X1 FILLER_10_862 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X16 FILLER_11_833 ();
 FILLCELL_X8 FILLER_11_849 ();
 FILLCELL_X4 FILLER_11_857 ();
 FILLCELL_X2 FILLER_11_861 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X4 FILLER_12_856 ();
 FILLCELL_X2 FILLER_12_860 ();
 FILLCELL_X1 FILLER_12_862 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X16 FILLER_13_833 ();
 FILLCELL_X8 FILLER_13_849 ();
 FILLCELL_X4 FILLER_13_857 ();
 FILLCELL_X2 FILLER_13_861 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X16 FILLER_14_385 ();
 FILLCELL_X8 FILLER_14_401 ();
 FILLCELL_X32 FILLER_14_423 ();
 FILLCELL_X32 FILLER_14_455 ();
 FILLCELL_X32 FILLER_14_487 ();
 FILLCELL_X32 FILLER_14_519 ();
 FILLCELL_X32 FILLER_14_551 ();
 FILLCELL_X32 FILLER_14_583 ();
 FILLCELL_X16 FILLER_14_615 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X4 FILLER_14_856 ();
 FILLCELL_X2 FILLER_14_860 ();
 FILLCELL_X1 FILLER_14_862 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X2 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_295 ();
 FILLCELL_X32 FILLER_15_327 ();
 FILLCELL_X8 FILLER_15_359 ();
 FILLCELL_X1 FILLER_15_367 ();
 FILLCELL_X8 FILLER_15_375 ();
 FILLCELL_X2 FILLER_15_383 ();
 FILLCELL_X4 FILLER_15_411 ();
 FILLCELL_X2 FILLER_15_415 ();
 FILLCELL_X1 FILLER_15_417 ();
 FILLCELL_X1 FILLER_15_425 ();
 FILLCELL_X4 FILLER_15_438 ();
 FILLCELL_X1 FILLER_15_442 ();
 FILLCELL_X4 FILLER_15_450 ();
 FILLCELL_X32 FILLER_15_461 ();
 FILLCELL_X32 FILLER_15_493 ();
 FILLCELL_X32 FILLER_15_525 ();
 FILLCELL_X32 FILLER_15_557 ();
 FILLCELL_X32 FILLER_15_589 ();
 FILLCELL_X32 FILLER_15_621 ();
 FILLCELL_X32 FILLER_15_653 ();
 FILLCELL_X32 FILLER_15_685 ();
 FILLCELL_X32 FILLER_15_717 ();
 FILLCELL_X32 FILLER_15_749 ();
 FILLCELL_X32 FILLER_15_781 ();
 FILLCELL_X32 FILLER_15_813 ();
 FILLCELL_X16 FILLER_15_845 ();
 FILLCELL_X2 FILLER_15_861 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X4 FILLER_16_289 ();
 FILLCELL_X2 FILLER_16_293 ();
 FILLCELL_X1 FILLER_16_295 ();
 FILLCELL_X32 FILLER_16_300 ();
 FILLCELL_X4 FILLER_16_346 ();
 FILLCELL_X1 FILLER_16_350 ();
 FILLCELL_X16 FILLER_16_358 ();
 FILLCELL_X4 FILLER_16_374 ();
 FILLCELL_X2 FILLER_16_378 ();
 FILLCELL_X4 FILLER_16_387 ();
 FILLCELL_X2 FILLER_16_391 ();
 FILLCELL_X1 FILLER_16_393 ();
 FILLCELL_X8 FILLER_16_401 ();
 FILLCELL_X2 FILLER_16_409 ();
 FILLCELL_X1 FILLER_16_411 ();
 FILLCELL_X8 FILLER_16_419 ();
 FILLCELL_X1 FILLER_16_427 ();
 FILLCELL_X16 FILLER_16_435 ();
 FILLCELL_X2 FILLER_16_451 ();
 FILLCELL_X32 FILLER_16_474 ();
 FILLCELL_X32 FILLER_16_506 ();
 FILLCELL_X32 FILLER_16_538 ();
 FILLCELL_X32 FILLER_16_570 ();
 FILLCELL_X16 FILLER_16_602 ();
 FILLCELL_X8 FILLER_16_618 ();
 FILLCELL_X4 FILLER_16_626 ();
 FILLCELL_X1 FILLER_16_630 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X4 FILLER_16_856 ();
 FILLCELL_X2 FILLER_16_860 ();
 FILLCELL_X1 FILLER_16_862 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X16 FILLER_17_321 ();
 FILLCELL_X8 FILLER_17_337 ();
 FILLCELL_X1 FILLER_17_359 ();
 FILLCELL_X32 FILLER_17_367 ();
 FILLCELL_X4 FILLER_17_404 ();
 FILLCELL_X1 FILLER_17_408 ();
 FILLCELL_X32 FILLER_17_416 ();
 FILLCELL_X32 FILLER_17_448 ();
 FILLCELL_X16 FILLER_17_480 ();
 FILLCELL_X4 FILLER_17_496 ();
 FILLCELL_X2 FILLER_17_500 ();
 FILLCELL_X32 FILLER_17_516 ();
 FILLCELL_X32 FILLER_17_548 ();
 FILLCELL_X32 FILLER_17_580 ();
 FILLCELL_X32 FILLER_17_612 ();
 FILLCELL_X32 FILLER_17_644 ();
 FILLCELL_X32 FILLER_17_676 ();
 FILLCELL_X32 FILLER_17_708 ();
 FILLCELL_X32 FILLER_17_740 ();
 FILLCELL_X32 FILLER_17_772 ();
 FILLCELL_X32 FILLER_17_804 ();
 FILLCELL_X16 FILLER_17_836 ();
 FILLCELL_X8 FILLER_17_852 ();
 FILLCELL_X2 FILLER_17_860 ();
 FILLCELL_X1 FILLER_17_862 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X16 FILLER_18_257 ();
 FILLCELL_X8 FILLER_18_273 ();
 FILLCELL_X4 FILLER_18_281 ();
 FILLCELL_X2 FILLER_18_285 ();
 FILLCELL_X1 FILLER_18_287 ();
 FILLCELL_X32 FILLER_18_292 ();
 FILLCELL_X4 FILLER_18_324 ();
 FILLCELL_X1 FILLER_18_328 ();
 FILLCELL_X8 FILLER_18_336 ();
 FILLCELL_X2 FILLER_18_351 ();
 FILLCELL_X1 FILLER_18_353 ();
 FILLCELL_X4 FILLER_18_361 ();
 FILLCELL_X1 FILLER_18_365 ();
 FILLCELL_X2 FILLER_18_373 ();
 FILLCELL_X1 FILLER_18_375 ();
 FILLCELL_X16 FILLER_18_383 ();
 FILLCELL_X4 FILLER_18_399 ();
 FILLCELL_X16 FILLER_18_410 ();
 FILLCELL_X8 FILLER_18_426 ();
 FILLCELL_X8 FILLER_18_441 ();
 FILLCELL_X2 FILLER_18_449 ();
 FILLCELL_X4 FILLER_18_458 ();
 FILLCELL_X2 FILLER_18_462 ();
 FILLCELL_X1 FILLER_18_464 ();
 FILLCELL_X8 FILLER_18_472 ();
 FILLCELL_X1 FILLER_18_480 ();
 FILLCELL_X1 FILLER_18_495 ();
 FILLCELL_X16 FILLER_18_503 ();
 FILLCELL_X4 FILLER_18_526 ();
 FILLCELL_X2 FILLER_18_530 ();
 FILLCELL_X1 FILLER_18_532 ();
 FILLCELL_X32 FILLER_18_538 ();
 FILLCELL_X32 FILLER_18_570 ();
 FILLCELL_X16 FILLER_18_602 ();
 FILLCELL_X8 FILLER_18_618 ();
 FILLCELL_X4 FILLER_18_626 ();
 FILLCELL_X1 FILLER_18_630 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X4 FILLER_18_856 ();
 FILLCELL_X2 FILLER_18_860 ();
 FILLCELL_X1 FILLER_18_862 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X4 FILLER_19_321 ();
 FILLCELL_X1 FILLER_19_325 ();
 FILLCELL_X4 FILLER_19_333 ();
 FILLCELL_X4 FILLER_19_344 ();
 FILLCELL_X2 FILLER_19_348 ();
 FILLCELL_X1 FILLER_19_350 ();
 FILLCELL_X16 FILLER_19_358 ();
 FILLCELL_X8 FILLER_19_374 ();
 FILLCELL_X1 FILLER_19_382 ();
 FILLCELL_X8 FILLER_19_390 ();
 FILLCELL_X4 FILLER_19_398 ();
 FILLCELL_X2 FILLER_19_402 ();
 FILLCELL_X2 FILLER_19_418 ();
 FILLCELL_X8 FILLER_19_434 ();
 FILLCELL_X4 FILLER_19_442 ();
 FILLCELL_X1 FILLER_19_446 ();
 FILLCELL_X8 FILLER_19_468 ();
 FILLCELL_X4 FILLER_19_476 ();
 FILLCELL_X2 FILLER_19_480 ();
 FILLCELL_X16 FILLER_19_492 ();
 FILLCELL_X4 FILLER_19_508 ();
 FILLCELL_X4 FILLER_19_526 ();
 FILLCELL_X4 FILLER_19_537 ();
 FILLCELL_X1 FILLER_19_541 ();
 FILLCELL_X32 FILLER_19_549 ();
 FILLCELL_X32 FILLER_19_581 ();
 FILLCELL_X32 FILLER_19_613 ();
 FILLCELL_X32 FILLER_19_645 ();
 FILLCELL_X32 FILLER_19_677 ();
 FILLCELL_X32 FILLER_19_709 ();
 FILLCELL_X32 FILLER_19_741 ();
 FILLCELL_X32 FILLER_19_773 ();
 FILLCELL_X32 FILLER_19_805 ();
 FILLCELL_X16 FILLER_19_837 ();
 FILLCELL_X8 FILLER_19_853 ();
 FILLCELL_X2 FILLER_19_861 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X8 FILLER_20_321 ();
 FILLCELL_X16 FILLER_20_336 ();
 FILLCELL_X8 FILLER_20_352 ();
 FILLCELL_X2 FILLER_20_360 ();
 FILLCELL_X4 FILLER_20_369 ();
 FILLCELL_X2 FILLER_20_373 ();
 FILLCELL_X1 FILLER_20_375 ();
 FILLCELL_X8 FILLER_20_383 ();
 FILLCELL_X4 FILLER_20_391 ();
 FILLCELL_X2 FILLER_20_395 ();
 FILLCELL_X1 FILLER_20_397 ();
 FILLCELL_X4 FILLER_20_405 ();
 FILLCELL_X1 FILLER_20_409 ();
 FILLCELL_X8 FILLER_20_417 ();
 FILLCELL_X4 FILLER_20_425 ();
 FILLCELL_X1 FILLER_20_429 ();
 FILLCELL_X8 FILLER_20_437 ();
 FILLCELL_X2 FILLER_20_445 ();
 FILLCELL_X32 FILLER_20_454 ();
 FILLCELL_X16 FILLER_20_486 ();
 FILLCELL_X2 FILLER_20_502 ();
 FILLCELL_X16 FILLER_20_518 ();
 FILLCELL_X8 FILLER_20_534 ();
 FILLCELL_X2 FILLER_20_542 ();
 FILLCELL_X1 FILLER_20_544 ();
 FILLCELL_X32 FILLER_20_552 ();
 FILLCELL_X32 FILLER_20_584 ();
 FILLCELL_X8 FILLER_20_616 ();
 FILLCELL_X4 FILLER_20_624 ();
 FILLCELL_X2 FILLER_20_628 ();
 FILLCELL_X1 FILLER_20_630 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X4 FILLER_20_856 ();
 FILLCELL_X2 FILLER_20_860 ();
 FILLCELL_X1 FILLER_20_862 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X16 FILLER_21_321 ();
 FILLCELL_X1 FILLER_21_337 ();
 FILLCELL_X1 FILLER_21_352 ();
 FILLCELL_X8 FILLER_21_360 ();
 FILLCELL_X4 FILLER_21_368 ();
 FILLCELL_X2 FILLER_21_372 ();
 FILLCELL_X1 FILLER_21_374 ();
 FILLCELL_X1 FILLER_21_396 ();
 FILLCELL_X32 FILLER_21_404 ();
 FILLCELL_X16 FILLER_21_436 ();
 FILLCELL_X8 FILLER_21_452 ();
 FILLCELL_X4 FILLER_21_472 ();
 FILLCELL_X4 FILLER_21_483 ();
 FILLCELL_X2 FILLER_21_487 ();
 FILLCELL_X1 FILLER_21_496 ();
 FILLCELL_X8 FILLER_21_500 ();
 FILLCELL_X4 FILLER_21_508 ();
 FILLCELL_X2 FILLER_21_519 ();
 FILLCELL_X32 FILLER_21_524 ();
 FILLCELL_X32 FILLER_21_556 ();
 FILLCELL_X32 FILLER_21_588 ();
 FILLCELL_X32 FILLER_21_620 ();
 FILLCELL_X32 FILLER_21_652 ();
 FILLCELL_X32 FILLER_21_684 ();
 FILLCELL_X32 FILLER_21_716 ();
 FILLCELL_X32 FILLER_21_748 ();
 FILLCELL_X32 FILLER_21_780 ();
 FILLCELL_X32 FILLER_21_812 ();
 FILLCELL_X16 FILLER_21_844 ();
 FILLCELL_X2 FILLER_21_860 ();
 FILLCELL_X1 FILLER_21_862 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X16 FILLER_22_321 ();
 FILLCELL_X4 FILLER_22_337 ();
 FILLCELL_X1 FILLER_22_341 ();
 FILLCELL_X4 FILLER_22_349 ();
 FILLCELL_X1 FILLER_22_353 ();
 FILLCELL_X2 FILLER_22_368 ();
 FILLCELL_X1 FILLER_22_384 ();
 FILLCELL_X2 FILLER_22_392 ();
 FILLCELL_X1 FILLER_22_394 ();
 FILLCELL_X4 FILLER_22_402 ();
 FILLCELL_X32 FILLER_22_413 ();
 FILLCELL_X16 FILLER_22_445 ();
 FILLCELL_X8 FILLER_22_461 ();
 FILLCELL_X4 FILLER_22_469 ();
 FILLCELL_X1 FILLER_22_473 ();
 FILLCELL_X8 FILLER_22_477 ();
 FILLCELL_X8 FILLER_22_506 ();
 FILLCELL_X1 FILLER_22_514 ();
 FILLCELL_X16 FILLER_22_522 ();
 FILLCELL_X2 FILLER_22_538 ();
 FILLCELL_X1 FILLER_22_540 ();
 FILLCELL_X4 FILLER_22_558 ();
 FILLCELL_X32 FILLER_22_572 ();
 FILLCELL_X16 FILLER_22_604 ();
 FILLCELL_X8 FILLER_22_620 ();
 FILLCELL_X2 FILLER_22_628 ();
 FILLCELL_X1 FILLER_22_630 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X4 FILLER_22_856 ();
 FILLCELL_X2 FILLER_22_860 ();
 FILLCELL_X1 FILLER_22_862 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X16 FILLER_23_353 ();
 FILLCELL_X8 FILLER_23_369 ();
 FILLCELL_X2 FILLER_23_377 ();
 FILLCELL_X4 FILLER_23_400 ();
 FILLCELL_X1 FILLER_23_411 ();
 FILLCELL_X2 FILLER_23_419 ();
 FILLCELL_X2 FILLER_23_435 ();
 FILLCELL_X1 FILLER_23_437 ();
 FILLCELL_X8 FILLER_23_445 ();
 FILLCELL_X4 FILLER_23_453 ();
 FILLCELL_X2 FILLER_23_457 ();
 FILLCELL_X8 FILLER_23_473 ();
 FILLCELL_X2 FILLER_23_481 ();
 FILLCELL_X1 FILLER_23_483 ();
 FILLCELL_X4 FILLER_23_491 ();
 FILLCELL_X2 FILLER_23_495 ();
 FILLCELL_X16 FILLER_23_500 ();
 FILLCELL_X1 FILLER_23_516 ();
 FILLCELL_X8 FILLER_23_531 ();
 FILLCELL_X4 FILLER_23_539 ();
 FILLCELL_X2 FILLER_23_543 ();
 FILLCELL_X32 FILLER_23_552 ();
 FILLCELL_X32 FILLER_23_584 ();
 FILLCELL_X32 FILLER_23_616 ();
 FILLCELL_X32 FILLER_23_648 ();
 FILLCELL_X32 FILLER_23_680 ();
 FILLCELL_X32 FILLER_23_712 ();
 FILLCELL_X32 FILLER_23_744 ();
 FILLCELL_X32 FILLER_23_776 ();
 FILLCELL_X32 FILLER_23_808 ();
 FILLCELL_X16 FILLER_23_840 ();
 FILLCELL_X4 FILLER_23_856 ();
 FILLCELL_X2 FILLER_23_860 ();
 FILLCELL_X1 FILLER_23_862 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X16 FILLER_24_321 ();
 FILLCELL_X4 FILLER_24_337 ();
 FILLCELL_X32 FILLER_24_348 ();
 FILLCELL_X32 FILLER_24_380 ();
 FILLCELL_X16 FILLER_24_412 ();
 FILLCELL_X1 FILLER_24_428 ();
 FILLCELL_X32 FILLER_24_436 ();
 FILLCELL_X2 FILLER_24_468 ();
 FILLCELL_X1 FILLER_24_470 ();
 FILLCELL_X8 FILLER_24_478 ();
 FILLCELL_X4 FILLER_24_486 ();
 FILLCELL_X1 FILLER_24_490 ();
 FILLCELL_X8 FILLER_24_498 ();
 FILLCELL_X4 FILLER_24_506 ();
 FILLCELL_X2 FILLER_24_510 ();
 FILLCELL_X1 FILLER_24_512 ();
 FILLCELL_X4 FILLER_24_520 ();
 FILLCELL_X4 FILLER_24_531 ();
 FILLCELL_X2 FILLER_24_535 ();
 FILLCELL_X1 FILLER_24_537 ();
 FILLCELL_X2 FILLER_24_545 ();
 FILLCELL_X4 FILLER_24_554 ();
 FILLCELL_X32 FILLER_24_576 ();
 FILLCELL_X16 FILLER_24_608 ();
 FILLCELL_X4 FILLER_24_624 ();
 FILLCELL_X2 FILLER_24_628 ();
 FILLCELL_X1 FILLER_24_630 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X4 FILLER_24_856 ();
 FILLCELL_X2 FILLER_24_860 ();
 FILLCELL_X1 FILLER_24_862 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X8 FILLER_25_321 ();
 FILLCELL_X2 FILLER_25_329 ();
 FILLCELL_X2 FILLER_25_352 ();
 FILLCELL_X8 FILLER_25_400 ();
 FILLCELL_X2 FILLER_25_408 ();
 FILLCELL_X8 FILLER_25_417 ();
 FILLCELL_X4 FILLER_25_425 ();
 FILLCELL_X2 FILLER_25_436 ();
 FILLCELL_X1 FILLER_25_438 ();
 FILLCELL_X8 FILLER_25_446 ();
 FILLCELL_X2 FILLER_25_454 ();
 FILLCELL_X4 FILLER_25_463 ();
 FILLCELL_X32 FILLER_25_474 ();
 FILLCELL_X2 FILLER_25_506 ();
 FILLCELL_X16 FILLER_25_515 ();
 FILLCELL_X2 FILLER_25_531 ();
 FILLCELL_X1 FILLER_25_533 ();
 FILLCELL_X8 FILLER_25_548 ();
 FILLCELL_X2 FILLER_25_556 ();
 FILLCELL_X4 FILLER_25_565 ();
 FILLCELL_X2 FILLER_25_569 ();
 FILLCELL_X1 FILLER_25_571 ();
 FILLCELL_X32 FILLER_25_576 ();
 FILLCELL_X32 FILLER_25_608 ();
 FILLCELL_X32 FILLER_25_640 ();
 FILLCELL_X32 FILLER_25_672 ();
 FILLCELL_X32 FILLER_25_704 ();
 FILLCELL_X32 FILLER_25_736 ();
 FILLCELL_X32 FILLER_25_768 ();
 FILLCELL_X32 FILLER_25_800 ();
 FILLCELL_X16 FILLER_25_832 ();
 FILLCELL_X8 FILLER_25_848 ();
 FILLCELL_X4 FILLER_25_856 ();
 FILLCELL_X2 FILLER_25_860 ();
 FILLCELL_X1 FILLER_25_862 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X4 FILLER_26_321 ();
 FILLCELL_X2 FILLER_26_325 ();
 FILLCELL_X32 FILLER_26_341 ();
 FILLCELL_X1 FILLER_26_373 ();
 FILLCELL_X4 FILLER_26_381 ();
 FILLCELL_X2 FILLER_26_385 ();
 FILLCELL_X8 FILLER_26_394 ();
 FILLCELL_X2 FILLER_26_402 ();
 FILLCELL_X1 FILLER_26_411 ();
 FILLCELL_X8 FILLER_26_419 ();
 FILLCELL_X2 FILLER_26_427 ();
 FILLCELL_X1 FILLER_26_429 ();
 FILLCELL_X16 FILLER_26_437 ();
 FILLCELL_X2 FILLER_26_453 ();
 FILLCELL_X16 FILLER_26_462 ();
 FILLCELL_X1 FILLER_26_478 ();
 FILLCELL_X1 FILLER_26_486 ();
 FILLCELL_X4 FILLER_26_494 ();
 FILLCELL_X2 FILLER_26_498 ();
 FILLCELL_X32 FILLER_26_507 ();
 FILLCELL_X16 FILLER_26_539 ();
 FILLCELL_X1 FILLER_26_555 ();
 FILLCELL_X32 FILLER_26_563 ();
 FILLCELL_X32 FILLER_26_595 ();
 FILLCELL_X4 FILLER_26_627 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X4 FILLER_26_856 ();
 FILLCELL_X2 FILLER_26_860 ();
 FILLCELL_X1 FILLER_26_862 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X16 FILLER_27_289 ();
 FILLCELL_X4 FILLER_27_305 ();
 FILLCELL_X1 FILLER_27_309 ();
 FILLCELL_X8 FILLER_27_317 ();
 FILLCELL_X2 FILLER_27_325 ();
 FILLCELL_X2 FILLER_27_362 ();
 FILLCELL_X1 FILLER_27_364 ();
 FILLCELL_X4 FILLER_27_372 ();
 FILLCELL_X2 FILLER_27_376 ();
 FILLCELL_X1 FILLER_27_378 ();
 FILLCELL_X4 FILLER_27_386 ();
 FILLCELL_X2 FILLER_27_390 ();
 FILLCELL_X32 FILLER_27_399 ();
 FILLCELL_X4 FILLER_27_431 ();
 FILLCELL_X1 FILLER_27_435 ();
 FILLCELL_X16 FILLER_27_450 ();
 FILLCELL_X8 FILLER_27_466 ();
 FILLCELL_X2 FILLER_27_474 ();
 FILLCELL_X1 FILLER_27_476 ();
 FILLCELL_X4 FILLER_27_484 ();
 FILLCELL_X2 FILLER_27_488 ();
 FILLCELL_X4 FILLER_27_497 ();
 FILLCELL_X4 FILLER_27_508 ();
 FILLCELL_X1 FILLER_27_512 ();
 FILLCELL_X8 FILLER_27_534 ();
 FILLCELL_X2 FILLER_27_542 ();
 FILLCELL_X2 FILLER_27_562 ();
 FILLCELL_X32 FILLER_27_578 ();
 FILLCELL_X32 FILLER_27_610 ();
 FILLCELL_X32 FILLER_27_642 ();
 FILLCELL_X32 FILLER_27_674 ();
 FILLCELL_X32 FILLER_27_706 ();
 FILLCELL_X32 FILLER_27_738 ();
 FILLCELL_X32 FILLER_27_770 ();
 FILLCELL_X32 FILLER_27_802 ();
 FILLCELL_X16 FILLER_27_834 ();
 FILLCELL_X8 FILLER_27_850 ();
 FILLCELL_X4 FILLER_27_858 ();
 FILLCELL_X1 FILLER_27_862 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X16 FILLER_28_321 ();
 FILLCELL_X8 FILLER_28_337 ();
 FILLCELL_X2 FILLER_28_345 ();
 FILLCELL_X8 FILLER_28_354 ();
 FILLCELL_X1 FILLER_28_362 ();
 FILLCELL_X2 FILLER_28_384 ();
 FILLCELL_X1 FILLER_28_393 ();
 FILLCELL_X16 FILLER_28_401 ();
 FILLCELL_X2 FILLER_28_417 ();
 FILLCELL_X8 FILLER_28_426 ();
 FILLCELL_X2 FILLER_28_434 ();
 FILLCELL_X4 FILLER_28_443 ();
 FILLCELL_X8 FILLER_28_458 ();
 FILLCELL_X1 FILLER_28_466 ();
 FILLCELL_X16 FILLER_28_488 ();
 FILLCELL_X2 FILLER_28_504 ();
 FILLCELL_X8 FILLER_28_517 ();
 FILLCELL_X4 FILLER_28_525 ();
 FILLCELL_X1 FILLER_28_529 ();
 FILLCELL_X4 FILLER_28_537 ();
 FILLCELL_X1 FILLER_28_541 ();
 FILLCELL_X16 FILLER_28_554 ();
 FILLCELL_X4 FILLER_28_570 ();
 FILLCELL_X32 FILLER_28_588 ();
 FILLCELL_X8 FILLER_28_620 ();
 FILLCELL_X2 FILLER_28_628 ();
 FILLCELL_X1 FILLER_28_630 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X4 FILLER_28_856 ();
 FILLCELL_X2 FILLER_28_860 ();
 FILLCELL_X1 FILLER_28_862 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X8 FILLER_29_385 ();
 FILLCELL_X4 FILLER_29_393 ();
 FILLCELL_X2 FILLER_29_406 ();
 FILLCELL_X8 FILLER_29_424 ();
 FILLCELL_X4 FILLER_29_432 ();
 FILLCELL_X4 FILLER_29_465 ();
 FILLCELL_X16 FILLER_29_476 ();
 FILLCELL_X8 FILLER_29_492 ();
 FILLCELL_X2 FILLER_29_500 ();
 FILLCELL_X16 FILLER_29_516 ();
 FILLCELL_X8 FILLER_29_532 ();
 FILLCELL_X4 FILLER_29_540 ();
 FILLCELL_X2 FILLER_29_544 ();
 FILLCELL_X1 FILLER_29_546 ();
 FILLCELL_X16 FILLER_29_554 ();
 FILLCELL_X8 FILLER_29_570 ();
 FILLCELL_X2 FILLER_29_578 ();
 FILLCELL_X2 FILLER_29_584 ();
 FILLCELL_X1 FILLER_29_586 ();
 FILLCELL_X32 FILLER_29_589 ();
 FILLCELL_X32 FILLER_29_621 ();
 FILLCELL_X32 FILLER_29_653 ();
 FILLCELL_X32 FILLER_29_685 ();
 FILLCELL_X32 FILLER_29_717 ();
 FILLCELL_X32 FILLER_29_749 ();
 FILLCELL_X32 FILLER_29_781 ();
 FILLCELL_X32 FILLER_29_813 ();
 FILLCELL_X16 FILLER_29_845 ();
 FILLCELL_X2 FILLER_29_861 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X4 FILLER_30_353 ();
 FILLCELL_X2 FILLER_30_357 ();
 FILLCELL_X1 FILLER_30_359 ();
 FILLCELL_X32 FILLER_30_374 ();
 FILLCELL_X16 FILLER_30_406 ();
 FILLCELL_X1 FILLER_30_422 ();
 FILLCELL_X8 FILLER_30_430 ();
 FILLCELL_X8 FILLER_30_447 ();
 FILLCELL_X16 FILLER_30_472 ();
 FILLCELL_X2 FILLER_30_488 ();
 FILLCELL_X2 FILLER_30_530 ();
 FILLCELL_X1 FILLER_30_532 ();
 FILLCELL_X2 FILLER_30_540 ();
 FILLCELL_X1 FILLER_30_542 ();
 FILLCELL_X1 FILLER_30_556 ();
 FILLCELL_X8 FILLER_30_560 ();
 FILLCELL_X4 FILLER_30_568 ();
 FILLCELL_X1 FILLER_30_572 ();
 FILLCELL_X32 FILLER_30_580 ();
 FILLCELL_X16 FILLER_30_612 ();
 FILLCELL_X2 FILLER_30_628 ();
 FILLCELL_X1 FILLER_30_630 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X4 FILLER_30_856 ();
 FILLCELL_X2 FILLER_30_860 ();
 FILLCELL_X1 FILLER_30_862 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X8 FILLER_31_353 ();
 FILLCELL_X4 FILLER_31_361 ();
 FILLCELL_X2 FILLER_31_365 ();
 FILLCELL_X8 FILLER_31_374 ();
 FILLCELL_X1 FILLER_31_382 ();
 FILLCELL_X32 FILLER_31_390 ();
 FILLCELL_X32 FILLER_31_422 ();
 FILLCELL_X16 FILLER_31_454 ();
 FILLCELL_X32 FILLER_31_474 ();
 FILLCELL_X8 FILLER_31_506 ();
 FILLCELL_X2 FILLER_31_514 ();
 FILLCELL_X8 FILLER_31_519 ();
 FILLCELL_X8 FILLER_31_536 ();
 FILLCELL_X4 FILLER_31_544 ();
 FILLCELL_X1 FILLER_31_548 ();
 FILLCELL_X2 FILLER_31_556 ();
 FILLCELL_X1 FILLER_31_558 ();
 FILLCELL_X16 FILLER_31_563 ();
 FILLCELL_X2 FILLER_31_579 ();
 FILLCELL_X1 FILLER_31_581 ();
 FILLCELL_X32 FILLER_31_589 ();
 FILLCELL_X32 FILLER_31_621 ();
 FILLCELL_X32 FILLER_31_653 ();
 FILLCELL_X32 FILLER_31_685 ();
 FILLCELL_X32 FILLER_31_717 ();
 FILLCELL_X32 FILLER_31_749 ();
 FILLCELL_X32 FILLER_31_781 ();
 FILLCELL_X32 FILLER_31_813 ();
 FILLCELL_X16 FILLER_31_845 ();
 FILLCELL_X2 FILLER_31_861 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X8 FILLER_32_321 ();
 FILLCELL_X4 FILLER_32_329 ();
 FILLCELL_X2 FILLER_32_333 ();
 FILLCELL_X1 FILLER_32_335 ();
 FILLCELL_X2 FILLER_32_343 ();
 FILLCELL_X2 FILLER_32_366 ();
 FILLCELL_X2 FILLER_32_382 ();
 FILLCELL_X1 FILLER_32_384 ();
 FILLCELL_X1 FILLER_32_392 ();
 FILLCELL_X2 FILLER_32_400 ();
 FILLCELL_X1 FILLER_32_402 ();
 FILLCELL_X1 FILLER_32_410 ();
 FILLCELL_X4 FILLER_32_418 ();
 FILLCELL_X4 FILLER_32_429 ();
 FILLCELL_X2 FILLER_32_433 ();
 FILLCELL_X1 FILLER_32_435 ();
 FILLCELL_X8 FILLER_32_454 ();
 FILLCELL_X4 FILLER_32_462 ();
 FILLCELL_X1 FILLER_32_478 ();
 FILLCELL_X4 FILLER_32_486 ();
 FILLCELL_X2 FILLER_32_490 ();
 FILLCELL_X1 FILLER_32_492 ();
 FILLCELL_X16 FILLER_32_500 ();
 FILLCELL_X1 FILLER_32_516 ();
 FILLCELL_X16 FILLER_32_524 ();
 FILLCELL_X2 FILLER_32_540 ();
 FILLCELL_X8 FILLER_32_546 ();
 FILLCELL_X4 FILLER_32_554 ();
 FILLCELL_X1 FILLER_32_558 ();
 FILLCELL_X4 FILLER_32_569 ();
 FILLCELL_X2 FILLER_32_573 ();
 FILLCELL_X32 FILLER_32_578 ();
 FILLCELL_X16 FILLER_32_610 ();
 FILLCELL_X4 FILLER_32_626 ();
 FILLCELL_X1 FILLER_32_630 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X4 FILLER_32_856 ();
 FILLCELL_X2 FILLER_32_860 ();
 FILLCELL_X1 FILLER_32_862 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X2 FILLER_33_321 ();
 FILLCELL_X1 FILLER_33_323 ();
 FILLCELL_X8 FILLER_33_331 ();
 FILLCELL_X2 FILLER_33_339 ();
 FILLCELL_X1 FILLER_33_341 ();
 FILLCELL_X2 FILLER_33_349 ();
 FILLCELL_X2 FILLER_33_365 ();
 FILLCELL_X2 FILLER_33_374 ();
 FILLCELL_X1 FILLER_33_376 ();
 FILLCELL_X4 FILLER_33_384 ();
 FILLCELL_X1 FILLER_33_388 ();
 FILLCELL_X4 FILLER_33_396 ();
 FILLCELL_X1 FILLER_33_400 ();
 FILLCELL_X2 FILLER_33_408 ();
 FILLCELL_X16 FILLER_33_417 ();
 FILLCELL_X8 FILLER_33_433 ();
 FILLCELL_X4 FILLER_33_441 ();
 FILLCELL_X2 FILLER_33_445 ();
 FILLCELL_X1 FILLER_33_447 ();
 FILLCELL_X16 FILLER_33_452 ();
 FILLCELL_X1 FILLER_33_468 ();
 FILLCELL_X8 FILLER_33_480 ();
 FILLCELL_X2 FILLER_33_488 ();
 FILLCELL_X1 FILLER_33_490 ();
 FILLCELL_X2 FILLER_33_498 ();
 FILLCELL_X2 FILLER_33_504 ();
 FILLCELL_X8 FILLER_33_511 ();
 FILLCELL_X2 FILLER_33_519 ();
 FILLCELL_X8 FILLER_33_535 ();
 FILLCELL_X4 FILLER_33_543 ();
 FILLCELL_X2 FILLER_33_554 ();
 FILLCELL_X1 FILLER_33_556 ();
 FILLCELL_X4 FILLER_33_568 ();
 FILLCELL_X2 FILLER_33_572 ();
 FILLCELL_X1 FILLER_33_581 ();
 FILLCELL_X32 FILLER_33_585 ();
 FILLCELL_X32 FILLER_33_617 ();
 FILLCELL_X32 FILLER_33_649 ();
 FILLCELL_X32 FILLER_33_681 ();
 FILLCELL_X32 FILLER_33_713 ();
 FILLCELL_X32 FILLER_33_745 ();
 FILLCELL_X32 FILLER_33_777 ();
 FILLCELL_X32 FILLER_33_809 ();
 FILLCELL_X16 FILLER_33_841 ();
 FILLCELL_X4 FILLER_33_857 ();
 FILLCELL_X2 FILLER_33_861 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X16 FILLER_34_289 ();
 FILLCELL_X8 FILLER_34_305 ();
 FILLCELL_X2 FILLER_34_320 ();
 FILLCELL_X2 FILLER_34_329 ();
 FILLCELL_X32 FILLER_34_345 ();
 FILLCELL_X32 FILLER_34_377 ();
 FILLCELL_X16 FILLER_34_409 ();
 FILLCELL_X8 FILLER_34_425 ();
 FILLCELL_X1 FILLER_34_433 ();
 FILLCELL_X32 FILLER_34_456 ();
 FILLCELL_X16 FILLER_34_488 ();
 FILLCELL_X4 FILLER_34_504 ();
 FILLCELL_X8 FILLER_34_510 ();
 FILLCELL_X4 FILLER_34_518 ();
 FILLCELL_X8 FILLER_34_540 ();
 FILLCELL_X1 FILLER_34_548 ();
 FILLCELL_X2 FILLER_34_558 ();
 FILLCELL_X1 FILLER_34_567 ();
 FILLCELL_X4 FILLER_34_570 ();
 FILLCELL_X1 FILLER_34_574 ();
 FILLCELL_X32 FILLER_34_582 ();
 FILLCELL_X16 FILLER_34_614 ();
 FILLCELL_X1 FILLER_34_630 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X4 FILLER_34_856 ();
 FILLCELL_X2 FILLER_34_860 ();
 FILLCELL_X1 FILLER_34_862 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X2 FILLER_35_289 ();
 FILLCELL_X1 FILLER_35_291 ();
 FILLCELL_X4 FILLER_35_341 ();
 FILLCELL_X4 FILLER_35_352 ();
 FILLCELL_X2 FILLER_35_356 ();
 FILLCELL_X32 FILLER_35_365 ();
 FILLCELL_X16 FILLER_35_397 ();
 FILLCELL_X4 FILLER_35_413 ();
 FILLCELL_X2 FILLER_35_417 ();
 FILLCELL_X16 FILLER_35_426 ();
 FILLCELL_X2 FILLER_35_442 ();
 FILLCELL_X2 FILLER_35_457 ();
 FILLCELL_X1 FILLER_35_459 ();
 FILLCELL_X32 FILLER_35_474 ();
 FILLCELL_X4 FILLER_35_506 ();
 FILLCELL_X2 FILLER_35_510 ();
 FILLCELL_X1 FILLER_35_512 ();
 FILLCELL_X8 FILLER_35_518 ();
 FILLCELL_X4 FILLER_35_526 ();
 FILLCELL_X2 FILLER_35_530 ();
 FILLCELL_X1 FILLER_35_536 ();
 FILLCELL_X2 FILLER_35_545 ();
 FILLCELL_X1 FILLER_35_547 ();
 FILLCELL_X2 FILLER_35_557 ();
 FILLCELL_X1 FILLER_35_559 ();
 FILLCELL_X32 FILLER_35_569 ();
 FILLCELL_X32 FILLER_35_601 ();
 FILLCELL_X32 FILLER_35_633 ();
 FILLCELL_X32 FILLER_35_665 ();
 FILLCELL_X32 FILLER_35_697 ();
 FILLCELL_X32 FILLER_35_729 ();
 FILLCELL_X32 FILLER_35_761 ();
 FILLCELL_X32 FILLER_35_793 ();
 FILLCELL_X32 FILLER_35_825 ();
 FILLCELL_X4 FILLER_35_857 ();
 FILLCELL_X2 FILLER_35_861 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X16 FILLER_36_289 ();
 FILLCELL_X8 FILLER_36_305 ();
 FILLCELL_X2 FILLER_36_313 ();
 FILLCELL_X4 FILLER_36_353 ();
 FILLCELL_X2 FILLER_36_357 ();
 FILLCELL_X32 FILLER_36_373 ();
 FILLCELL_X8 FILLER_36_405 ();
 FILLCELL_X4 FILLER_36_420 ();
 FILLCELL_X2 FILLER_36_424 ();
 FILLCELL_X2 FILLER_36_433 ();
 FILLCELL_X2 FILLER_36_440 ();
 FILLCELL_X16 FILLER_36_451 ();
 FILLCELL_X8 FILLER_36_467 ();
 FILLCELL_X4 FILLER_36_475 ();
 FILLCELL_X2 FILLER_36_486 ();
 FILLCELL_X8 FILLER_36_495 ();
 FILLCELL_X2 FILLER_36_503 ();
 FILLCELL_X2 FILLER_36_512 ();
 FILLCELL_X1 FILLER_36_514 ();
 FILLCELL_X4 FILLER_36_522 ();
 FILLCELL_X2 FILLER_36_526 ();
 FILLCELL_X1 FILLER_36_528 ();
 FILLCELL_X2 FILLER_36_532 ();
 FILLCELL_X4 FILLER_36_537 ();
 FILLCELL_X2 FILLER_36_541 ();
 FILLCELL_X1 FILLER_36_543 ();
 FILLCELL_X2 FILLER_36_548 ();
 FILLCELL_X2 FILLER_36_560 ();
 FILLCELL_X4 FILLER_36_571 ();
 FILLCELL_X4 FILLER_36_586 ();
 FILLCELL_X32 FILLER_36_597 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X4 FILLER_36_856 ();
 FILLCELL_X2 FILLER_36_860 ();
 FILLCELL_X1 FILLER_36_862 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X16 FILLER_37_289 ();
 FILLCELL_X8 FILLER_37_305 ();
 FILLCELL_X8 FILLER_37_320 ();
 FILLCELL_X1 FILLER_37_328 ();
 FILLCELL_X32 FILLER_37_343 ();
 FILLCELL_X4 FILLER_37_375 ();
 FILLCELL_X2 FILLER_37_379 ();
 FILLCELL_X8 FILLER_37_402 ();
 FILLCELL_X2 FILLER_37_410 ();
 FILLCELL_X8 FILLER_37_437 ();
 FILLCELL_X1 FILLER_37_445 ();
 FILLCELL_X16 FILLER_37_448 ();
 FILLCELL_X1 FILLER_37_464 ();
 FILLCELL_X4 FILLER_37_467 ();
 FILLCELL_X16 FILLER_37_475 ();
 FILLCELL_X8 FILLER_37_491 ();
 FILLCELL_X4 FILLER_37_499 ();
 FILLCELL_X2 FILLER_37_503 ();
 FILLCELL_X2 FILLER_37_509 ();
 FILLCELL_X4 FILLER_37_518 ();
 FILLCELL_X2 FILLER_37_522 ();
 FILLCELL_X2 FILLER_37_542 ();
 FILLCELL_X16 FILLER_37_556 ();
 FILLCELL_X4 FILLER_37_572 ();
 FILLCELL_X2 FILLER_37_579 ();
 FILLCELL_X1 FILLER_37_581 ();
 FILLCELL_X32 FILLER_37_585 ();
 FILLCELL_X32 FILLER_37_617 ();
 FILLCELL_X32 FILLER_37_649 ();
 FILLCELL_X32 FILLER_37_681 ();
 FILLCELL_X32 FILLER_37_713 ();
 FILLCELL_X32 FILLER_37_745 ();
 FILLCELL_X32 FILLER_37_777 ();
 FILLCELL_X32 FILLER_37_809 ();
 FILLCELL_X16 FILLER_37_841 ();
 FILLCELL_X4 FILLER_37_857 ();
 FILLCELL_X2 FILLER_37_861 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X16 FILLER_38_289 ();
 FILLCELL_X4 FILLER_38_305 ();
 FILLCELL_X2 FILLER_38_309 ();
 FILLCELL_X1 FILLER_38_311 ();
 FILLCELL_X4 FILLER_38_319 ();
 FILLCELL_X2 FILLER_38_323 ();
 FILLCELL_X2 FILLER_38_339 ();
 FILLCELL_X16 FILLER_38_350 ();
 FILLCELL_X8 FILLER_38_366 ();
 FILLCELL_X4 FILLER_38_374 ();
 FILLCELL_X1 FILLER_38_378 ();
 FILLCELL_X16 FILLER_38_386 ();
 FILLCELL_X1 FILLER_38_402 ();
 FILLCELL_X4 FILLER_38_424 ();
 FILLCELL_X2 FILLER_38_428 ();
 FILLCELL_X1 FILLER_38_430 ();
 FILLCELL_X8 FILLER_38_435 ();
 FILLCELL_X4 FILLER_38_443 ();
 FILLCELL_X1 FILLER_38_447 ();
 FILLCELL_X8 FILLER_38_455 ();
 FILLCELL_X32 FILLER_38_472 ();
 FILLCELL_X8 FILLER_38_504 ();
 FILLCELL_X4 FILLER_38_515 ();
 FILLCELL_X2 FILLER_38_519 ();
 FILLCELL_X1 FILLER_38_521 ();
 FILLCELL_X4 FILLER_38_534 ();
 FILLCELL_X1 FILLER_38_538 ();
 FILLCELL_X4 FILLER_38_544 ();
 FILLCELL_X2 FILLER_38_548 ();
 FILLCELL_X2 FILLER_38_559 ();
 FILLCELL_X1 FILLER_38_561 ();
 FILLCELL_X4 FILLER_38_569 ();
 FILLCELL_X32 FILLER_38_580 ();
 FILLCELL_X16 FILLER_38_612 ();
 FILLCELL_X2 FILLER_38_628 ();
 FILLCELL_X1 FILLER_38_630 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X4 FILLER_38_856 ();
 FILLCELL_X2 FILLER_38_860 ();
 FILLCELL_X1 FILLER_38_862 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X4 FILLER_39_289 ();
 FILLCELL_X1 FILLER_39_293 ();
 FILLCELL_X4 FILLER_39_307 ();
 FILLCELL_X2 FILLER_39_318 ();
 FILLCELL_X1 FILLER_39_320 ();
 FILLCELL_X16 FILLER_39_328 ();
 FILLCELL_X4 FILLER_39_344 ();
 FILLCELL_X1 FILLER_39_348 ();
 FILLCELL_X8 FILLER_39_356 ();
 FILLCELL_X4 FILLER_39_364 ();
 FILLCELL_X1 FILLER_39_368 ();
 FILLCELL_X4 FILLER_39_376 ();
 FILLCELL_X16 FILLER_39_385 ();
 FILLCELL_X8 FILLER_39_401 ();
 FILLCELL_X4 FILLER_39_409 ();
 FILLCELL_X2 FILLER_39_420 ();
 FILLCELL_X4 FILLER_39_451 ();
 FILLCELL_X2 FILLER_39_455 ();
 FILLCELL_X1 FILLER_39_457 ();
 FILLCELL_X8 FILLER_39_464 ();
 FILLCELL_X4 FILLER_39_472 ();
 FILLCELL_X2 FILLER_39_476 ();
 FILLCELL_X1 FILLER_39_478 ();
 FILLCELL_X1 FILLER_39_483 ();
 FILLCELL_X4 FILLER_39_488 ();
 FILLCELL_X1 FILLER_39_496 ();
 FILLCELL_X4 FILLER_39_508 ();
 FILLCELL_X1 FILLER_39_512 ();
 FILLCELL_X2 FILLER_39_520 ();
 FILLCELL_X4 FILLER_39_536 ();
 FILLCELL_X8 FILLER_39_547 ();
 FILLCELL_X8 FILLER_39_558 ();
 FILLCELL_X2 FILLER_39_566 ();
 FILLCELL_X1 FILLER_39_568 ();
 FILLCELL_X1 FILLER_39_571 ();
 FILLCELL_X8 FILLER_39_575 ();
 FILLCELL_X4 FILLER_39_583 ();
 FILLCELL_X32 FILLER_39_595 ();
 FILLCELL_X32 FILLER_39_627 ();
 FILLCELL_X32 FILLER_39_659 ();
 FILLCELL_X32 FILLER_39_691 ();
 FILLCELL_X32 FILLER_39_723 ();
 FILLCELL_X32 FILLER_39_755 ();
 FILLCELL_X32 FILLER_39_787 ();
 FILLCELL_X32 FILLER_39_819 ();
 FILLCELL_X8 FILLER_39_851 ();
 FILLCELL_X4 FILLER_39_859 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X16 FILLER_40_257 ();
 FILLCELL_X8 FILLER_40_273 ();
 FILLCELL_X4 FILLER_40_281 ();
 FILLCELL_X4 FILLER_40_311 ();
 FILLCELL_X1 FILLER_40_315 ();
 FILLCELL_X8 FILLER_40_332 ();
 FILLCELL_X1 FILLER_40_340 ();
 FILLCELL_X32 FILLER_40_369 ();
 FILLCELL_X16 FILLER_40_401 ();
 FILLCELL_X8 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_428 ();
 FILLCELL_X2 FILLER_40_460 ();
 FILLCELL_X1 FILLER_40_462 ();
 FILLCELL_X8 FILLER_40_466 ();
 FILLCELL_X4 FILLER_40_502 ();
 FILLCELL_X2 FILLER_40_506 ();
 FILLCELL_X1 FILLER_40_508 ();
 FILLCELL_X4 FILLER_40_513 ();
 FILLCELL_X2 FILLER_40_517 ();
 FILLCELL_X1 FILLER_40_524 ();
 FILLCELL_X1 FILLER_40_540 ();
 FILLCELL_X2 FILLER_40_547 ();
 FILLCELL_X8 FILLER_40_556 ();
 FILLCELL_X4 FILLER_40_564 ();
 FILLCELL_X2 FILLER_40_568 ();
 FILLCELL_X1 FILLER_40_584 ();
 FILLCELL_X1 FILLER_40_592 ();
 FILLCELL_X32 FILLER_40_597 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X4 FILLER_40_856 ();
 FILLCELL_X2 FILLER_40_860 ();
 FILLCELL_X1 FILLER_40_862 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X16 FILLER_41_289 ();
 FILLCELL_X4 FILLER_41_305 ();
 FILLCELL_X2 FILLER_41_330 ();
 FILLCELL_X16 FILLER_41_339 ();
 FILLCELL_X8 FILLER_41_355 ();
 FILLCELL_X1 FILLER_41_377 ();
 FILLCELL_X8 FILLER_41_392 ();
 FILLCELL_X4 FILLER_41_400 ();
 FILLCELL_X2 FILLER_41_404 ();
 FILLCELL_X8 FILLER_41_427 ();
 FILLCELL_X2 FILLER_41_435 ();
 FILLCELL_X1 FILLER_41_437 ();
 FILLCELL_X16 FILLER_41_441 ();
 FILLCELL_X2 FILLER_41_457 ();
 FILLCELL_X4 FILLER_41_470 ();
 FILLCELL_X2 FILLER_41_474 ();
 FILLCELL_X2 FILLER_41_513 ();
 FILLCELL_X1 FILLER_41_515 ();
 FILLCELL_X4 FILLER_41_519 ();
 FILLCELL_X2 FILLER_41_523 ();
 FILLCELL_X1 FILLER_41_536 ();
 FILLCELL_X2 FILLER_41_541 ();
 FILLCELL_X2 FILLER_41_550 ();
 FILLCELL_X1 FILLER_41_552 ();
 FILLCELL_X8 FILLER_41_564 ();
 FILLCELL_X1 FILLER_41_572 ();
 FILLCELL_X2 FILLER_41_576 ();
 FILLCELL_X1 FILLER_41_578 ();
 FILLCELL_X32 FILLER_41_603 ();
 FILLCELL_X32 FILLER_41_635 ();
 FILLCELL_X32 FILLER_41_667 ();
 FILLCELL_X32 FILLER_41_699 ();
 FILLCELL_X32 FILLER_41_731 ();
 FILLCELL_X32 FILLER_41_763 ();
 FILLCELL_X32 FILLER_41_795 ();
 FILLCELL_X32 FILLER_41_827 ();
 FILLCELL_X4 FILLER_41_859 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X16 FILLER_42_257 ();
 FILLCELL_X8 FILLER_42_273 ();
 FILLCELL_X2 FILLER_42_281 ();
 FILLCELL_X16 FILLER_42_330 ();
 FILLCELL_X4 FILLER_42_353 ();
 FILLCELL_X8 FILLER_42_378 ();
 FILLCELL_X4 FILLER_42_386 ();
 FILLCELL_X1 FILLER_42_390 ();
 FILLCELL_X16 FILLER_42_398 ();
 FILLCELL_X4 FILLER_42_414 ();
 FILLCELL_X4 FILLER_42_421 ();
 FILLCELL_X2 FILLER_42_425 ();
 FILLCELL_X2 FILLER_42_438 ();
 FILLCELL_X4 FILLER_42_454 ();
 FILLCELL_X2 FILLER_42_458 ();
 FILLCELL_X4 FILLER_42_470 ();
 FILLCELL_X4 FILLER_42_478 ();
 FILLCELL_X8 FILLER_42_489 ();
 FILLCELL_X4 FILLER_42_497 ();
 FILLCELL_X2 FILLER_42_501 ();
 FILLCELL_X4 FILLER_42_506 ();
 FILLCELL_X2 FILLER_42_510 ();
 FILLCELL_X8 FILLER_42_552 ();
 FILLCELL_X4 FILLER_42_560 ();
 FILLCELL_X1 FILLER_42_564 ();
 FILLCELL_X4 FILLER_42_572 ();
 FILLCELL_X2 FILLER_42_576 ();
 FILLCELL_X1 FILLER_42_578 ();
 FILLCELL_X32 FILLER_42_594 ();
 FILLCELL_X4 FILLER_42_626 ();
 FILLCELL_X1 FILLER_42_630 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X4 FILLER_42_856 ();
 FILLCELL_X2 FILLER_42_860 ();
 FILLCELL_X1 FILLER_42_862 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X4 FILLER_43_289 ();
 FILLCELL_X1 FILLER_43_293 ();
 FILLCELL_X4 FILLER_43_310 ();
 FILLCELL_X2 FILLER_43_314 ();
 FILLCELL_X1 FILLER_43_316 ();
 FILLCELL_X8 FILLER_43_338 ();
 FILLCELL_X2 FILLER_43_346 ();
 FILLCELL_X4 FILLER_43_376 ();
 FILLCELL_X2 FILLER_43_380 ();
 FILLCELL_X16 FILLER_43_389 ();
 FILLCELL_X2 FILLER_43_405 ();
 FILLCELL_X8 FILLER_43_414 ();
 FILLCELL_X4 FILLER_43_422 ();
 FILLCELL_X16 FILLER_43_444 ();
 FILLCELL_X2 FILLER_43_460 ();
 FILLCELL_X1 FILLER_43_462 ();
 FILLCELL_X8 FILLER_43_468 ();
 FILLCELL_X2 FILLER_43_476 ();
 FILLCELL_X1 FILLER_43_478 ();
 FILLCELL_X4 FILLER_43_497 ();
 FILLCELL_X4 FILLER_43_504 ();
 FILLCELL_X4 FILLER_43_519 ();
 FILLCELL_X2 FILLER_43_523 ();
 FILLCELL_X1 FILLER_43_525 ();
 FILLCELL_X2 FILLER_43_548 ();
 FILLCELL_X16 FILLER_43_558 ();
 FILLCELL_X8 FILLER_43_574 ();
 FILLCELL_X4 FILLER_43_582 ();
 FILLCELL_X1 FILLER_43_586 ();
 FILLCELL_X32 FILLER_43_591 ();
 FILLCELL_X32 FILLER_43_623 ();
 FILLCELL_X32 FILLER_43_655 ();
 FILLCELL_X32 FILLER_43_687 ();
 FILLCELL_X32 FILLER_43_719 ();
 FILLCELL_X32 FILLER_43_751 ();
 FILLCELL_X32 FILLER_43_783 ();
 FILLCELL_X8 FILLER_43_815 ();
 FILLCELL_X1 FILLER_43_823 ();
 FILLCELL_X32 FILLER_43_827 ();
 FILLCELL_X4 FILLER_43_859 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X16 FILLER_44_289 ();
 FILLCELL_X4 FILLER_44_305 ();
 FILLCELL_X2 FILLER_44_309 ();
 FILLCELL_X8 FILLER_44_325 ();
 FILLCELL_X4 FILLER_44_333 ();
 FILLCELL_X4 FILLER_44_344 ();
 FILLCELL_X2 FILLER_44_348 ();
 FILLCELL_X1 FILLER_44_350 ();
 FILLCELL_X2 FILLER_44_367 ();
 FILLCELL_X4 FILLER_44_383 ();
 FILLCELL_X8 FILLER_44_401 ();
 FILLCELL_X4 FILLER_44_409 ();
 FILLCELL_X1 FILLER_44_413 ();
 FILLCELL_X4 FILLER_44_421 ();
 FILLCELL_X2 FILLER_44_425 ();
 FILLCELL_X1 FILLER_44_427 ();
 FILLCELL_X4 FILLER_44_438 ();
 FILLCELL_X2 FILLER_44_442 ();
 FILLCELL_X1 FILLER_44_444 ();
 FILLCELL_X4 FILLER_44_456 ();
 FILLCELL_X1 FILLER_44_460 ();
 FILLCELL_X4 FILLER_44_466 ();
 FILLCELL_X16 FILLER_44_490 ();
 FILLCELL_X4 FILLER_44_517 ();
 FILLCELL_X1 FILLER_44_521 ();
 FILLCELL_X8 FILLER_44_525 ();
 FILLCELL_X4 FILLER_44_533 ();
 FILLCELL_X1 FILLER_44_537 ();
 FILLCELL_X4 FILLER_44_541 ();
 FILLCELL_X1 FILLER_44_545 ();
 FILLCELL_X4 FILLER_44_564 ();
 FILLCELL_X2 FILLER_44_568 ();
 FILLCELL_X1 FILLER_44_570 ();
 FILLCELL_X4 FILLER_44_578 ();
 FILLCELL_X2 FILLER_44_582 ();
 FILLCELL_X1 FILLER_44_584 ();
 FILLCELL_X32 FILLER_44_591 ();
 FILLCELL_X8 FILLER_44_623 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X4 FILLER_44_856 ();
 FILLCELL_X2 FILLER_44_860 ();
 FILLCELL_X1 FILLER_44_862 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X16 FILLER_45_289 ();
 FILLCELL_X8 FILLER_45_305 ();
 FILLCELL_X4 FILLER_45_313 ();
 FILLCELL_X2 FILLER_45_317 ();
 FILLCELL_X1 FILLER_45_319 ();
 FILLCELL_X1 FILLER_45_334 ();
 FILLCELL_X1 FILLER_45_349 ();
 FILLCELL_X1 FILLER_45_363 ();
 FILLCELL_X8 FILLER_45_371 ();
 FILLCELL_X4 FILLER_45_379 ();
 FILLCELL_X2 FILLER_45_383 ();
 FILLCELL_X1 FILLER_45_385 ();
 FILLCELL_X16 FILLER_45_393 ();
 FILLCELL_X4 FILLER_45_409 ();
 FILLCELL_X2 FILLER_45_413 ();
 FILLCELL_X1 FILLER_45_415 ();
 FILLCELL_X8 FILLER_45_425 ();
 FILLCELL_X2 FILLER_45_433 ();
 FILLCELL_X1 FILLER_45_435 ();
 FILLCELL_X2 FILLER_45_445 ();
 FILLCELL_X8 FILLER_45_454 ();
 FILLCELL_X4 FILLER_45_462 ();
 FILLCELL_X4 FILLER_45_482 ();
 FILLCELL_X2 FILLER_45_486 ();
 FILLCELL_X1 FILLER_45_488 ();
 FILLCELL_X32 FILLER_45_500 ();
 FILLCELL_X8 FILLER_45_532 ();
 FILLCELL_X2 FILLER_45_540 ();
 FILLCELL_X1 FILLER_45_542 ();
 FILLCELL_X4 FILLER_45_549 ();
 FILLCELL_X1 FILLER_45_553 ();
 FILLCELL_X32 FILLER_45_557 ();
 FILLCELL_X32 FILLER_45_589 ();
 FILLCELL_X32 FILLER_45_621 ();
 FILLCELL_X32 FILLER_45_653 ();
 FILLCELL_X32 FILLER_45_685 ();
 FILLCELL_X32 FILLER_45_717 ();
 FILLCELL_X32 FILLER_45_749 ();
 FILLCELL_X32 FILLER_45_781 ();
 FILLCELL_X32 FILLER_45_813 ();
 FILLCELL_X16 FILLER_45_845 ();
 FILLCELL_X2 FILLER_45_861 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X16 FILLER_46_289 ();
 FILLCELL_X4 FILLER_46_305 ();
 FILLCELL_X2 FILLER_46_309 ();
 FILLCELL_X1 FILLER_46_311 ();
 FILLCELL_X16 FILLER_46_328 ();
 FILLCELL_X8 FILLER_46_344 ();
 FILLCELL_X4 FILLER_46_352 ();
 FILLCELL_X2 FILLER_46_356 ();
 FILLCELL_X1 FILLER_46_358 ();
 FILLCELL_X8 FILLER_46_366 ();
 FILLCELL_X4 FILLER_46_374 ();
 FILLCELL_X2 FILLER_46_378 ();
 FILLCELL_X16 FILLER_46_387 ();
 FILLCELL_X8 FILLER_46_403 ();
 FILLCELL_X4 FILLER_46_411 ();
 FILLCELL_X1 FILLER_46_415 ();
 FILLCELL_X8 FILLER_46_423 ();
 FILLCELL_X2 FILLER_46_431 ();
 FILLCELL_X1 FILLER_46_433 ();
 FILLCELL_X8 FILLER_46_441 ();
 FILLCELL_X2 FILLER_46_449 ();
 FILLCELL_X4 FILLER_46_454 ();
 FILLCELL_X2 FILLER_46_458 ();
 FILLCELL_X2 FILLER_46_465 ();
 FILLCELL_X8 FILLER_46_472 ();
 FILLCELL_X2 FILLER_46_511 ();
 FILLCELL_X2 FILLER_46_524 ();
 FILLCELL_X2 FILLER_46_533 ();
 FILLCELL_X4 FILLER_46_549 ();
 FILLCELL_X1 FILLER_46_582 ();
 FILLCELL_X32 FILLER_46_586 ();
 FILLCELL_X8 FILLER_46_618 ();
 FILLCELL_X4 FILLER_46_626 ();
 FILLCELL_X1 FILLER_46_630 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X16 FILLER_46_824 ();
 FILLCELL_X8 FILLER_46_840 ();
 FILLCELL_X4 FILLER_46_848 ();
 FILLCELL_X2 FILLER_46_852 ();
 FILLCELL_X1 FILLER_46_854 ();
 FILLCELL_X4 FILLER_46_858 ();
 FILLCELL_X1 FILLER_46_862 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X8 FILLER_47_289 ();
 FILLCELL_X4 FILLER_47_297 ();
 FILLCELL_X8 FILLER_47_308 ();
 FILLCELL_X1 FILLER_47_316 ();
 FILLCELL_X8 FILLER_47_324 ();
 FILLCELL_X1 FILLER_47_332 ();
 FILLCELL_X16 FILLER_47_340 ();
 FILLCELL_X8 FILLER_47_370 ();
 FILLCELL_X4 FILLER_47_378 ();
 FILLCELL_X2 FILLER_47_382 ();
 FILLCELL_X4 FILLER_47_398 ();
 FILLCELL_X2 FILLER_47_402 ();
 FILLCELL_X1 FILLER_47_404 ();
 FILLCELL_X2 FILLER_47_412 ();
 FILLCELL_X2 FILLER_47_418 ();
 FILLCELL_X32 FILLER_47_427 ();
 FILLCELL_X8 FILLER_47_459 ();
 FILLCELL_X4 FILLER_47_467 ();
 FILLCELL_X2 FILLER_47_471 ();
 FILLCELL_X8 FILLER_47_478 ();
 FILLCELL_X2 FILLER_47_486 ();
 FILLCELL_X4 FILLER_47_499 ();
 FILLCELL_X2 FILLER_47_503 ();
 FILLCELL_X2 FILLER_47_512 ();
 FILLCELL_X2 FILLER_47_539 ();
 FILLCELL_X1 FILLER_47_541 ();
 FILLCELL_X2 FILLER_47_561 ();
 FILLCELL_X16 FILLER_47_570 ();
 FILLCELL_X1 FILLER_47_586 ();
 FILLCELL_X2 FILLER_47_592 ();
 FILLCELL_X1 FILLER_47_594 ();
 FILLCELL_X32 FILLER_47_599 ();
 FILLCELL_X32 FILLER_47_631 ();
 FILLCELL_X32 FILLER_47_663 ();
 FILLCELL_X32 FILLER_47_695 ();
 FILLCELL_X32 FILLER_47_727 ();
 FILLCELL_X32 FILLER_47_759 ();
 FILLCELL_X32 FILLER_47_791 ();
 FILLCELL_X32 FILLER_47_823 ();
 FILLCELL_X8 FILLER_47_855 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X8 FILLER_48_289 ();
 FILLCELL_X2 FILLER_48_297 ();
 FILLCELL_X4 FILLER_48_313 ();
 FILLCELL_X1 FILLER_48_317 ();
 FILLCELL_X16 FILLER_48_339 ();
 FILLCELL_X8 FILLER_48_355 ();
 FILLCELL_X4 FILLER_48_363 ();
 FILLCELL_X1 FILLER_48_367 ();
 FILLCELL_X4 FILLER_48_375 ();
 FILLCELL_X32 FILLER_48_386 ();
 FILLCELL_X16 FILLER_48_418 ();
 FILLCELL_X4 FILLER_48_434 ();
 FILLCELL_X1 FILLER_48_438 ();
 FILLCELL_X1 FILLER_48_443 ();
 FILLCELL_X8 FILLER_48_452 ();
 FILLCELL_X2 FILLER_48_460 ();
 FILLCELL_X1 FILLER_48_462 ();
 FILLCELL_X8 FILLER_48_474 ();
 FILLCELL_X4 FILLER_48_484 ();
 FILLCELL_X1 FILLER_48_488 ();
 FILLCELL_X4 FILLER_48_500 ();
 FILLCELL_X1 FILLER_48_504 ();
 FILLCELL_X2 FILLER_48_518 ();
 FILLCELL_X1 FILLER_48_520 ();
 FILLCELL_X2 FILLER_48_547 ();
 FILLCELL_X8 FILLER_48_551 ();
 FILLCELL_X4 FILLER_48_559 ();
 FILLCELL_X2 FILLER_48_580 ();
 FILLCELL_X1 FILLER_48_582 ();
 FILLCELL_X16 FILLER_48_612 ();
 FILLCELL_X2 FILLER_48_628 ();
 FILLCELL_X1 FILLER_48_630 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_827 ();
 FILLCELL_X4 FILLER_48_859 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X8 FILLER_49_289 ();
 FILLCELL_X4 FILLER_49_297 ();
 FILLCELL_X2 FILLER_49_301 ();
 FILLCELL_X2 FILLER_49_310 ();
 FILLCELL_X2 FILLER_49_319 ();
 FILLCELL_X1 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_338 ();
 FILLCELL_X32 FILLER_49_370 ();
 FILLCELL_X8 FILLER_49_402 ();
 FILLCELL_X4 FILLER_49_410 ();
 FILLCELL_X2 FILLER_49_414 ();
 FILLCELL_X1 FILLER_49_416 ();
 FILLCELL_X16 FILLER_49_424 ();
 FILLCELL_X2 FILLER_49_468 ();
 FILLCELL_X8 FILLER_49_472 ();
 FILLCELL_X32 FILLER_49_487 ();
 FILLCELL_X4 FILLER_49_519 ();
 FILLCELL_X1 FILLER_49_523 ();
 FILLCELL_X8 FILLER_49_531 ();
 FILLCELL_X4 FILLER_49_539 ();
 FILLCELL_X1 FILLER_49_543 ();
 FILLCELL_X4 FILLER_49_548 ();
 FILLCELL_X2 FILLER_49_552 ();
 FILLCELL_X2 FILLER_49_561 ();
 FILLCELL_X1 FILLER_49_580 ();
 FILLCELL_X1 FILLER_49_603 ();
 FILLCELL_X32 FILLER_49_607 ();
 FILLCELL_X32 FILLER_49_639 ();
 FILLCELL_X32 FILLER_49_671 ();
 FILLCELL_X32 FILLER_49_703 ();
 FILLCELL_X32 FILLER_49_735 ();
 FILLCELL_X32 FILLER_49_767 ();
 FILLCELL_X16 FILLER_49_799 ();
 FILLCELL_X8 FILLER_49_815 ();
 FILLCELL_X1 FILLER_49_823 ();
 FILLCELL_X32 FILLER_49_827 ();
 FILLCELL_X4 FILLER_49_859 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X4 FILLER_50_289 ();
 FILLCELL_X2 FILLER_50_293 ();
 FILLCELL_X16 FILLER_50_309 ();
 FILLCELL_X8 FILLER_50_325 ();
 FILLCELL_X4 FILLER_50_333 ();
 FILLCELL_X2 FILLER_50_337 ();
 FILLCELL_X1 FILLER_50_339 ();
 FILLCELL_X32 FILLER_50_347 ();
 FILLCELL_X2 FILLER_50_379 ();
 FILLCELL_X4 FILLER_50_388 ();
 FILLCELL_X2 FILLER_50_392 ();
 FILLCELL_X1 FILLER_50_394 ();
 FILLCELL_X4 FILLER_50_409 ();
 FILLCELL_X4 FILLER_50_420 ();
 FILLCELL_X1 FILLER_50_424 ();
 FILLCELL_X2 FILLER_50_443 ();
 FILLCELL_X1 FILLER_50_445 ();
 FILLCELL_X1 FILLER_50_457 ();
 FILLCELL_X1 FILLER_50_462 ();
 FILLCELL_X4 FILLER_50_467 ();
 FILLCELL_X1 FILLER_50_471 ();
 FILLCELL_X16 FILLER_50_486 ();
 FILLCELL_X8 FILLER_50_502 ();
 FILLCELL_X1 FILLER_50_510 ();
 FILLCELL_X1 FILLER_50_518 ();
 FILLCELL_X2 FILLER_50_523 ();
 FILLCELL_X2 FILLER_50_541 ();
 FILLCELL_X4 FILLER_50_561 ();
 FILLCELL_X1 FILLER_50_565 ();
 FILLCELL_X32 FILLER_50_591 ();
 FILLCELL_X8 FILLER_50_623 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X8 FILLER_50_824 ();
 FILLCELL_X2 FILLER_50_836 ();
 FILLCELL_X16 FILLER_50_841 ();
 FILLCELL_X4 FILLER_50_857 ();
 FILLCELL_X2 FILLER_50_861 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X8 FILLER_51_289 ();
 FILLCELL_X2 FILLER_51_297 ();
 FILLCELL_X8 FILLER_51_320 ();
 FILLCELL_X32 FILLER_51_342 ();
 FILLCELL_X2 FILLER_51_374 ();
 FILLCELL_X32 FILLER_51_383 ();
 FILLCELL_X4 FILLER_51_415 ();
 FILLCELL_X8 FILLER_51_422 ();
 FILLCELL_X1 FILLER_51_430 ();
 FILLCELL_X8 FILLER_51_438 ();
 FILLCELL_X4 FILLER_51_446 ();
 FILLCELL_X2 FILLER_51_450 ();
 FILLCELL_X1 FILLER_51_452 ();
 FILLCELL_X16 FILLER_51_456 ();
 FILLCELL_X2 FILLER_51_472 ();
 FILLCELL_X1 FILLER_51_474 ();
 FILLCELL_X2 FILLER_51_490 ();
 FILLCELL_X2 FILLER_51_495 ();
 FILLCELL_X1 FILLER_51_500 ();
 FILLCELL_X8 FILLER_51_518 ();
 FILLCELL_X1 FILLER_51_526 ();
 FILLCELL_X8 FILLER_51_552 ();
 FILLCELL_X4 FILLER_51_560 ();
 FILLCELL_X2 FILLER_51_564 ();
 FILLCELL_X32 FILLER_51_591 ();
 FILLCELL_X32 FILLER_51_623 ();
 FILLCELL_X32 FILLER_51_655 ();
 FILLCELL_X32 FILLER_51_687 ();
 FILLCELL_X32 FILLER_51_719 ();
 FILLCELL_X32 FILLER_51_751 ();
 FILLCELL_X32 FILLER_51_783 ();
 FILLCELL_X32 FILLER_51_815 ();
 FILLCELL_X8 FILLER_51_847 ();
 FILLCELL_X2 FILLER_51_855 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X8 FILLER_52_289 ();
 FILLCELL_X4 FILLER_52_306 ();
 FILLCELL_X8 FILLER_52_338 ();
 FILLCELL_X4 FILLER_52_346 ();
 FILLCELL_X2 FILLER_52_350 ();
 FILLCELL_X1 FILLER_52_352 ();
 FILLCELL_X4 FILLER_52_360 ();
 FILLCELL_X2 FILLER_52_364 ();
 FILLCELL_X1 FILLER_52_366 ();
 FILLCELL_X2 FILLER_52_374 ();
 FILLCELL_X4 FILLER_52_383 ();
 FILLCELL_X32 FILLER_52_394 ();
 FILLCELL_X8 FILLER_52_426 ();
 FILLCELL_X4 FILLER_52_434 ();
 FILLCELL_X1 FILLER_52_438 ();
 FILLCELL_X8 FILLER_52_441 ();
 FILLCELL_X4 FILLER_52_449 ();
 FILLCELL_X4 FILLER_52_460 ();
 FILLCELL_X2 FILLER_52_464 ();
 FILLCELL_X2 FILLER_52_473 ();
 FILLCELL_X1 FILLER_52_475 ();
 FILLCELL_X16 FILLER_52_482 ();
 FILLCELL_X2 FILLER_52_498 ();
 FILLCELL_X1 FILLER_52_500 ();
 FILLCELL_X4 FILLER_52_512 ();
 FILLCELL_X2 FILLER_52_516 ();
 FILLCELL_X2 FILLER_52_529 ();
 FILLCELL_X1 FILLER_52_531 ();
 FILLCELL_X2 FILLER_52_557 ();
 FILLCELL_X1 FILLER_52_559 ();
 FILLCELL_X1 FILLER_52_567 ();
 FILLCELL_X32 FILLER_52_588 ();
 FILLCELL_X8 FILLER_52_620 ();
 FILLCELL_X2 FILLER_52_628 ();
 FILLCELL_X1 FILLER_52_630 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X32 FILLER_52_760 ();
 FILLCELL_X16 FILLER_52_792 ();
 FILLCELL_X8 FILLER_52_808 ();
 FILLCELL_X4 FILLER_52_816 ();
 FILLCELL_X2 FILLER_52_820 ();
 FILLCELL_X16 FILLER_52_825 ();
 FILLCELL_X4 FILLER_52_841 ();
 FILLCELL_X8 FILLER_52_848 ();
 FILLCELL_X4 FILLER_52_856 ();
 FILLCELL_X2 FILLER_52_860 ();
 FILLCELL_X1 FILLER_52_862 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X8 FILLER_53_289 ();
 FILLCELL_X1 FILLER_53_311 ();
 FILLCELL_X4 FILLER_53_319 ();
 FILLCELL_X1 FILLER_53_323 ();
 FILLCELL_X4 FILLER_53_333 ();
 FILLCELL_X32 FILLER_53_346 ();
 FILLCELL_X8 FILLER_53_378 ();
 FILLCELL_X4 FILLER_53_393 ();
 FILLCELL_X2 FILLER_53_397 ();
 FILLCELL_X1 FILLER_53_399 ();
 FILLCELL_X1 FILLER_53_407 ();
 FILLCELL_X4 FILLER_53_420 ();
 FILLCELL_X2 FILLER_53_424 ();
 FILLCELL_X1 FILLER_53_426 ();
 FILLCELL_X1 FILLER_53_434 ();
 FILLCELL_X4 FILLER_53_452 ();
 FILLCELL_X2 FILLER_53_456 ();
 FILLCELL_X8 FILLER_53_462 ();
 FILLCELL_X2 FILLER_53_470 ();
 FILLCELL_X1 FILLER_53_472 ();
 FILLCELL_X8 FILLER_53_482 ();
 FILLCELL_X2 FILLER_53_490 ();
 FILLCELL_X1 FILLER_53_492 ();
 FILLCELL_X8 FILLER_53_510 ();
 FILLCELL_X4 FILLER_53_529 ();
 FILLCELL_X1 FILLER_53_533 ();
 FILLCELL_X16 FILLER_53_541 ();
 FILLCELL_X8 FILLER_53_557 ();
 FILLCELL_X2 FILLER_53_565 ();
 FILLCELL_X32 FILLER_53_584 ();
 FILLCELL_X32 FILLER_53_616 ();
 FILLCELL_X32 FILLER_53_648 ();
 FILLCELL_X32 FILLER_53_680 ();
 FILLCELL_X32 FILLER_53_712 ();
 FILLCELL_X32 FILLER_53_744 ();
 FILLCELL_X32 FILLER_53_776 ();
 FILLCELL_X16 FILLER_53_808 ();
 FILLCELL_X8 FILLER_53_827 ();
 FILLCELL_X2 FILLER_53_835 ();
 FILLCELL_X8 FILLER_53_840 ();
 FILLCELL_X8 FILLER_53_851 ();
 FILLCELL_X4 FILLER_53_859 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X16 FILLER_54_257 ();
 FILLCELL_X8 FILLER_54_273 ();
 FILLCELL_X2 FILLER_54_281 ();
 FILLCELL_X2 FILLER_54_332 ();
 FILLCELL_X1 FILLER_54_334 ();
 FILLCELL_X4 FILLER_54_349 ();
 FILLCELL_X2 FILLER_54_353 ();
 FILLCELL_X1 FILLER_54_355 ();
 FILLCELL_X16 FILLER_54_363 ();
 FILLCELL_X8 FILLER_54_379 ();
 FILLCELL_X2 FILLER_54_394 ();
 FILLCELL_X1 FILLER_54_396 ();
 FILLCELL_X2 FILLER_54_404 ();
 FILLCELL_X2 FILLER_54_417 ();
 FILLCELL_X2 FILLER_54_456 ();
 FILLCELL_X8 FILLER_54_472 ();
 FILLCELL_X2 FILLER_54_480 ();
 FILLCELL_X1 FILLER_54_482 ();
 FILLCELL_X2 FILLER_54_519 ();
 FILLCELL_X8 FILLER_54_536 ();
 FILLCELL_X2 FILLER_54_544 ();
 FILLCELL_X1 FILLER_54_546 ();
 FILLCELL_X4 FILLER_54_554 ();
 FILLCELL_X2 FILLER_54_558 ();
 FILLCELL_X1 FILLER_54_560 ();
 FILLCELL_X4 FILLER_54_568 ();
 FILLCELL_X2 FILLER_54_572 ();
 FILLCELL_X4 FILLER_54_578 ();
 FILLCELL_X1 FILLER_54_582 ();
 FILLCELL_X32 FILLER_54_594 ();
 FILLCELL_X4 FILLER_54_626 ();
 FILLCELL_X1 FILLER_54_630 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X32 FILLER_54_728 ();
 FILLCELL_X32 FILLER_54_760 ();
 FILLCELL_X32 FILLER_54_792 ();
 FILLCELL_X16 FILLER_54_824 ();
 FILLCELL_X8 FILLER_54_840 ();
 FILLCELL_X4 FILLER_54_848 ();
 FILLCELL_X4 FILLER_54_856 ();
 FILLCELL_X2 FILLER_54_860 ();
 FILLCELL_X1 FILLER_54_862 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X16 FILLER_55_289 ();
 FILLCELL_X4 FILLER_55_305 ();
 FILLCELL_X2 FILLER_55_309 ();
 FILLCELL_X1 FILLER_55_311 ();
 FILLCELL_X2 FILLER_55_319 ();
 FILLCELL_X1 FILLER_55_321 ();
 FILLCELL_X2 FILLER_55_329 ();
 FILLCELL_X1 FILLER_55_331 ();
 FILLCELL_X16 FILLER_55_339 ();
 FILLCELL_X4 FILLER_55_355 ();
 FILLCELL_X2 FILLER_55_359 ();
 FILLCELL_X8 FILLER_55_368 ();
 FILLCELL_X2 FILLER_55_376 ();
 FILLCELL_X1 FILLER_55_378 ();
 FILLCELL_X16 FILLER_55_386 ();
 FILLCELL_X4 FILLER_55_402 ();
 FILLCELL_X1 FILLER_55_406 ();
 FILLCELL_X1 FILLER_55_414 ();
 FILLCELL_X8 FILLER_55_422 ();
 FILLCELL_X1 FILLER_55_430 ();
 FILLCELL_X16 FILLER_55_451 ();
 FILLCELL_X1 FILLER_55_467 ();
 FILLCELL_X2 FILLER_55_472 ();
 FILLCELL_X4 FILLER_55_480 ();
 FILLCELL_X4 FILLER_55_491 ();
 FILLCELL_X1 FILLER_55_495 ();
 FILLCELL_X16 FILLER_55_500 ();
 FILLCELL_X4 FILLER_55_516 ();
 FILLCELL_X1 FILLER_55_520 ();
 FILLCELL_X2 FILLER_55_544 ();
 FILLCELL_X1 FILLER_55_546 ();
 FILLCELL_X4 FILLER_55_556 ();
 FILLCELL_X8 FILLER_55_576 ();
 FILLCELL_X32 FILLER_55_587 ();
 FILLCELL_X32 FILLER_55_619 ();
 FILLCELL_X32 FILLER_55_651 ();
 FILLCELL_X32 FILLER_55_683 ();
 FILLCELL_X32 FILLER_55_715 ();
 FILLCELL_X32 FILLER_55_747 ();
 FILLCELL_X32 FILLER_55_779 ();
 FILLCELL_X8 FILLER_55_811 ();
 FILLCELL_X4 FILLER_55_819 ();
 FILLCELL_X32 FILLER_55_826 ();
 FILLCELL_X4 FILLER_55_858 ();
 FILLCELL_X1 FILLER_55_862 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X8 FILLER_56_289 ();
 FILLCELL_X1 FILLER_56_297 ();
 FILLCELL_X4 FILLER_56_305 ();
 FILLCELL_X2 FILLER_56_309 ();
 FILLCELL_X1 FILLER_56_311 ();
 FILLCELL_X4 FILLER_56_319 ();
 FILLCELL_X1 FILLER_56_323 ();
 FILLCELL_X16 FILLER_56_338 ();
 FILLCELL_X4 FILLER_56_354 ();
 FILLCELL_X2 FILLER_56_358 ();
 FILLCELL_X1 FILLER_56_360 ();
 FILLCELL_X32 FILLER_56_368 ();
 FILLCELL_X16 FILLER_56_400 ();
 FILLCELL_X4 FILLER_56_416 ();
 FILLCELL_X16 FILLER_56_431 ();
 FILLCELL_X8 FILLER_56_447 ();
 FILLCELL_X4 FILLER_56_455 ();
 FILLCELL_X2 FILLER_56_459 ();
 FILLCELL_X8 FILLER_56_464 ();
 FILLCELL_X4 FILLER_56_472 ();
 FILLCELL_X1 FILLER_56_476 ();
 FILLCELL_X2 FILLER_56_482 ();
 FILLCELL_X2 FILLER_56_488 ();
 FILLCELL_X2 FILLER_56_497 ();
 FILLCELL_X1 FILLER_56_499 ();
 FILLCELL_X16 FILLER_56_507 ();
 FILLCELL_X2 FILLER_56_523 ();
 FILLCELL_X1 FILLER_56_525 ();
 FILLCELL_X2 FILLER_56_539 ();
 FILLCELL_X8 FILLER_56_558 ();
 FILLCELL_X4 FILLER_56_566 ();
 FILLCELL_X2 FILLER_56_570 ();
 FILLCELL_X1 FILLER_56_572 ();
 FILLCELL_X2 FILLER_56_592 ();
 FILLCELL_X1 FILLER_56_594 ();
 FILLCELL_X16 FILLER_56_602 ();
 FILLCELL_X8 FILLER_56_618 ();
 FILLCELL_X4 FILLER_56_626 ();
 FILLCELL_X1 FILLER_56_630 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X32 FILLER_56_760 ();
 FILLCELL_X32 FILLER_56_792 ();
 FILLCELL_X4 FILLER_56_824 ();
 FILLCELL_X1 FILLER_56_828 ();
 FILLCELL_X1 FILLER_56_832 ();
 FILLCELL_X8 FILLER_56_836 ();
 FILLCELL_X2 FILLER_56_847 ();
 FILLCELL_X1 FILLER_56_849 ();
 FILLCELL_X8 FILLER_56_853 ();
 FILLCELL_X2 FILLER_56_861 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X16 FILLER_57_289 ();
 FILLCELL_X4 FILLER_57_305 ();
 FILLCELL_X2 FILLER_57_309 ();
 FILLCELL_X1 FILLER_57_311 ();
 FILLCELL_X4 FILLER_57_326 ();
 FILLCELL_X2 FILLER_57_330 ();
 FILLCELL_X16 FILLER_57_346 ();
 FILLCELL_X1 FILLER_57_362 ();
 FILLCELL_X32 FILLER_57_370 ();
 FILLCELL_X8 FILLER_57_402 ();
 FILLCELL_X2 FILLER_57_410 ();
 FILLCELL_X1 FILLER_57_443 ();
 FILLCELL_X2 FILLER_57_458 ();
 FILLCELL_X1 FILLER_57_460 ();
 FILLCELL_X8 FILLER_57_479 ();
 FILLCELL_X8 FILLER_57_496 ();
 FILLCELL_X4 FILLER_57_504 ();
 FILLCELL_X2 FILLER_57_508 ();
 FILLCELL_X1 FILLER_57_510 ();
 FILLCELL_X4 FILLER_57_530 ();
 FILLCELL_X2 FILLER_57_534 ();
 FILLCELL_X2 FILLER_57_543 ();
 FILLCELL_X16 FILLER_57_548 ();
 FILLCELL_X2 FILLER_57_564 ();
 FILLCELL_X1 FILLER_57_566 ();
 FILLCELL_X4 FILLER_57_570 ();
 FILLCELL_X2 FILLER_57_574 ();
 FILLCELL_X1 FILLER_57_576 ();
 FILLCELL_X1 FILLER_57_581 ();
 FILLCELL_X32 FILLER_57_593 ();
 FILLCELL_X32 FILLER_57_625 ();
 FILLCELL_X32 FILLER_57_657 ();
 FILLCELL_X32 FILLER_57_689 ();
 FILLCELL_X32 FILLER_57_721 ();
 FILLCELL_X32 FILLER_57_753 ();
 FILLCELL_X32 FILLER_57_785 ();
 FILLCELL_X4 FILLER_57_817 ();
 FILLCELL_X2 FILLER_57_821 ();
 FILLCELL_X1 FILLER_57_823 ();
 FILLCELL_X32 FILLER_57_828 ();
 FILLCELL_X2 FILLER_57_860 ();
 FILLCELL_X1 FILLER_57_862 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X8 FILLER_58_257 ();
 FILLCELL_X4 FILLER_58_265 ();
 FILLCELL_X1 FILLER_58_269 ();
 FILLCELL_X8 FILLER_58_303 ();
 FILLCELL_X4 FILLER_58_311 ();
 FILLCELL_X2 FILLER_58_315 ();
 FILLCELL_X32 FILLER_58_320 ();
 FILLCELL_X32 FILLER_58_352 ();
 FILLCELL_X16 FILLER_58_384 ();
 FILLCELL_X2 FILLER_58_400 ();
 FILLCELL_X1 FILLER_58_402 ();
 FILLCELL_X16 FILLER_58_410 ();
 FILLCELL_X4 FILLER_58_426 ();
 FILLCELL_X2 FILLER_58_430 ();
 FILLCELL_X1 FILLER_58_443 ();
 FILLCELL_X2 FILLER_58_447 ();
 FILLCELL_X1 FILLER_58_449 ();
 FILLCELL_X4 FILLER_58_466 ();
 FILLCELL_X1 FILLER_58_474 ();
 FILLCELL_X2 FILLER_58_489 ();
 FILLCELL_X4 FILLER_58_494 ();
 FILLCELL_X2 FILLER_58_507 ();
 FILLCELL_X1 FILLER_58_516 ();
 FILLCELL_X1 FILLER_58_534 ();
 FILLCELL_X1 FILLER_58_572 ();
 FILLCELL_X16 FILLER_58_580 ();
 FILLCELL_X16 FILLER_58_601 ();
 FILLCELL_X8 FILLER_58_617 ();
 FILLCELL_X4 FILLER_58_625 ();
 FILLCELL_X2 FILLER_58_629 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X4 FILLER_58_856 ();
 FILLCELL_X2 FILLER_58_860 ();
 FILLCELL_X1 FILLER_58_862 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X4 FILLER_59_321 ();
 FILLCELL_X1 FILLER_59_325 ();
 FILLCELL_X8 FILLER_59_333 ();
 FILLCELL_X4 FILLER_59_341 ();
 FILLCELL_X2 FILLER_59_345 ();
 FILLCELL_X32 FILLER_59_368 ();
 FILLCELL_X4 FILLER_59_400 ();
 FILLCELL_X16 FILLER_59_409 ();
 FILLCELL_X1 FILLER_59_425 ();
 FILLCELL_X8 FILLER_59_437 ();
 FILLCELL_X4 FILLER_59_445 ();
 FILLCELL_X2 FILLER_59_449 ();
 FILLCELL_X16 FILLER_59_472 ();
 FILLCELL_X4 FILLER_59_488 ();
 FILLCELL_X1 FILLER_59_492 ();
 FILLCELL_X4 FILLER_59_500 ();
 FILLCELL_X1 FILLER_59_523 ();
 FILLCELL_X4 FILLER_59_531 ();
 FILLCELL_X1 FILLER_59_535 ();
 FILLCELL_X32 FILLER_59_552 ();
 FILLCELL_X32 FILLER_59_584 ();
 FILLCELL_X32 FILLER_59_616 ();
 FILLCELL_X32 FILLER_59_648 ();
 FILLCELL_X32 FILLER_59_680 ();
 FILLCELL_X32 FILLER_59_712 ();
 FILLCELL_X32 FILLER_59_744 ();
 FILLCELL_X32 FILLER_59_776 ();
 FILLCELL_X32 FILLER_59_808 ();
 FILLCELL_X16 FILLER_59_840 ();
 FILLCELL_X4 FILLER_59_856 ();
 FILLCELL_X2 FILLER_59_860 ();
 FILLCELL_X1 FILLER_59_862 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X4 FILLER_60_321 ();
 FILLCELL_X16 FILLER_60_332 ();
 FILLCELL_X1 FILLER_60_369 ();
 FILLCELL_X8 FILLER_60_377 ();
 FILLCELL_X4 FILLER_60_385 ();
 FILLCELL_X2 FILLER_60_389 ();
 FILLCELL_X1 FILLER_60_391 ();
 FILLCELL_X16 FILLER_60_399 ();
 FILLCELL_X2 FILLER_60_415 ();
 FILLCELL_X1 FILLER_60_417 ();
 FILLCELL_X2 FILLER_60_425 ();
 FILLCELL_X4 FILLER_60_448 ();
 FILLCELL_X2 FILLER_60_470 ();
 FILLCELL_X2 FILLER_60_479 ();
 FILLCELL_X8 FILLER_60_490 ();
 FILLCELL_X2 FILLER_60_498 ();
 FILLCELL_X1 FILLER_60_500 ();
 FILLCELL_X2 FILLER_60_519 ();
 FILLCELL_X32 FILLER_60_532 ();
 FILLCELL_X32 FILLER_60_564 ();
 FILLCELL_X32 FILLER_60_596 ();
 FILLCELL_X2 FILLER_60_628 ();
 FILLCELL_X1 FILLER_60_630 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X32 FILLER_60_760 ();
 FILLCELL_X32 FILLER_60_792 ();
 FILLCELL_X32 FILLER_60_824 ();
 FILLCELL_X4 FILLER_60_856 ();
 FILLCELL_X2 FILLER_60_860 ();
 FILLCELL_X1 FILLER_60_862 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X16 FILLER_61_353 ();
 FILLCELL_X8 FILLER_61_369 ();
 FILLCELL_X1 FILLER_61_377 ();
 FILLCELL_X16 FILLER_61_385 ();
 FILLCELL_X2 FILLER_61_401 ();
 FILLCELL_X2 FILLER_61_417 ();
 FILLCELL_X8 FILLER_61_440 ();
 FILLCELL_X2 FILLER_61_455 ();
 FILLCELL_X4 FILLER_61_469 ();
 FILLCELL_X4 FILLER_61_478 ();
 FILLCELL_X2 FILLER_61_489 ();
 FILLCELL_X1 FILLER_61_491 ();
 FILLCELL_X2 FILLER_61_499 ();
 FILLCELL_X8 FILLER_61_506 ();
 FILLCELL_X2 FILLER_61_514 ();
 FILLCELL_X2 FILLER_61_521 ();
 FILLCELL_X32 FILLER_61_530 ();
 FILLCELL_X32 FILLER_61_562 ();
 FILLCELL_X32 FILLER_61_594 ();
 FILLCELL_X32 FILLER_61_626 ();
 FILLCELL_X32 FILLER_61_658 ();
 FILLCELL_X32 FILLER_61_690 ();
 FILLCELL_X32 FILLER_61_722 ();
 FILLCELL_X32 FILLER_61_754 ();
 FILLCELL_X32 FILLER_61_786 ();
 FILLCELL_X32 FILLER_61_818 ();
 FILLCELL_X8 FILLER_61_850 ();
 FILLCELL_X4 FILLER_61_858 ();
 FILLCELL_X1 FILLER_61_862 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X32 FILLER_62_129 ();
 FILLCELL_X32 FILLER_62_161 ();
 FILLCELL_X32 FILLER_62_193 ();
 FILLCELL_X32 FILLER_62_225 ();
 FILLCELL_X32 FILLER_62_257 ();
 FILLCELL_X32 FILLER_62_289 ();
 FILLCELL_X32 FILLER_62_321 ();
 FILLCELL_X32 FILLER_62_353 ();
 FILLCELL_X16 FILLER_62_385 ();
 FILLCELL_X8 FILLER_62_401 ();
 FILLCELL_X4 FILLER_62_409 ();
 FILLCELL_X1 FILLER_62_413 ();
 FILLCELL_X8 FILLER_62_432 ();
 FILLCELL_X4 FILLER_62_440 ();
 FILLCELL_X2 FILLER_62_444 ();
 FILLCELL_X1 FILLER_62_446 ();
 FILLCELL_X8 FILLER_62_461 ();
 FILLCELL_X4 FILLER_62_469 ();
 FILLCELL_X4 FILLER_62_478 ();
 FILLCELL_X2 FILLER_62_482 ();
 FILLCELL_X4 FILLER_62_505 ();
 FILLCELL_X1 FILLER_62_509 ();
 FILLCELL_X32 FILLER_62_513 ();
 FILLCELL_X32 FILLER_62_545 ();
 FILLCELL_X32 FILLER_62_577 ();
 FILLCELL_X16 FILLER_62_609 ();
 FILLCELL_X4 FILLER_62_625 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X4 FILLER_62_856 ();
 FILLCELL_X2 FILLER_62_860 ();
 FILLCELL_X1 FILLER_62_862 ();
 FILLCELL_X16 FILLER_63_1 ();
 FILLCELL_X4 FILLER_63_17 ();
 FILLCELL_X1 FILLER_63_21 ();
 FILLCELL_X32 FILLER_63_27 ();
 FILLCELL_X32 FILLER_63_59 ();
 FILLCELL_X32 FILLER_63_91 ();
 FILLCELL_X32 FILLER_63_123 ();
 FILLCELL_X32 FILLER_63_155 ();
 FILLCELL_X32 FILLER_63_187 ();
 FILLCELL_X32 FILLER_63_219 ();
 FILLCELL_X32 FILLER_63_251 ();
 FILLCELL_X32 FILLER_63_283 ();
 FILLCELL_X32 FILLER_63_315 ();
 FILLCELL_X16 FILLER_63_347 ();
 FILLCELL_X8 FILLER_63_363 ();
 FILLCELL_X4 FILLER_63_371 ();
 FILLCELL_X1 FILLER_63_375 ();
 FILLCELL_X2 FILLER_63_385 ();
 FILLCELL_X1 FILLER_63_387 ();
 FILLCELL_X16 FILLER_63_411 ();
 FILLCELL_X8 FILLER_63_427 ();
 FILLCELL_X4 FILLER_63_435 ();
 FILLCELL_X8 FILLER_63_449 ();
 FILLCELL_X2 FILLER_63_457 ();
 FILLCELL_X4 FILLER_63_464 ();
 FILLCELL_X1 FILLER_63_468 ();
 FILLCELL_X4 FILLER_63_494 ();
 FILLCELL_X2 FILLER_63_511 ();
 FILLCELL_X1 FILLER_63_513 ();
 FILLCELL_X8 FILLER_63_523 ();
 FILLCELL_X4 FILLER_63_540 ();
 FILLCELL_X1 FILLER_63_544 ();
 FILLCELL_X32 FILLER_63_550 ();
 FILLCELL_X32 FILLER_63_582 ();
 FILLCELL_X32 FILLER_63_614 ();
 FILLCELL_X32 FILLER_63_646 ();
 FILLCELL_X32 FILLER_63_678 ();
 FILLCELL_X32 FILLER_63_710 ();
 FILLCELL_X32 FILLER_63_742 ();
 FILLCELL_X32 FILLER_63_774 ();
 FILLCELL_X32 FILLER_63_806 ();
 FILLCELL_X16 FILLER_63_838 ();
 FILLCELL_X8 FILLER_63_854 ();
 FILLCELL_X1 FILLER_63_862 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X8 FILLER_64_385 ();
 FILLCELL_X2 FILLER_64_393 ();
 FILLCELL_X8 FILLER_64_415 ();
 FILLCELL_X4 FILLER_64_423 ();
 FILLCELL_X2 FILLER_64_427 ();
 FILLCELL_X1 FILLER_64_441 ();
 FILLCELL_X4 FILLER_64_448 ();
 FILLCELL_X2 FILLER_64_457 ();
 FILLCELL_X1 FILLER_64_463 ();
 FILLCELL_X1 FILLER_64_480 ();
 FILLCELL_X8 FILLER_64_508 ();
 FILLCELL_X4 FILLER_64_516 ();
 FILLCELL_X32 FILLER_64_527 ();
 FILLCELL_X32 FILLER_64_559 ();
 FILLCELL_X32 FILLER_64_591 ();
 FILLCELL_X8 FILLER_64_623 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X32 FILLER_64_760 ();
 FILLCELL_X32 FILLER_64_792 ();
 FILLCELL_X32 FILLER_64_824 ();
 FILLCELL_X4 FILLER_64_856 ();
 FILLCELL_X2 FILLER_64_860 ();
 FILLCELL_X1 FILLER_64_862 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X8 FILLER_65_417 ();
 FILLCELL_X1 FILLER_65_425 ();
 FILLCELL_X1 FILLER_65_429 ();
 FILLCELL_X1 FILLER_65_437 ();
 FILLCELL_X1 FILLER_65_455 ();
 FILLCELL_X2 FILLER_65_463 ();
 FILLCELL_X4 FILLER_65_472 ();
 FILLCELL_X4 FILLER_65_486 ();
 FILLCELL_X1 FILLER_65_490 ();
 FILLCELL_X4 FILLER_65_504 ();
 FILLCELL_X32 FILLER_65_515 ();
 FILLCELL_X1 FILLER_65_547 ();
 FILLCELL_X32 FILLER_65_553 ();
 FILLCELL_X32 FILLER_65_585 ();
 FILLCELL_X32 FILLER_65_617 ();
 FILLCELL_X32 FILLER_65_649 ();
 FILLCELL_X32 FILLER_65_681 ();
 FILLCELL_X32 FILLER_65_713 ();
 FILLCELL_X32 FILLER_65_745 ();
 FILLCELL_X32 FILLER_65_777 ();
 FILLCELL_X32 FILLER_65_809 ();
 FILLCELL_X16 FILLER_65_841 ();
 FILLCELL_X4 FILLER_65_857 ();
 FILLCELL_X2 FILLER_65_861 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X32 FILLER_66_353 ();
 FILLCELL_X32 FILLER_66_385 ();
 FILLCELL_X8 FILLER_66_417 ();
 FILLCELL_X4 FILLER_66_425 ();
 FILLCELL_X2 FILLER_66_429 ();
 FILLCELL_X1 FILLER_66_431 ();
 FILLCELL_X2 FILLER_66_449 ();
 FILLCELL_X1 FILLER_66_451 ();
 FILLCELL_X2 FILLER_66_455 ();
 FILLCELL_X1 FILLER_66_457 ();
 FILLCELL_X2 FILLER_66_461 ();
 FILLCELL_X1 FILLER_66_463 ();
 FILLCELL_X2 FILLER_66_487 ();
 FILLCELL_X2 FILLER_66_496 ();
 FILLCELL_X1 FILLER_66_498 ();
 FILLCELL_X32 FILLER_66_503 ();
 FILLCELL_X32 FILLER_66_535 ();
 FILLCELL_X32 FILLER_66_567 ();
 FILLCELL_X32 FILLER_66_599 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X32 FILLER_66_760 ();
 FILLCELL_X32 FILLER_66_792 ();
 FILLCELL_X32 FILLER_66_824 ();
 FILLCELL_X4 FILLER_66_856 ();
 FILLCELL_X2 FILLER_66_860 ();
 FILLCELL_X1 FILLER_66_862 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X16 FILLER_67_417 ();
 FILLCELL_X4 FILLER_67_433 ();
 FILLCELL_X2 FILLER_67_437 ();
 FILLCELL_X1 FILLER_67_439 ();
 FILLCELL_X32 FILLER_67_454 ();
 FILLCELL_X4 FILLER_67_486 ();
 FILLCELL_X1 FILLER_67_490 ();
 FILLCELL_X32 FILLER_67_498 ();
 FILLCELL_X16 FILLER_67_530 ();
 FILLCELL_X32 FILLER_67_560 ();
 FILLCELL_X32 FILLER_67_592 ();
 FILLCELL_X32 FILLER_67_624 ();
 FILLCELL_X32 FILLER_67_656 ();
 FILLCELL_X32 FILLER_67_688 ();
 FILLCELL_X32 FILLER_67_720 ();
 FILLCELL_X32 FILLER_67_752 ();
 FILLCELL_X32 FILLER_67_784 ();
 FILLCELL_X32 FILLER_67_816 ();
 FILLCELL_X8 FILLER_67_848 ();
 FILLCELL_X4 FILLER_67_856 ();
 FILLCELL_X2 FILLER_67_860 ();
 FILLCELL_X1 FILLER_67_862 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X2 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_308 ();
 FILLCELL_X32 FILLER_68_340 ();
 FILLCELL_X32 FILLER_68_372 ();
 FILLCELL_X32 FILLER_68_404 ();
 FILLCELL_X4 FILLER_68_436 ();
 FILLCELL_X2 FILLER_68_440 ();
 FILLCELL_X1 FILLER_68_442 ();
 FILLCELL_X32 FILLER_68_450 ();
 FILLCELL_X32 FILLER_68_482 ();
 FILLCELL_X32 FILLER_68_514 ();
 FILLCELL_X32 FILLER_68_546 ();
 FILLCELL_X32 FILLER_68_578 ();
 FILLCELL_X16 FILLER_68_610 ();
 FILLCELL_X4 FILLER_68_626 ();
 FILLCELL_X1 FILLER_68_630 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X32 FILLER_68_760 ();
 FILLCELL_X32 FILLER_68_792 ();
 FILLCELL_X32 FILLER_68_824 ();
 FILLCELL_X4 FILLER_68_856 ();
 FILLCELL_X2 FILLER_68_860 ();
 FILLCELL_X1 FILLER_68_862 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X32 FILLER_69_449 ();
 FILLCELL_X32 FILLER_69_481 ();
 FILLCELL_X32 FILLER_69_513 ();
 FILLCELL_X32 FILLER_69_545 ();
 FILLCELL_X32 FILLER_69_577 ();
 FILLCELL_X32 FILLER_69_609 ();
 FILLCELL_X32 FILLER_69_641 ();
 FILLCELL_X32 FILLER_69_673 ();
 FILLCELL_X32 FILLER_69_705 ();
 FILLCELL_X32 FILLER_69_737 ();
 FILLCELL_X32 FILLER_69_769 ();
 FILLCELL_X32 FILLER_69_801 ();
 FILLCELL_X16 FILLER_69_833 ();
 FILLCELL_X8 FILLER_69_849 ();
 FILLCELL_X4 FILLER_69_857 ();
 FILLCELL_X2 FILLER_69_861 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X16 FILLER_70_353 ();
 FILLCELL_X4 FILLER_70_369 ();
 FILLCELL_X32 FILLER_70_380 ();
 FILLCELL_X32 FILLER_70_412 ();
 FILLCELL_X32 FILLER_70_444 ();
 FILLCELL_X32 FILLER_70_476 ();
 FILLCELL_X32 FILLER_70_508 ();
 FILLCELL_X32 FILLER_70_540 ();
 FILLCELL_X32 FILLER_70_572 ();
 FILLCELL_X16 FILLER_70_604 ();
 FILLCELL_X8 FILLER_70_620 ();
 FILLCELL_X2 FILLER_70_628 ();
 FILLCELL_X1 FILLER_70_630 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X32 FILLER_70_760 ();
 FILLCELL_X32 FILLER_70_792 ();
 FILLCELL_X32 FILLER_70_824 ();
 FILLCELL_X4 FILLER_70_856 ();
 FILLCELL_X2 FILLER_70_860 ();
 FILLCELL_X1 FILLER_70_862 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X32 FILLER_71_449 ();
 FILLCELL_X32 FILLER_71_481 ();
 FILLCELL_X32 FILLER_71_513 ();
 FILLCELL_X32 FILLER_71_545 ();
 FILLCELL_X32 FILLER_71_577 ();
 FILLCELL_X32 FILLER_71_609 ();
 FILLCELL_X32 FILLER_71_641 ();
 FILLCELL_X32 FILLER_71_673 ();
 FILLCELL_X32 FILLER_71_705 ();
 FILLCELL_X32 FILLER_71_737 ();
 FILLCELL_X32 FILLER_71_769 ();
 FILLCELL_X32 FILLER_71_801 ();
 FILLCELL_X16 FILLER_71_833 ();
 FILLCELL_X8 FILLER_71_849 ();
 FILLCELL_X4 FILLER_71_857 ();
 FILLCELL_X2 FILLER_71_861 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X32 FILLER_72_353 ();
 FILLCELL_X32 FILLER_72_385 ();
 FILLCELL_X32 FILLER_72_417 ();
 FILLCELL_X32 FILLER_72_449 ();
 FILLCELL_X32 FILLER_72_481 ();
 FILLCELL_X32 FILLER_72_513 ();
 FILLCELL_X32 FILLER_72_545 ();
 FILLCELL_X32 FILLER_72_577 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X32 FILLER_72_760 ();
 FILLCELL_X32 FILLER_72_792 ();
 FILLCELL_X32 FILLER_72_824 ();
 FILLCELL_X4 FILLER_72_856 ();
 FILLCELL_X2 FILLER_72_860 ();
 FILLCELL_X1 FILLER_72_862 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X32 FILLER_73_385 ();
 FILLCELL_X32 FILLER_73_417 ();
 FILLCELL_X32 FILLER_73_449 ();
 FILLCELL_X32 FILLER_73_481 ();
 FILLCELL_X32 FILLER_73_513 ();
 FILLCELL_X32 FILLER_73_545 ();
 FILLCELL_X32 FILLER_73_577 ();
 FILLCELL_X32 FILLER_73_609 ();
 FILLCELL_X32 FILLER_73_641 ();
 FILLCELL_X32 FILLER_73_673 ();
 FILLCELL_X32 FILLER_73_705 ();
 FILLCELL_X32 FILLER_73_737 ();
 FILLCELL_X32 FILLER_73_769 ();
 FILLCELL_X32 FILLER_73_801 ();
 FILLCELL_X16 FILLER_73_833 ();
 FILLCELL_X8 FILLER_73_849 ();
 FILLCELL_X4 FILLER_73_857 ();
 FILLCELL_X2 FILLER_73_861 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X32 FILLER_74_353 ();
 FILLCELL_X32 FILLER_74_385 ();
 FILLCELL_X32 FILLER_74_417 ();
 FILLCELL_X32 FILLER_74_449 ();
 FILLCELL_X32 FILLER_74_481 ();
 FILLCELL_X32 FILLER_74_513 ();
 FILLCELL_X32 FILLER_74_545 ();
 FILLCELL_X32 FILLER_74_577 ();
 FILLCELL_X16 FILLER_74_609 ();
 FILLCELL_X4 FILLER_74_625 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X32 FILLER_74_760 ();
 FILLCELL_X32 FILLER_74_792 ();
 FILLCELL_X32 FILLER_74_824 ();
 FILLCELL_X4 FILLER_74_856 ();
 FILLCELL_X2 FILLER_74_860 ();
 FILLCELL_X1 FILLER_74_862 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X32 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_513 ();
 FILLCELL_X32 FILLER_75_545 ();
 FILLCELL_X32 FILLER_75_577 ();
 FILLCELL_X32 FILLER_75_609 ();
 FILLCELL_X32 FILLER_75_641 ();
 FILLCELL_X32 FILLER_75_673 ();
 FILLCELL_X32 FILLER_75_705 ();
 FILLCELL_X32 FILLER_75_737 ();
 FILLCELL_X32 FILLER_75_769 ();
 FILLCELL_X32 FILLER_75_801 ();
 FILLCELL_X16 FILLER_75_833 ();
 FILLCELL_X8 FILLER_75_849 ();
 FILLCELL_X4 FILLER_75_857 ();
 FILLCELL_X2 FILLER_75_861 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X32 FILLER_76_449 ();
 FILLCELL_X32 FILLER_76_481 ();
 FILLCELL_X32 FILLER_76_513 ();
 FILLCELL_X32 FILLER_76_545 ();
 FILLCELL_X32 FILLER_76_577 ();
 FILLCELL_X16 FILLER_76_609 ();
 FILLCELL_X4 FILLER_76_625 ();
 FILLCELL_X2 FILLER_76_629 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X32 FILLER_76_760 ();
 FILLCELL_X32 FILLER_76_792 ();
 FILLCELL_X32 FILLER_76_824 ();
 FILLCELL_X4 FILLER_76_856 ();
 FILLCELL_X2 FILLER_76_860 ();
 FILLCELL_X1 FILLER_76_862 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X32 FILLER_77_769 ();
 FILLCELL_X32 FILLER_77_801 ();
 FILLCELL_X16 FILLER_77_833 ();
 FILLCELL_X8 FILLER_77_849 ();
 FILLCELL_X4 FILLER_77_857 ();
 FILLCELL_X2 FILLER_77_861 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X32 FILLER_78_760 ();
 FILLCELL_X32 FILLER_78_792 ();
 FILLCELL_X32 FILLER_78_824 ();
 FILLCELL_X4 FILLER_78_856 ();
 FILLCELL_X2 FILLER_78_860 ();
 FILLCELL_X1 FILLER_78_862 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X32 FILLER_79_769 ();
 FILLCELL_X32 FILLER_79_801 ();
 FILLCELL_X16 FILLER_79_833 ();
 FILLCELL_X8 FILLER_79_849 ();
 FILLCELL_X4 FILLER_79_857 ();
 FILLCELL_X2 FILLER_79_861 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X32 FILLER_80_760 ();
 FILLCELL_X32 FILLER_80_792 ();
 FILLCELL_X32 FILLER_80_824 ();
 FILLCELL_X4 FILLER_80_856 ();
 FILLCELL_X2 FILLER_80_860 ();
 FILLCELL_X1 FILLER_80_862 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X32 FILLER_81_769 ();
 FILLCELL_X32 FILLER_81_801 ();
 FILLCELL_X16 FILLER_81_833 ();
 FILLCELL_X8 FILLER_81_849 ();
 FILLCELL_X4 FILLER_81_857 ();
 FILLCELL_X2 FILLER_81_861 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X32 FILLER_82_760 ();
 FILLCELL_X32 FILLER_82_792 ();
 FILLCELL_X32 FILLER_82_824 ();
 FILLCELL_X4 FILLER_82_856 ();
 FILLCELL_X2 FILLER_82_860 ();
 FILLCELL_X1 FILLER_82_862 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X32 FILLER_83_769 ();
 FILLCELL_X32 FILLER_83_801 ();
 FILLCELL_X16 FILLER_83_833 ();
 FILLCELL_X8 FILLER_83_849 ();
 FILLCELL_X4 FILLER_83_857 ();
 FILLCELL_X2 FILLER_83_861 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X32 FILLER_84_760 ();
 FILLCELL_X32 FILLER_84_792 ();
 FILLCELL_X32 FILLER_84_824 ();
 FILLCELL_X4 FILLER_84_856 ();
 FILLCELL_X2 FILLER_84_860 ();
 FILLCELL_X1 FILLER_84_862 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X32 FILLER_85_769 ();
 FILLCELL_X32 FILLER_85_801 ();
 FILLCELL_X16 FILLER_85_833 ();
 FILLCELL_X8 FILLER_85_849 ();
 FILLCELL_X4 FILLER_85_857 ();
 FILLCELL_X2 FILLER_85_861 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X32 FILLER_86_760 ();
 FILLCELL_X32 FILLER_86_792 ();
 FILLCELL_X32 FILLER_86_824 ();
 FILLCELL_X4 FILLER_86_856 ();
 FILLCELL_X2 FILLER_86_860 ();
 FILLCELL_X1 FILLER_86_862 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X32 FILLER_87_769 ();
 FILLCELL_X32 FILLER_87_801 ();
 FILLCELL_X16 FILLER_87_833 ();
 FILLCELL_X8 FILLER_87_849 ();
 FILLCELL_X4 FILLER_87_857 ();
 FILLCELL_X2 FILLER_87_861 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X32 FILLER_88_760 ();
 FILLCELL_X32 FILLER_88_792 ();
 FILLCELL_X32 FILLER_88_824 ();
 FILLCELL_X4 FILLER_88_856 ();
 FILLCELL_X2 FILLER_88_860 ();
 FILLCELL_X1 FILLER_88_862 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X32 FILLER_89_769 ();
 FILLCELL_X32 FILLER_89_801 ();
 FILLCELL_X16 FILLER_89_833 ();
 FILLCELL_X8 FILLER_89_849 ();
 FILLCELL_X4 FILLER_89_857 ();
 FILLCELL_X2 FILLER_89_861 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X32 FILLER_90_760 ();
 FILLCELL_X32 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_824 ();
 FILLCELL_X4 FILLER_90_856 ();
 FILLCELL_X2 FILLER_90_860 ();
 FILLCELL_X1 FILLER_90_862 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X32 FILLER_91_769 ();
 FILLCELL_X32 FILLER_91_801 ();
 FILLCELL_X16 FILLER_91_833 ();
 FILLCELL_X8 FILLER_91_849 ();
 FILLCELL_X4 FILLER_91_857 ();
 FILLCELL_X2 FILLER_91_861 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X32 FILLER_92_760 ();
 FILLCELL_X32 FILLER_92_792 ();
 FILLCELL_X32 FILLER_92_824 ();
 FILLCELL_X4 FILLER_92_856 ();
 FILLCELL_X2 FILLER_92_860 ();
 FILLCELL_X1 FILLER_92_862 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X32 FILLER_93_769 ();
 FILLCELL_X32 FILLER_93_801 ();
 FILLCELL_X16 FILLER_93_833 ();
 FILLCELL_X8 FILLER_93_849 ();
 FILLCELL_X4 FILLER_93_857 ();
 FILLCELL_X2 FILLER_93_861 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X32 FILLER_94_760 ();
 FILLCELL_X32 FILLER_94_792 ();
 FILLCELL_X32 FILLER_94_824 ();
 FILLCELL_X4 FILLER_94_856 ();
 FILLCELL_X2 FILLER_94_860 ();
 FILLCELL_X1 FILLER_94_862 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X32 FILLER_95_353 ();
 FILLCELL_X32 FILLER_95_385 ();
 FILLCELL_X32 FILLER_95_417 ();
 FILLCELL_X32 FILLER_95_449 ();
 FILLCELL_X32 FILLER_95_481 ();
 FILLCELL_X32 FILLER_95_513 ();
 FILLCELL_X32 FILLER_95_545 ();
 FILLCELL_X32 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_609 ();
 FILLCELL_X32 FILLER_95_641 ();
 FILLCELL_X32 FILLER_95_673 ();
 FILLCELL_X32 FILLER_95_705 ();
 FILLCELL_X32 FILLER_95_737 ();
 FILLCELL_X32 FILLER_95_769 ();
 FILLCELL_X32 FILLER_95_801 ();
 FILLCELL_X16 FILLER_95_833 ();
 FILLCELL_X8 FILLER_95_849 ();
 FILLCELL_X4 FILLER_95_857 ();
 FILLCELL_X2 FILLER_95_861 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X32 FILLER_96_760 ();
 FILLCELL_X32 FILLER_96_792 ();
 FILLCELL_X32 FILLER_96_824 ();
 FILLCELL_X4 FILLER_96_856 ();
 FILLCELL_X2 FILLER_96_860 ();
 FILLCELL_X1 FILLER_96_862 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X32 FILLER_97_321 ();
 FILLCELL_X32 FILLER_97_353 ();
 FILLCELL_X32 FILLER_97_385 ();
 FILLCELL_X32 FILLER_97_417 ();
 FILLCELL_X32 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_481 ();
 FILLCELL_X32 FILLER_97_513 ();
 FILLCELL_X32 FILLER_97_545 ();
 FILLCELL_X32 FILLER_97_577 ();
 FILLCELL_X32 FILLER_97_609 ();
 FILLCELL_X32 FILLER_97_641 ();
 FILLCELL_X32 FILLER_97_673 ();
 FILLCELL_X32 FILLER_97_705 ();
 FILLCELL_X32 FILLER_97_737 ();
 FILLCELL_X32 FILLER_97_769 ();
 FILLCELL_X32 FILLER_97_801 ();
 FILLCELL_X16 FILLER_97_833 ();
 FILLCELL_X8 FILLER_97_849 ();
 FILLCELL_X4 FILLER_97_857 ();
 FILLCELL_X2 FILLER_97_861 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X32 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_193 ();
 FILLCELL_X32 FILLER_98_225 ();
 FILLCELL_X32 FILLER_98_257 ();
 FILLCELL_X32 FILLER_98_289 ();
 FILLCELL_X32 FILLER_98_321 ();
 FILLCELL_X32 FILLER_98_353 ();
 FILLCELL_X32 FILLER_98_385 ();
 FILLCELL_X32 FILLER_98_417 ();
 FILLCELL_X32 FILLER_98_449 ();
 FILLCELL_X32 FILLER_98_481 ();
 FILLCELL_X32 FILLER_98_513 ();
 FILLCELL_X32 FILLER_98_545 ();
 FILLCELL_X32 FILLER_98_577 ();
 FILLCELL_X16 FILLER_98_609 ();
 FILLCELL_X4 FILLER_98_625 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X32 FILLER_98_824 ();
 FILLCELL_X4 FILLER_98_856 ();
 FILLCELL_X2 FILLER_98_860 ();
 FILLCELL_X1 FILLER_98_862 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X32 FILLER_99_769 ();
 FILLCELL_X32 FILLER_99_801 ();
 FILLCELL_X16 FILLER_99_833 ();
 FILLCELL_X8 FILLER_99_849 ();
 FILLCELL_X4 FILLER_99_857 ();
 FILLCELL_X2 FILLER_99_861 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X32 FILLER_100_760 ();
 FILLCELL_X32 FILLER_100_792 ();
 FILLCELL_X32 FILLER_100_824 ();
 FILLCELL_X4 FILLER_100_856 ();
 FILLCELL_X2 FILLER_100_860 ();
 FILLCELL_X1 FILLER_100_862 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X32 FILLER_101_769 ();
 FILLCELL_X32 FILLER_101_801 ();
 FILLCELL_X16 FILLER_101_833 ();
 FILLCELL_X8 FILLER_101_849 ();
 FILLCELL_X4 FILLER_101_857 ();
 FILLCELL_X2 FILLER_101_861 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X32 FILLER_102_792 ();
 FILLCELL_X32 FILLER_102_824 ();
 FILLCELL_X4 FILLER_102_856 ();
 FILLCELL_X2 FILLER_102_860 ();
 FILLCELL_X1 FILLER_102_862 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X32 FILLER_103_769 ();
 FILLCELL_X32 FILLER_103_801 ();
 FILLCELL_X16 FILLER_103_833 ();
 FILLCELL_X8 FILLER_103_849 ();
 FILLCELL_X4 FILLER_103_857 ();
 FILLCELL_X2 FILLER_103_861 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X32 FILLER_104_385 ();
 FILLCELL_X32 FILLER_104_417 ();
 FILLCELL_X32 FILLER_104_449 ();
 FILLCELL_X32 FILLER_104_481 ();
 FILLCELL_X32 FILLER_104_513 ();
 FILLCELL_X32 FILLER_104_545 ();
 FILLCELL_X32 FILLER_104_577 ();
 FILLCELL_X16 FILLER_104_609 ();
 FILLCELL_X4 FILLER_104_625 ();
 FILLCELL_X2 FILLER_104_629 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X32 FILLER_104_760 ();
 FILLCELL_X32 FILLER_104_792 ();
 FILLCELL_X32 FILLER_104_824 ();
 FILLCELL_X4 FILLER_104_856 ();
 FILLCELL_X2 FILLER_104_860 ();
 FILLCELL_X1 FILLER_104_862 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_385 ();
 FILLCELL_X32 FILLER_105_417 ();
 FILLCELL_X32 FILLER_105_449 ();
 FILLCELL_X32 FILLER_105_481 ();
 FILLCELL_X32 FILLER_105_513 ();
 FILLCELL_X32 FILLER_105_545 ();
 FILLCELL_X32 FILLER_105_577 ();
 FILLCELL_X32 FILLER_105_609 ();
 FILLCELL_X32 FILLER_105_641 ();
 FILLCELL_X32 FILLER_105_673 ();
 FILLCELL_X32 FILLER_105_705 ();
 FILLCELL_X32 FILLER_105_737 ();
 FILLCELL_X32 FILLER_105_769 ();
 FILLCELL_X32 FILLER_105_801 ();
 FILLCELL_X16 FILLER_105_833 ();
 FILLCELL_X8 FILLER_105_849 ();
 FILLCELL_X4 FILLER_105_857 ();
 FILLCELL_X2 FILLER_105_861 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X32 FILLER_106_481 ();
 FILLCELL_X32 FILLER_106_513 ();
 FILLCELL_X32 FILLER_106_545 ();
 FILLCELL_X32 FILLER_106_577 ();
 FILLCELL_X16 FILLER_106_609 ();
 FILLCELL_X4 FILLER_106_625 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X32 FILLER_106_792 ();
 FILLCELL_X32 FILLER_106_824 ();
 FILLCELL_X4 FILLER_106_856 ();
 FILLCELL_X2 FILLER_106_860 ();
 FILLCELL_X1 FILLER_106_862 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X32 FILLER_107_577 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X32 FILLER_107_801 ();
 FILLCELL_X16 FILLER_107_833 ();
 FILLCELL_X8 FILLER_107_849 ();
 FILLCELL_X4 FILLER_107_857 ();
 FILLCELL_X2 FILLER_107_861 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X32 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_760 ();
 FILLCELL_X32 FILLER_108_792 ();
 FILLCELL_X32 FILLER_108_824 ();
 FILLCELL_X4 FILLER_108_856 ();
 FILLCELL_X2 FILLER_108_860 ();
 FILLCELL_X1 FILLER_108_862 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X32 FILLER_109_385 ();
 FILLCELL_X32 FILLER_109_417 ();
 FILLCELL_X32 FILLER_109_449 ();
 FILLCELL_X32 FILLER_109_481 ();
 FILLCELL_X32 FILLER_109_513 ();
 FILLCELL_X32 FILLER_109_545 ();
 FILLCELL_X32 FILLER_109_577 ();
 FILLCELL_X32 FILLER_109_609 ();
 FILLCELL_X32 FILLER_109_641 ();
 FILLCELL_X32 FILLER_109_673 ();
 FILLCELL_X32 FILLER_109_705 ();
 FILLCELL_X32 FILLER_109_737 ();
 FILLCELL_X32 FILLER_109_769 ();
 FILLCELL_X32 FILLER_109_801 ();
 FILLCELL_X16 FILLER_109_833 ();
 FILLCELL_X8 FILLER_109_849 ();
 FILLCELL_X4 FILLER_109_857 ();
 FILLCELL_X2 FILLER_109_861 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X32 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_321 ();
 FILLCELL_X32 FILLER_110_353 ();
 FILLCELL_X32 FILLER_110_385 ();
 FILLCELL_X32 FILLER_110_417 ();
 FILLCELL_X32 FILLER_110_449 ();
 FILLCELL_X32 FILLER_110_481 ();
 FILLCELL_X32 FILLER_110_513 ();
 FILLCELL_X32 FILLER_110_545 ();
 FILLCELL_X32 FILLER_110_577 ();
 FILLCELL_X16 FILLER_110_609 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X32 FILLER_110_696 ();
 FILLCELL_X32 FILLER_110_728 ();
 FILLCELL_X32 FILLER_110_760 ();
 FILLCELL_X32 FILLER_110_792 ();
 FILLCELL_X32 FILLER_110_824 ();
 FILLCELL_X4 FILLER_110_856 ();
 FILLCELL_X2 FILLER_110_860 ();
 FILLCELL_X1 FILLER_110_862 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X32 FILLER_111_289 ();
 FILLCELL_X32 FILLER_111_321 ();
 FILLCELL_X32 FILLER_111_353 ();
 FILLCELL_X32 FILLER_111_385 ();
 FILLCELL_X32 FILLER_111_417 ();
 FILLCELL_X32 FILLER_111_449 ();
 FILLCELL_X32 FILLER_111_481 ();
 FILLCELL_X32 FILLER_111_513 ();
 FILLCELL_X32 FILLER_111_545 ();
 FILLCELL_X32 FILLER_111_577 ();
 FILLCELL_X32 FILLER_111_609 ();
 FILLCELL_X32 FILLER_111_641 ();
 FILLCELL_X32 FILLER_111_673 ();
 FILLCELL_X32 FILLER_111_705 ();
 FILLCELL_X32 FILLER_111_737 ();
 FILLCELL_X32 FILLER_111_769 ();
 FILLCELL_X32 FILLER_111_801 ();
 FILLCELL_X16 FILLER_111_833 ();
 FILLCELL_X8 FILLER_111_849 ();
 FILLCELL_X4 FILLER_111_857 ();
 FILLCELL_X2 FILLER_111_861 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X32 FILLER_112_225 ();
 FILLCELL_X32 FILLER_112_257 ();
 FILLCELL_X32 FILLER_112_289 ();
 FILLCELL_X32 FILLER_112_321 ();
 FILLCELL_X32 FILLER_112_353 ();
 FILLCELL_X32 FILLER_112_385 ();
 FILLCELL_X32 FILLER_112_417 ();
 FILLCELL_X32 FILLER_112_449 ();
 FILLCELL_X32 FILLER_112_481 ();
 FILLCELL_X32 FILLER_112_513 ();
 FILLCELL_X32 FILLER_112_545 ();
 FILLCELL_X32 FILLER_112_577 ();
 FILLCELL_X16 FILLER_112_609 ();
 FILLCELL_X4 FILLER_112_625 ();
 FILLCELL_X2 FILLER_112_629 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X32 FILLER_112_696 ();
 FILLCELL_X32 FILLER_112_728 ();
 FILLCELL_X32 FILLER_112_760 ();
 FILLCELL_X32 FILLER_112_792 ();
 FILLCELL_X32 FILLER_112_824 ();
 FILLCELL_X4 FILLER_112_856 ();
 FILLCELL_X2 FILLER_112_860 ();
 FILLCELL_X1 FILLER_112_862 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X32 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_193 ();
 FILLCELL_X32 FILLER_113_225 ();
 FILLCELL_X32 FILLER_113_257 ();
 FILLCELL_X32 FILLER_113_289 ();
 FILLCELL_X32 FILLER_113_321 ();
 FILLCELL_X32 FILLER_113_353 ();
 FILLCELL_X32 FILLER_113_385 ();
 FILLCELL_X32 FILLER_113_417 ();
 FILLCELL_X32 FILLER_113_449 ();
 FILLCELL_X32 FILLER_113_481 ();
 FILLCELL_X32 FILLER_113_513 ();
 FILLCELL_X32 FILLER_113_545 ();
 FILLCELL_X32 FILLER_113_577 ();
 FILLCELL_X32 FILLER_113_609 ();
 FILLCELL_X32 FILLER_113_641 ();
 FILLCELL_X32 FILLER_113_673 ();
 FILLCELL_X32 FILLER_113_705 ();
 FILLCELL_X32 FILLER_113_737 ();
 FILLCELL_X32 FILLER_113_769 ();
 FILLCELL_X32 FILLER_113_801 ();
 FILLCELL_X16 FILLER_113_833 ();
 FILLCELL_X8 FILLER_113_849 ();
 FILLCELL_X4 FILLER_113_857 ();
 FILLCELL_X2 FILLER_113_861 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X32 FILLER_114_225 ();
 FILLCELL_X32 FILLER_114_257 ();
 FILLCELL_X32 FILLER_114_289 ();
 FILLCELL_X32 FILLER_114_321 ();
 FILLCELL_X32 FILLER_114_353 ();
 FILLCELL_X32 FILLER_114_385 ();
 FILLCELL_X32 FILLER_114_417 ();
 FILLCELL_X32 FILLER_114_449 ();
 FILLCELL_X32 FILLER_114_481 ();
 FILLCELL_X32 FILLER_114_513 ();
 FILLCELL_X32 FILLER_114_545 ();
 FILLCELL_X32 FILLER_114_577 ();
 FILLCELL_X16 FILLER_114_609 ();
 FILLCELL_X4 FILLER_114_625 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X32 FILLER_114_664 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X32 FILLER_114_760 ();
 FILLCELL_X32 FILLER_114_792 ();
 FILLCELL_X32 FILLER_114_824 ();
 FILLCELL_X4 FILLER_114_856 ();
 FILLCELL_X2 FILLER_114_860 ();
 FILLCELL_X1 FILLER_114_862 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X32 FILLER_115_321 ();
 FILLCELL_X32 FILLER_115_353 ();
 FILLCELL_X32 FILLER_115_385 ();
 FILLCELL_X32 FILLER_115_417 ();
 FILLCELL_X32 FILLER_115_449 ();
 FILLCELL_X8 FILLER_115_481 ();
 FILLCELL_X4 FILLER_115_489 ();
 FILLCELL_X32 FILLER_115_496 ();
 FILLCELL_X32 FILLER_115_531 ();
 FILLCELL_X16 FILLER_115_563 ();
 FILLCELL_X8 FILLER_115_579 ();
 FILLCELL_X32 FILLER_115_590 ();
 FILLCELL_X32 FILLER_115_622 ();
 FILLCELL_X32 FILLER_115_654 ();
 FILLCELL_X32 FILLER_115_686 ();
 FILLCELL_X32 FILLER_115_718 ();
 FILLCELL_X32 FILLER_115_750 ();
 FILLCELL_X32 FILLER_115_782 ();
 FILLCELL_X32 FILLER_115_814 ();
 FILLCELL_X16 FILLER_115_846 ();
 FILLCELL_X1 FILLER_115_862 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X32 FILLER_116_321 ();
 FILLCELL_X32 FILLER_116_353 ();
 FILLCELL_X32 FILLER_116_385 ();
 FILLCELL_X32 FILLER_116_417 ();
 FILLCELL_X4 FILLER_116_449 ();
 FILLCELL_X2 FILLER_116_453 ();
 FILLCELL_X1 FILLER_116_455 ();
 FILLCELL_X4 FILLER_116_459 ();
 FILLCELL_X2 FILLER_116_463 ();
 FILLCELL_X16 FILLER_116_478 ();
 FILLCELL_X2 FILLER_116_494 ();
 FILLCELL_X4 FILLER_116_499 ();
 FILLCELL_X2 FILLER_116_503 ();
 FILLCELL_X4 FILLER_116_508 ();
 FILLCELL_X1 FILLER_116_512 ();
 FILLCELL_X16 FILLER_116_517 ();
 FILLCELL_X2 FILLER_116_533 ();
 FILLCELL_X16 FILLER_116_538 ();
 FILLCELL_X8 FILLER_116_554 ();
 FILLCELL_X1 FILLER_116_562 ();
 FILLCELL_X4 FILLER_116_566 ();
 FILLCELL_X2 FILLER_116_570 ();
 FILLCELL_X32 FILLER_116_575 ();
 FILLCELL_X16 FILLER_116_607 ();
 FILLCELL_X8 FILLER_116_623 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X32 FILLER_116_728 ();
 FILLCELL_X32 FILLER_116_760 ();
 FILLCELL_X32 FILLER_116_792 ();
 FILLCELL_X32 FILLER_116_824 ();
 FILLCELL_X4 FILLER_116_856 ();
 FILLCELL_X2 FILLER_116_860 ();
 FILLCELL_X1 FILLER_116_862 ();
endmodule
