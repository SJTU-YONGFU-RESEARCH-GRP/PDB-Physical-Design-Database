module configurable_lfsr (clk,
    enable,
    load_seed,
    rst_n,
    serial_out,
    parallel_out,
    seed,
    tap_pattern);
 input clk;
 input enable;
 input load_seed;
 input rst_n;
 output serial_out;
 output [7:0] parallel_out;
 input [7:0] seed;
 input [7:0] tap_pattern;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X2 _059_ (.A(net1),
    .ZN(_008_));
 CLKBUF_X3 _060_ (.A(load_seed),
    .Z(_009_));
 INV_X2 _061_ (.A(_009_),
    .ZN(_010_));
 NOR2_X1 _062_ (.A1(_010_),
    .A2(net2),
    .ZN(_011_));
 CLKBUF_X3 _063_ (.A(enable),
    .Z(_012_));
 MUX2_X1 _064_ (.A(net26),
    .B(net19),
    .S(_012_),
    .Z(_013_));
 NOR2_X1 _065_ (.A1(_009_),
    .A2(_013_),
    .ZN(_014_));
 NOR3_X1 _066_ (.A1(_008_),
    .A2(_011_),
    .A3(_014_),
    .ZN(_000_));
 NOR2_X1 _067_ (.A1(_010_),
    .A2(net3),
    .ZN(_015_));
 MUX2_X1 _068_ (.A(net19),
    .B(net20),
    .S(_012_),
    .Z(_016_));
 NOR2_X1 _069_ (.A1(_009_),
    .A2(_016_),
    .ZN(_017_));
 NOR3_X1 _070_ (.A1(_008_),
    .A2(_015_),
    .A3(_017_),
    .ZN(_001_));
 NOR2_X1 _071_ (.A1(_010_),
    .A2(net4),
    .ZN(_018_));
 MUX2_X1 _072_ (.A(net20),
    .B(net21),
    .S(_012_),
    .Z(_019_));
 NOR2_X1 _073_ (.A1(_009_),
    .A2(_019_),
    .ZN(_020_));
 NOR3_X1 _074_ (.A1(_008_),
    .A2(_018_),
    .A3(_020_),
    .ZN(_002_));
 NOR2_X1 _075_ (.A1(_010_),
    .A2(net5),
    .ZN(_021_));
 MUX2_X1 _076_ (.A(net21),
    .B(net22),
    .S(_012_),
    .Z(_022_));
 NOR2_X1 _077_ (.A1(_009_),
    .A2(_022_),
    .ZN(_023_));
 NOR3_X1 _078_ (.A1(_008_),
    .A2(_021_),
    .A3(_023_),
    .ZN(_003_));
 NOR2_X1 _079_ (.A1(_010_),
    .A2(net6),
    .ZN(_024_));
 MUX2_X1 _080_ (.A(net22),
    .B(net23),
    .S(_012_),
    .Z(_025_));
 NOR2_X1 _081_ (.A1(_009_),
    .A2(_025_),
    .ZN(_026_));
 NOR3_X1 _082_ (.A1(_008_),
    .A2(_024_),
    .A3(_026_),
    .ZN(_004_));
 NOR2_X1 _083_ (.A1(_010_),
    .A2(net7),
    .ZN(_027_));
 MUX2_X1 _084_ (.A(net23),
    .B(net24),
    .S(_012_),
    .Z(_028_));
 NOR2_X1 _085_ (.A1(_009_),
    .A2(_028_),
    .ZN(_029_));
 NOR3_X1 _086_ (.A1(_008_),
    .A2(_027_),
    .A3(_029_),
    .ZN(_005_));
 NOR2_X1 _087_ (.A1(_010_),
    .A2(net8),
    .ZN(_030_));
 MUX2_X1 _088_ (.A(net24),
    .B(net25),
    .S(_012_),
    .Z(_031_));
 NOR2_X1 _089_ (.A1(_009_),
    .A2(_031_),
    .ZN(_032_));
 NOR3_X1 _090_ (.A1(_008_),
    .A2(_030_),
    .A3(_032_),
    .ZN(_006_));
 NOR2_X1 _091_ (.A1(_009_),
    .A2(_012_),
    .ZN(_033_));
 AOI22_X1 _092_ (.A1(_009_),
    .A2(net9),
    .B1(_033_),
    .B2(net25),
    .ZN(_034_));
 NAND2_X1 _093_ (.A1(net23),
    .A2(net15),
    .ZN(_035_));
 NAND2_X1 _094_ (.A1(net21),
    .A2(net13),
    .ZN(_036_));
 XOR2_X1 _095_ (.A(_035_),
    .B(_036_),
    .Z(_037_));
 NAND2_X1 _096_ (.A1(net24),
    .A2(net16),
    .ZN(_038_));
 NAND2_X1 _097_ (.A1(net22),
    .A2(net14),
    .ZN(_039_));
 XNOR2_X1 _098_ (.A(_038_),
    .B(_039_),
    .ZN(_040_));
 XNOR2_X1 _099_ (.A(_037_),
    .B(_040_),
    .ZN(_041_));
 NAND2_X1 _100_ (.A1(net19),
    .A2(net11),
    .ZN(_042_));
 NAND2_X1 _101_ (.A1(net10),
    .A2(net26),
    .ZN(_043_));
 XOR2_X1 _102_ (.A(_042_),
    .B(_043_),
    .Z(_044_));
 NAND2_X1 _103_ (.A1(net25),
    .A2(net17),
    .ZN(_045_));
 NAND2_X1 _104_ (.A1(net20),
    .A2(net12),
    .ZN(_046_));
 XNOR2_X1 _105_ (.A(_045_),
    .B(_046_),
    .ZN(_047_));
 XNOR2_X1 _106_ (.A(_044_),
    .B(_047_),
    .ZN(_048_));
 XNOR2_X1 _107_ (.A(_041_),
    .B(_048_),
    .ZN(_049_));
 NAND3_X1 _108_ (.A1(_010_),
    .A2(_012_),
    .A3(net1),
    .ZN(_050_));
 OAI22_X1 _109_ (.A1(_008_),
    .A2(_034_),
    .B1(_049_),
    .B2(_050_),
    .ZN(_007_));
 BUF_X1 _110_ (.A(net26),
    .Z(net18));
 DFF_X1 \shift_reg[0]$_SDFFE_PN0P_  (.D(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net26),
    .QN(_058_));
 DFF_X1 \shift_reg[1]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net19),
    .QN(_057_));
 DFF_X1 \shift_reg[2]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net20),
    .QN(_056_));
 DFF_X1 \shift_reg[3]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net21),
    .QN(_055_));
 DFF_X1 \shift_reg[4]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net22),
    .QN(_054_));
 DFF_X1 \shift_reg[5]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net23),
    .QN(_053_));
 DFF_X1 \shift_reg[6]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net24),
    .QN(_052_));
 DFF_X1 \shift_reg[7]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net25),
    .QN(_051_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_41 ();
 BUF_X1 input1 (.A(rst_n),
    .Z(net1));
 BUF_X1 input2 (.A(seed[0]),
    .Z(net2));
 BUF_X1 input3 (.A(seed[1]),
    .Z(net3));
 BUF_X1 input4 (.A(seed[2]),
    .Z(net4));
 BUF_X1 input5 (.A(seed[3]),
    .Z(net5));
 BUF_X1 input6 (.A(seed[4]),
    .Z(net6));
 BUF_X1 input7 (.A(seed[5]),
    .Z(net7));
 BUF_X1 input8 (.A(seed[6]),
    .Z(net8));
 BUF_X1 input9 (.A(seed[7]),
    .Z(net9));
 BUF_X1 input10 (.A(tap_pattern[0]),
    .Z(net10));
 BUF_X1 input11 (.A(tap_pattern[1]),
    .Z(net11));
 BUF_X1 input12 (.A(tap_pattern[2]),
    .Z(net12));
 BUF_X1 input13 (.A(tap_pattern[3]),
    .Z(net13));
 BUF_X1 input14 (.A(tap_pattern[4]),
    .Z(net14));
 BUF_X1 input15 (.A(tap_pattern[5]),
    .Z(net15));
 BUF_X1 input16 (.A(tap_pattern[6]),
    .Z(net16));
 BUF_X1 input17 (.A(tap_pattern[7]),
    .Z(net17));
 BUF_X1 output18 (.A(net18),
    .Z(parallel_out[0]));
 BUF_X1 output19 (.A(net19),
    .Z(parallel_out[1]));
 BUF_X1 output20 (.A(net20),
    .Z(parallel_out[2]));
 BUF_X1 output21 (.A(net21),
    .Z(parallel_out[3]));
 BUF_X1 output22 (.A(net22),
    .Z(parallel_out[4]));
 BUF_X1 output23 (.A(net23),
    .Z(parallel_out[5]));
 BUF_X1 output24 (.A(net24),
    .Z(parallel_out[6]));
 BUF_X1 output25 (.A(net25),
    .Z(parallel_out[7]));
 BUF_X1 output26 (.A(net26),
    .Z(serial_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_33 ();
 FILLCELL_X4 FILLER_0_41 ();
 FILLCELL_X1 FILLER_0_45 ();
 FILLCELL_X4 FILLER_0_49 ();
 FILLCELL_X8 FILLER_0_56 ();
 FILLCELL_X1 FILLER_0_64 ();
 FILLCELL_X8 FILLER_0_68 ();
 FILLCELL_X4 FILLER_0_76 ();
 FILLCELL_X32 FILLER_0_83 ();
 FILLCELL_X32 FILLER_0_115 ();
 FILLCELL_X8 FILLER_0_147 ();
 FILLCELL_X4 FILLER_0_155 ();
 FILLCELL_X2 FILLER_0_159 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X4 FILLER_1_65 ();
 FILLCELL_X16 FILLER_1_75 ();
 FILLCELL_X8 FILLER_1_91 ();
 FILLCELL_X2 FILLER_1_99 ();
 FILLCELL_X1 FILLER_1_101 ();
 FILLCELL_X32 FILLER_1_105 ();
 FILLCELL_X16 FILLER_1_137 ();
 FILLCELL_X8 FILLER_1_153 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X4 FILLER_2_49 ();
 FILLCELL_X2 FILLER_2_53 ();
 FILLCELL_X8 FILLER_2_58 ();
 FILLCELL_X4 FILLER_2_66 ();
 FILLCELL_X2 FILLER_2_70 ();
 FILLCELL_X32 FILLER_2_75 ();
 FILLCELL_X32 FILLER_2_107 ();
 FILLCELL_X16 FILLER_2_139 ();
 FILLCELL_X4 FILLER_2_155 ();
 FILLCELL_X2 FILLER_2_159 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X8 FILLER_5_33 ();
 FILLCELL_X4 FILLER_5_41 ();
 FILLCELL_X1 FILLER_5_45 ();
 FILLCELL_X16 FILLER_5_49 ();
 FILLCELL_X8 FILLER_5_65 ();
 FILLCELL_X4 FILLER_5_73 ();
 FILLCELL_X2 FILLER_5_77 ();
 FILLCELL_X32 FILLER_5_82 ();
 FILLCELL_X32 FILLER_5_114 ();
 FILLCELL_X8 FILLER_5_146 ();
 FILLCELL_X4 FILLER_5_154 ();
 FILLCELL_X2 FILLER_5_158 ();
 FILLCELL_X1 FILLER_5_160 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X8 FILLER_6_33 ();
 FILLCELL_X4 FILLER_6_41 ();
 FILLCELL_X2 FILLER_6_45 ();
 FILLCELL_X4 FILLER_6_51 ();
 FILLCELL_X1 FILLER_6_55 ();
 FILLCELL_X16 FILLER_6_59 ();
 FILLCELL_X2 FILLER_6_75 ();
 FILLCELL_X1 FILLER_6_77 ();
 FILLCELL_X4 FILLER_6_82 ();
 FILLCELL_X2 FILLER_6_89 ();
 FILLCELL_X1 FILLER_6_91 ();
 FILLCELL_X32 FILLER_6_95 ();
 FILLCELL_X16 FILLER_6_127 ();
 FILLCELL_X4 FILLER_6_143 ();
 FILLCELL_X1 FILLER_6_147 ();
 FILLCELL_X8 FILLER_6_151 ();
 FILLCELL_X2 FILLER_6_159 ();
 FILLCELL_X8 FILLER_7_4 ();
 FILLCELL_X4 FILLER_7_12 ();
 FILLCELL_X2 FILLER_7_23 ();
 FILLCELL_X4 FILLER_7_35 ();
 FILLCELL_X1 FILLER_7_63 ();
 FILLCELL_X1 FILLER_7_81 ();
 FILLCELL_X1 FILLER_7_89 ();
 FILLCELL_X32 FILLER_7_94 ();
 FILLCELL_X8 FILLER_7_126 ();
 FILLCELL_X2 FILLER_7_134 ();
 FILLCELL_X16 FILLER_7_139 ();
 FILLCELL_X4 FILLER_7_155 ();
 FILLCELL_X2 FILLER_7_159 ();
 FILLCELL_X2 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_3 ();
 FILLCELL_X32 FILLER_8_27 ();
 FILLCELL_X4 FILLER_8_59 ();
 FILLCELL_X4 FILLER_8_69 ();
 FILLCELL_X2 FILLER_8_73 ();
 FILLCELL_X32 FILLER_8_102 ();
 FILLCELL_X8 FILLER_8_134 ();
 FILLCELL_X2 FILLER_8_142 ();
 FILLCELL_X1 FILLER_8_144 ();
 FILLCELL_X8 FILLER_8_148 ();
 FILLCELL_X4 FILLER_8_156 ();
 FILLCELL_X1 FILLER_8_160 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X2 FILLER_9_49 ();
 FILLCELL_X1 FILLER_9_51 ();
 FILLCELL_X4 FILLER_9_58 ();
 FILLCELL_X16 FILLER_9_68 ();
 FILLCELL_X4 FILLER_9_84 ();
 FILLCELL_X2 FILLER_9_94 ();
 FILLCELL_X1 FILLER_9_96 ();
 FILLCELL_X32 FILLER_9_100 ();
 FILLCELL_X8 FILLER_9_132 ();
 FILLCELL_X4 FILLER_9_140 ();
 FILLCELL_X2 FILLER_9_144 ();
 FILLCELL_X8 FILLER_9_149 ();
 FILLCELL_X4 FILLER_9_157 ();
 FILLCELL_X1 FILLER_10_1 ();
 FILLCELL_X8 FILLER_10_8 ();
 FILLCELL_X2 FILLER_10_16 ();
 FILLCELL_X4 FILLER_10_21 ();
 FILLCELL_X32 FILLER_10_37 ();
 FILLCELL_X16 FILLER_10_69 ();
 FILLCELL_X8 FILLER_10_85 ();
 FILLCELL_X2 FILLER_10_93 ();
 FILLCELL_X32 FILLER_10_100 ();
 FILLCELL_X4 FILLER_10_132 ();
 FILLCELL_X2 FILLER_10_136 ();
 FILLCELL_X1 FILLER_10_138 ();
 FILLCELL_X8 FILLER_10_151 ();
 FILLCELL_X2 FILLER_10_159 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_9 ();
 FILLCELL_X8 FILLER_11_36 ();
 FILLCELL_X2 FILLER_11_44 ();
 FILLCELL_X1 FILLER_11_46 ();
 FILLCELL_X4 FILLER_11_50 ();
 FILLCELL_X16 FILLER_11_66 ();
 FILLCELL_X4 FILLER_11_82 ();
 FILLCELL_X2 FILLER_11_86 ();
 FILLCELL_X1 FILLER_11_88 ();
 FILLCELL_X2 FILLER_11_99 ();
 FILLCELL_X32 FILLER_11_108 ();
 FILLCELL_X4 FILLER_11_140 ();
 FILLCELL_X2 FILLER_11_144 ();
 FILLCELL_X2 FILLER_11_149 ();
 FILLCELL_X4 FILLER_11_154 ();
 FILLCELL_X2 FILLER_11_158 ();
 FILLCELL_X1 FILLER_11_160 ();
 FILLCELL_X2 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_3 ();
 FILLCELL_X4 FILLER_12_7 ();
 FILLCELL_X1 FILLER_12_11 ();
 FILLCELL_X1 FILLER_12_20 ();
 FILLCELL_X16 FILLER_12_25 ();
 FILLCELL_X8 FILLER_12_41 ();
 FILLCELL_X4 FILLER_12_49 ();
 FILLCELL_X2 FILLER_12_53 ();
 FILLCELL_X1 FILLER_12_55 ();
 FILLCELL_X16 FILLER_12_63 ();
 FILLCELL_X4 FILLER_12_79 ();
 FILLCELL_X1 FILLER_12_83 ();
 FILLCELL_X32 FILLER_12_108 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X16 FILLER_13_33 ();
 FILLCELL_X2 FILLER_13_49 ();
 FILLCELL_X1 FILLER_13_51 ();
 FILLCELL_X2 FILLER_13_69 ();
 FILLCELL_X32 FILLER_13_95 ();
 FILLCELL_X16 FILLER_13_127 ();
 FILLCELL_X4 FILLER_13_143 ();
 FILLCELL_X2 FILLER_13_147 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X16 FILLER_14_33 ();
 FILLCELL_X4 FILLER_14_49 ();
 FILLCELL_X2 FILLER_14_53 ();
 FILLCELL_X1 FILLER_14_55 ();
 FILLCELL_X16 FILLER_14_59 ();
 FILLCELL_X4 FILLER_14_75 ();
 FILLCELL_X2 FILLER_14_79 ();
 FILLCELL_X1 FILLER_14_81 ();
 FILLCELL_X2 FILLER_14_87 ();
 FILLCELL_X32 FILLER_14_92 ();
 FILLCELL_X32 FILLER_14_124 ();
 FILLCELL_X4 FILLER_14_156 ();
 FILLCELL_X1 FILLER_14_160 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X16 FILLER_20_33 ();
 FILLCELL_X4 FILLER_20_49 ();
 FILLCELL_X2 FILLER_20_53 ();
 FILLCELL_X16 FILLER_20_58 ();
 FILLCELL_X8 FILLER_20_74 ();
 FILLCELL_X4 FILLER_20_82 ();
 FILLCELL_X2 FILLER_20_86 ();
 FILLCELL_X8 FILLER_20_91 ();
 FILLCELL_X2 FILLER_20_99 ();
 FILLCELL_X32 FILLER_20_104 ();
 FILLCELL_X16 FILLER_20_136 ();
 FILLCELL_X8 FILLER_20_152 ();
 FILLCELL_X1 FILLER_20_160 ();
endmodule
