module uart (clk,
    m_axis_tready,
    m_axis_tvalid,
    rst,
    rx_busy,
    rx_frame_error,
    rx_overrun_error,
    rxd,
    s_axis_tready,
    s_axis_tvalid,
    tx_busy,
    txd,
    m_axis_tdata,
    prescale,
    s_axis_tdata);
 input clk;
 input m_axis_tready;
 output m_axis_tvalid;
 input rst;
 output rx_busy;
 output rx_frame_error;
 output rx_overrun_error;
 input rxd;
 output s_axis_tready;
 input s_axis_tvalid;
 output tx_busy;
 output txd;
 output [7:0] m_axis_tdata;
 input [15:0] prescale;
 input [7:0] s_axis_tdata;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire \uart_rx_inst.bit_cnt[0] ;
 wire \uart_rx_inst.bit_cnt[1] ;
 wire \uart_rx_inst.bit_cnt[2] ;
 wire \uart_rx_inst.bit_cnt[3] ;
 wire \uart_rx_inst.data_reg[0] ;
 wire \uart_rx_inst.data_reg[1] ;
 wire \uart_rx_inst.data_reg[2] ;
 wire \uart_rx_inst.data_reg[3] ;
 wire \uart_rx_inst.data_reg[4] ;
 wire \uart_rx_inst.data_reg[5] ;
 wire \uart_rx_inst.data_reg[6] ;
 wire \uart_rx_inst.data_reg[7] ;
 wire \uart_rx_inst.prescale_reg[0] ;
 wire \uart_rx_inst.prescale_reg[10] ;
 wire \uart_rx_inst.prescale_reg[11] ;
 wire \uart_rx_inst.prescale_reg[12] ;
 wire \uart_rx_inst.prescale_reg[13] ;
 wire \uart_rx_inst.prescale_reg[14] ;
 wire \uart_rx_inst.prescale_reg[15] ;
 wire \uart_rx_inst.prescale_reg[16] ;
 wire \uart_rx_inst.prescale_reg[17] ;
 wire \uart_rx_inst.prescale_reg[18] ;
 wire \uart_rx_inst.prescale_reg[1] ;
 wire \uart_rx_inst.prescale_reg[2] ;
 wire \uart_rx_inst.prescale_reg[3] ;
 wire \uart_rx_inst.prescale_reg[4] ;
 wire \uart_rx_inst.prescale_reg[5] ;
 wire \uart_rx_inst.prescale_reg[6] ;
 wire \uart_rx_inst.prescale_reg[7] ;
 wire \uart_rx_inst.prescale_reg[8] ;
 wire \uart_rx_inst.prescale_reg[9] ;
 wire \uart_rx_inst.rxd_reg ;
 wire \uart_tx_inst.bit_cnt[0] ;
 wire \uart_tx_inst.bit_cnt[1] ;
 wire \uart_tx_inst.bit_cnt[2] ;
 wire \uart_tx_inst.bit_cnt[3] ;
 wire \uart_tx_inst.data_reg[0] ;
 wire \uart_tx_inst.data_reg[1] ;
 wire \uart_tx_inst.data_reg[2] ;
 wire \uart_tx_inst.data_reg[3] ;
 wire \uart_tx_inst.data_reg[4] ;
 wire \uart_tx_inst.data_reg[5] ;
 wire \uart_tx_inst.data_reg[6] ;
 wire \uart_tx_inst.data_reg[7] ;
 wire \uart_tx_inst.data_reg[8] ;
 wire \uart_tx_inst.prescale_reg[0] ;
 wire \uart_tx_inst.prescale_reg[10] ;
 wire \uart_tx_inst.prescale_reg[11] ;
 wire \uart_tx_inst.prescale_reg[12] ;
 wire \uart_tx_inst.prescale_reg[13] ;
 wire \uart_tx_inst.prescale_reg[14] ;
 wire \uart_tx_inst.prescale_reg[15] ;
 wire \uart_tx_inst.prescale_reg[16] ;
 wire \uart_tx_inst.prescale_reg[17] ;
 wire \uart_tx_inst.prescale_reg[18] ;
 wire \uart_tx_inst.prescale_reg[1] ;
 wire \uart_tx_inst.prescale_reg[2] ;
 wire \uart_tx_inst.prescale_reg[3] ;
 wire \uart_tx_inst.prescale_reg[4] ;
 wire \uart_tx_inst.prescale_reg[5] ;
 wire \uart_tx_inst.prescale_reg[6] ;
 wire \uart_tx_inst.prescale_reg[7] ;
 wire \uart_tx_inst.prescale_reg[8] ;
 wire \uart_tx_inst.prescale_reg[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 BUF_X2 _0608_ (.A(prescale[0]),
    .Z(_0081_));
 INV_X1 _0609_ (.A(_0081_),
    .ZN(_0592_));
 INV_X1 _0610_ (.A(net6),
    .ZN(_0593_));
 BUF_X4 _0611_ (.A(rst),
    .Z(_0082_));
 INV_X4 _0612_ (.A(_0082_),
    .ZN(_0083_));
 BUF_X2 _0613_ (.A(\uart_rx_inst.bit_cnt[2] ),
    .Z(_0084_));
 CLKBUF_X2 _0614_ (.A(_0602_),
    .Z(_0085_));
 NOR2_X1 _0615_ (.A1(_0600_),
    .A2(_0085_),
    .ZN(_0086_));
 OAI21_X2 _0616_ (.A(\uart_rx_inst.bit_cnt[3] ),
    .B1(_0084_),
    .B2(_0086_),
    .ZN(_0087_));
 NOR2_X2 _0617_ (.A1(\uart_rx_inst.bit_cnt[3] ),
    .A2(_0084_),
    .ZN(_0088_));
 BUF_X2 _0618_ (.A(_0000_),
    .Z(_0089_));
 INV_X1 _0619_ (.A(_0089_),
    .ZN(_0090_));
 BUF_X1 _0620_ (.A(_0598_),
    .Z(_0091_));
 AND2_X1 _0621_ (.A1(_0090_),
    .A2(_0091_),
    .ZN(_0092_));
 NOR2_X1 _0622_ (.A1(\uart_rx_inst.bit_cnt[1] ),
    .A2(_0091_),
    .ZN(_0093_));
 OAI21_X4 _0623_ (.A(_0088_),
    .B1(_0092_),
    .B2(_0093_),
    .ZN(_0094_));
 NOR2_X4 _0624_ (.A1(\uart_rx_inst.prescale_reg[4] ),
    .A2(\uart_rx_inst.prescale_reg[3] ),
    .ZN(_0095_));
 BUF_X2 _0625_ (.A(\uart_rx_inst.prescale_reg[2] ),
    .Z(_0096_));
 NOR3_X4 _0626_ (.A1(_0096_),
    .A2(\uart_rx_inst.prescale_reg[1] ),
    .A3(\uart_rx_inst.prescale_reg[0] ),
    .ZN(_0097_));
 BUF_X2 _0627_ (.A(\uart_rx_inst.prescale_reg[5] ),
    .Z(_0098_));
 NOR4_X4 _0628_ (.A1(\uart_rx_inst.prescale_reg[7] ),
    .A2(\uart_rx_inst.prescale_reg[8] ),
    .A3(\uart_rx_inst.prescale_reg[6] ),
    .A4(_0098_),
    .ZN(_0099_));
 NOR2_X2 _0629_ (.A1(\uart_rx_inst.prescale_reg[9] ),
    .A2(\uart_rx_inst.prescale_reg[10] ),
    .ZN(_0100_));
 NAND4_X4 _0630_ (.A1(_0095_),
    .A2(_0097_),
    .A3(_0099_),
    .A4(_0100_),
    .ZN(_0101_));
 BUF_X1 _0631_ (.A(\uart_rx_inst.prescale_reg[14] ),
    .Z(_0102_));
 BUF_X2 _0632_ (.A(\uart_rx_inst.prescale_reg[11] ),
    .Z(_0103_));
 OR3_X2 _0633_ (.A1(\uart_rx_inst.prescale_reg[13] ),
    .A2(_0103_),
    .A3(\uart_rx_inst.prescale_reg[12] ),
    .ZN(_0104_));
 OR3_X1 _0634_ (.A1(\uart_rx_inst.prescale_reg[17] ),
    .A2(\uart_rx_inst.prescale_reg[18] ),
    .A3(\uart_rx_inst.prescale_reg[16] ),
    .ZN(_0105_));
 OR4_X2 _0635_ (.A1(\uart_rx_inst.prescale_reg[15] ),
    .A2(_0102_),
    .A3(_0104_),
    .A4(_0105_),
    .ZN(_0106_));
 NOR2_X4 _0636_ (.A1(_0101_),
    .A2(_0106_),
    .ZN(_0107_));
 NAND4_X4 _0637_ (.A1(_0083_),
    .A2(_0087_),
    .A3(_0094_),
    .A4(_0107_),
    .ZN(_0108_));
 BUF_X2 _0638_ (.A(_0108_),
    .Z(_0109_));
 NAND2_X1 _0639_ (.A1(\uart_rx_inst.data_reg[0] ),
    .A2(_0109_),
    .ZN(_0110_));
 NAND2_X1 _0640_ (.A1(_0091_),
    .A2(_0088_),
    .ZN(_0111_));
 CLKBUF_X3 _0641_ (.A(_0111_),
    .Z(_0112_));
 CLKBUF_X3 _0642_ (.A(_0112_),
    .Z(_0113_));
 NAND2_X1 _0643_ (.A1(\uart_rx_inst.data_reg[1] ),
    .A2(_0113_),
    .ZN(_0114_));
 OAI21_X1 _0644_ (.A(_0110_),
    .B1(_0114_),
    .B2(_0109_),
    .ZN(_0007_));
 NAND2_X1 _0645_ (.A1(\uart_rx_inst.data_reg[1] ),
    .A2(_0109_),
    .ZN(_0115_));
 NAND2_X1 _0646_ (.A1(\uart_rx_inst.data_reg[2] ),
    .A2(_0113_),
    .ZN(_0116_));
 OAI21_X1 _0647_ (.A(_0115_),
    .B1(_0116_),
    .B2(_0109_),
    .ZN(_0008_));
 NAND2_X1 _0648_ (.A1(\uart_rx_inst.data_reg[2] ),
    .A2(_0109_),
    .ZN(_0117_));
 NAND2_X1 _0649_ (.A1(\uart_rx_inst.data_reg[3] ),
    .A2(_0113_),
    .ZN(_0118_));
 OAI21_X1 _0650_ (.A(_0117_),
    .B1(_0118_),
    .B2(_0109_),
    .ZN(_0009_));
 NAND2_X1 _0651_ (.A1(\uart_rx_inst.data_reg[3] ),
    .A2(_0108_),
    .ZN(_0119_));
 NAND2_X1 _0652_ (.A1(\uart_rx_inst.data_reg[4] ),
    .A2(_0113_),
    .ZN(_0120_));
 OAI21_X1 _0653_ (.A(_0119_),
    .B1(_0120_),
    .B2(_0109_),
    .ZN(_0010_));
 NAND2_X1 _0654_ (.A1(\uart_rx_inst.data_reg[4] ),
    .A2(_0108_),
    .ZN(_0121_));
 NAND2_X1 _0655_ (.A1(\uart_rx_inst.data_reg[5] ),
    .A2(_0113_),
    .ZN(_0122_));
 OAI21_X1 _0656_ (.A(_0121_),
    .B1(_0122_),
    .B2(_0109_),
    .ZN(_0011_));
 NAND2_X1 _0657_ (.A1(\uart_rx_inst.data_reg[5] ),
    .A2(_0108_),
    .ZN(_0123_));
 NAND2_X1 _0658_ (.A1(\uart_rx_inst.data_reg[6] ),
    .A2(_0113_),
    .ZN(_0124_));
 OAI21_X1 _0659_ (.A(_0123_),
    .B1(_0124_),
    .B2(_0109_),
    .ZN(_0012_));
 NAND2_X1 _0660_ (.A1(\uart_rx_inst.data_reg[6] ),
    .A2(_0108_),
    .ZN(_0125_));
 NAND2_X1 _0661_ (.A1(\uart_rx_inst.data_reg[7] ),
    .A2(_0113_),
    .ZN(_0126_));
 OAI21_X1 _0662_ (.A(_0125_),
    .B1(_0126_),
    .B2(_0109_),
    .ZN(_0013_));
 INV_X1 _0663_ (.A(\uart_rx_inst.rxd_reg ),
    .ZN(_0127_));
 AND2_X2 _0664_ (.A1(_0091_),
    .A2(_0088_),
    .ZN(_0128_));
 CLKBUF_X3 _0665_ (.A(_0128_),
    .Z(_0129_));
 NOR2_X1 _0666_ (.A1(_0127_),
    .A2(_0129_),
    .ZN(_0130_));
 MUX2_X1 _0667_ (.A(_0130_),
    .B(\uart_rx_inst.data_reg[7] ),
    .S(_0108_),
    .Z(_0014_));
 BUF_X2 _0668_ (.A(\uart_tx_inst.bit_cnt[2] ),
    .Z(_0131_));
 CLKBUF_X3 _0669_ (.A(\uart_tx_inst.bit_cnt[1] ),
    .Z(_0132_));
 CLKBUF_X3 _0670_ (.A(\uart_tx_inst.bit_cnt[0] ),
    .Z(_0133_));
 NOR4_X4 _0671_ (.A1(_0131_),
    .A2(\uart_tx_inst.bit_cnt[3] ),
    .A3(_0132_),
    .A4(_0133_),
    .ZN(_0134_));
 CLKBUF_X3 _0672_ (.A(_0134_),
    .Z(_0135_));
 MUX2_X1 _0673_ (.A(\uart_tx_inst.data_reg[1] ),
    .B(net9),
    .S(_0135_),
    .Z(_0136_));
 NOR2_X1 _0674_ (.A1(\uart_tx_inst.prescale_reg[10] ),
    .A2(\uart_tx_inst.prescale_reg[9] ),
    .ZN(_0137_));
 CLKBUF_X2 _0675_ (.A(\uart_tx_inst.prescale_reg[6] ),
    .Z(_0138_));
 NOR3_X2 _0676_ (.A1(\uart_tx_inst.prescale_reg[8] ),
    .A2(\uart_tx_inst.prescale_reg[7] ),
    .A3(_0138_),
    .ZN(_0139_));
 BUF_X2 _0677_ (.A(\uart_tx_inst.prescale_reg[2] ),
    .Z(_0140_));
 NOR4_X2 _0678_ (.A1(\uart_tx_inst.prescale_reg[3] ),
    .A2(\uart_tx_inst.prescale_reg[1] ),
    .A3(_0140_),
    .A4(\uart_tx_inst.prescale_reg[0] ),
    .ZN(_0141_));
 BUF_X2 _0679_ (.A(\uart_tx_inst.prescale_reg[4] ),
    .Z(_0142_));
 NOR2_X1 _0680_ (.A1(\uart_tx_inst.prescale_reg[5] ),
    .A2(_0142_),
    .ZN(_0143_));
 AND4_X2 _0681_ (.A1(_0137_),
    .A2(_0139_),
    .A3(_0141_),
    .A4(_0143_),
    .ZN(_0144_));
 OR3_X2 _0682_ (.A1(\uart_tx_inst.prescale_reg[13] ),
    .A2(\uart_tx_inst.prescale_reg[12] ),
    .A3(\uart_tx_inst.prescale_reg[11] ),
    .ZN(_0145_));
 NOR3_X4 _0683_ (.A1(\uart_tx_inst.prescale_reg[15] ),
    .A2(\uart_tx_inst.prescale_reg[14] ),
    .A3(_0145_),
    .ZN(_0146_));
 INV_X1 _0684_ (.A(net17),
    .ZN(_0147_));
 NAND2_X4 _0685_ (.A1(_0147_),
    .A2(_0134_),
    .ZN(_0148_));
 OR2_X1 _0686_ (.A1(\uart_tx_inst.prescale_reg[17] ),
    .A2(\uart_tx_inst.prescale_reg[16] ),
    .ZN(_0149_));
 NOR2_X2 _0687_ (.A1(\uart_tx_inst.prescale_reg[18] ),
    .A2(_0149_),
    .ZN(_0150_));
 NAND4_X4 _0688_ (.A1(_0144_),
    .A2(_0146_),
    .A3(_0148_),
    .A4(_0150_),
    .ZN(_0151_));
 NOR3_X4 _0689_ (.A1(_0131_),
    .A2(\uart_tx_inst.bit_cnt[3] ),
    .A3(_0132_),
    .ZN(_0152_));
 AND2_X2 _0690_ (.A1(_0133_),
    .A2(_0152_),
    .ZN(_0153_));
 BUF_X4 _0691_ (.A(_0153_),
    .Z(_0154_));
 NOR3_X4 _0692_ (.A1(_0082_),
    .A2(_0151_),
    .A3(_0154_),
    .ZN(_0155_));
 MUX2_X1 _0693_ (.A(\uart_tx_inst.data_reg[0] ),
    .B(_0136_),
    .S(_0155_),
    .Z(_0051_));
 MUX2_X1 _0694_ (.A(\uart_tx_inst.data_reg[2] ),
    .B(net10),
    .S(_0135_),
    .Z(_0156_));
 MUX2_X1 _0695_ (.A(\uart_tx_inst.data_reg[1] ),
    .B(_0156_),
    .S(_0155_),
    .Z(_0052_));
 MUX2_X1 _0696_ (.A(\uart_tx_inst.data_reg[3] ),
    .B(net11),
    .S(_0135_),
    .Z(_0157_));
 MUX2_X1 _0697_ (.A(\uart_tx_inst.data_reg[2] ),
    .B(_0157_),
    .S(_0155_),
    .Z(_0053_));
 MUX2_X1 _0698_ (.A(\uart_tx_inst.data_reg[4] ),
    .B(net12),
    .S(_0135_),
    .Z(_0158_));
 MUX2_X1 _0699_ (.A(\uart_tx_inst.data_reg[3] ),
    .B(_0158_),
    .S(_0155_),
    .Z(_0054_));
 MUX2_X1 _0700_ (.A(\uart_tx_inst.data_reg[5] ),
    .B(net13),
    .S(_0135_),
    .Z(_0159_));
 MUX2_X1 _0701_ (.A(\uart_tx_inst.data_reg[4] ),
    .B(_0159_),
    .S(_0155_),
    .Z(_0055_));
 MUX2_X1 _0702_ (.A(\uart_tx_inst.data_reg[6] ),
    .B(net14),
    .S(_0135_),
    .Z(_0160_));
 MUX2_X1 _0703_ (.A(\uart_tx_inst.data_reg[5] ),
    .B(_0160_),
    .S(_0155_),
    .Z(_0056_));
 MUX2_X1 _0704_ (.A(\uart_tx_inst.data_reg[7] ),
    .B(net15),
    .S(_0134_),
    .Z(_0161_));
 MUX2_X1 _0705_ (.A(\uart_tx_inst.data_reg[6] ),
    .B(_0161_),
    .S(_0155_),
    .Z(_0057_));
 MUX2_X1 _0706_ (.A(\uart_tx_inst.data_reg[8] ),
    .B(net16),
    .S(_0134_),
    .Z(_0162_));
 MUX2_X1 _0707_ (.A(\uart_tx_inst.data_reg[7] ),
    .B(_0162_),
    .S(_0155_),
    .Z(_0058_));
 AND3_X1 _0708_ (.A1(_0144_),
    .A2(_0146_),
    .A3(_0150_),
    .ZN(_0163_));
 CLKBUF_X3 _0709_ (.A(_0163_),
    .Z(_0164_));
 NAND2_X1 _0710_ (.A1(_0083_),
    .A2(_0164_),
    .ZN(_0165_));
 OAI21_X1 _0711_ (.A(\uart_tx_inst.data_reg[8] ),
    .B1(_0152_),
    .B2(_0165_),
    .ZN(_0166_));
 NAND2_X1 _0712_ (.A1(net17),
    .A2(_0135_),
    .ZN(_0167_));
 OAI21_X1 _0713_ (.A(_0166_),
    .B1(_0167_),
    .B2(_0165_),
    .ZN(_0059_));
 CLKBUF_X3 _0714_ (.A(_0083_),
    .Z(_0168_));
 INV_X1 _0715_ (.A(\uart_rx_inst.bit_cnt[3] ),
    .ZN(_0169_));
 OR2_X1 _0716_ (.A1(_0600_),
    .A2(_0085_),
    .ZN(_0170_));
 INV_X1 _0717_ (.A(_0084_),
    .ZN(_0171_));
 AOI211_X2 _0718_ (.A(_0169_),
    .B(_0127_),
    .C1(_0170_),
    .C2(_0171_),
    .ZN(_0172_));
 OR2_X2 _0719_ (.A1(_0128_),
    .A2(_0172_),
    .ZN(_0173_));
 NOR2_X1 _0720_ (.A1(\uart_rx_inst.bit_cnt[0] ),
    .A2(_0173_),
    .ZN(_0174_));
 OR2_X2 _0721_ (.A1(\uart_rx_inst.bit_cnt[1] ),
    .A2(_0091_),
    .ZN(_0175_));
 NOR2_X1 _0722_ (.A1(_0085_),
    .A2(_0175_),
    .ZN(_0176_));
 OAI21_X1 _0723_ (.A(_0088_),
    .B1(_0092_),
    .B2(_0176_),
    .ZN(_0177_));
 NAND2_X1 _0724_ (.A1(_0107_),
    .A2(_0177_),
    .ZN(_0178_));
 MUX2_X1 _0725_ (.A(_0174_),
    .B(\uart_rx_inst.bit_cnt[0] ),
    .S(_0178_),
    .Z(_0179_));
 AND2_X1 _0726_ (.A1(_0168_),
    .A2(_0179_),
    .ZN(_0002_));
 OAI21_X1 _0727_ (.A(_0112_),
    .B1(_0172_),
    .B2(_0599_),
    .ZN(_0180_));
 MUX2_X1 _0728_ (.A(_0180_),
    .B(\uart_rx_inst.bit_cnt[1] ),
    .S(_0178_),
    .Z(_0181_));
 AND2_X1 _0729_ (.A1(_0168_),
    .A2(_0181_),
    .ZN(_0003_));
 CLKBUF_X3 _0730_ (.A(_0082_),
    .Z(_0182_));
 OR2_X1 _0731_ (.A1(_0101_),
    .A2(_0106_),
    .ZN(_0183_));
 BUF_X4 _0732_ (.A(_0183_),
    .Z(_0184_));
 CLKBUF_X3 _0733_ (.A(_0184_),
    .Z(_0185_));
 NOR2_X1 _0734_ (.A1(_0600_),
    .A2(_0172_),
    .ZN(_0186_));
 OAI21_X1 _0735_ (.A(_0084_),
    .B1(_0185_),
    .B2(_0186_),
    .ZN(_0187_));
 NAND2_X1 _0736_ (.A1(_0600_),
    .A2(_0112_),
    .ZN(_0188_));
 OR3_X1 _0737_ (.A1(_0084_),
    .A2(_0178_),
    .A3(_0188_),
    .ZN(_0189_));
 AOI21_X1 _0738_ (.A(_0182_),
    .B1(_0187_),
    .B2(_0189_),
    .ZN(_0004_));
 NOR3_X1 _0739_ (.A1(_0084_),
    .A2(\uart_rx_inst.bit_cnt[1] ),
    .A3(\uart_rx_inst.bit_cnt[0] ),
    .ZN(_0190_));
 XOR2_X1 _0740_ (.A(_0001_),
    .B(_0190_),
    .Z(_0191_));
 OAI21_X1 _0741_ (.A(_0112_),
    .B1(_0172_),
    .B2(_0191_),
    .ZN(_0192_));
 MUX2_X1 _0742_ (.A(_0192_),
    .B(\uart_rx_inst.bit_cnt[3] ),
    .S(_0178_),
    .Z(_0193_));
 AND2_X1 _0743_ (.A1(_0168_),
    .A2(_0193_),
    .ZN(_0005_));
 NOR2_X2 _0744_ (.A1(_0184_),
    .A2(_0111_),
    .ZN(_0194_));
 MUX2_X1 _0745_ (.A(net27),
    .B(_0089_),
    .S(_0194_),
    .Z(_0195_));
 AND2_X1 _0746_ (.A1(_0168_),
    .A2(_0195_),
    .ZN(_0006_));
 INV_X1 _0747_ (.A(_0088_),
    .ZN(_0196_));
 NOR2_X4 _0748_ (.A1(_0196_),
    .A2(_0175_),
    .ZN(_0197_));
 NAND3_X1 _0749_ (.A1(_0089_),
    .A2(_0085_),
    .A3(_0197_),
    .ZN(_0198_));
 NOR3_X1 _0750_ (.A1(_0182_),
    .A2(_0185_),
    .A3(_0198_),
    .ZN(_0015_));
 AND3_X1 _0751_ (.A1(_0090_),
    .A2(\uart_rx_inst.bit_cnt[0] ),
    .A3(_0001_),
    .ZN(_0199_));
 NAND3_X4 _0752_ (.A1(_0107_),
    .A2(_0197_),
    .A3(_0199_),
    .ZN(_0200_));
 NAND2_X1 _0753_ (.A1(net18),
    .A2(_0200_),
    .ZN(_0201_));
 AND3_X1 _0754_ (.A1(_0107_),
    .A2(_0197_),
    .A3(_0199_),
    .ZN(_0202_));
 BUF_X2 _0755_ (.A(_0202_),
    .Z(_0203_));
 NAND2_X1 _0756_ (.A1(\uart_rx_inst.data_reg[0] ),
    .A2(_0203_),
    .ZN(_0204_));
 AOI21_X1 _0757_ (.A(_0182_),
    .B1(_0201_),
    .B2(_0204_),
    .ZN(_0016_));
 NAND2_X1 _0758_ (.A1(net19),
    .A2(_0200_),
    .ZN(_0205_));
 NAND2_X1 _0759_ (.A1(\uart_rx_inst.data_reg[1] ),
    .A2(_0203_),
    .ZN(_0206_));
 AOI21_X1 _0760_ (.A(_0182_),
    .B1(_0205_),
    .B2(_0206_),
    .ZN(_0017_));
 NAND2_X1 _0761_ (.A1(net20),
    .A2(_0200_),
    .ZN(_0207_));
 NAND2_X1 _0762_ (.A1(\uart_rx_inst.data_reg[2] ),
    .A2(_0203_),
    .ZN(_0208_));
 AOI21_X1 _0763_ (.A(_0182_),
    .B1(_0207_),
    .B2(_0208_),
    .ZN(_0018_));
 CLKBUF_X3 _0764_ (.A(_0082_),
    .Z(_0209_));
 NAND2_X1 _0765_ (.A1(net21),
    .A2(_0200_),
    .ZN(_0210_));
 NAND2_X1 _0766_ (.A1(\uart_rx_inst.data_reg[3] ),
    .A2(_0203_),
    .ZN(_0211_));
 AOI21_X1 _0767_ (.A(_0209_),
    .B1(_0210_),
    .B2(_0211_),
    .ZN(_0019_));
 NAND2_X1 _0768_ (.A1(net22),
    .A2(_0200_),
    .ZN(_0212_));
 NAND2_X1 _0769_ (.A1(\uart_rx_inst.data_reg[4] ),
    .A2(_0203_),
    .ZN(_0213_));
 AOI21_X1 _0770_ (.A(_0209_),
    .B1(_0212_),
    .B2(_0213_),
    .ZN(_0020_));
 NAND2_X1 _0771_ (.A1(net23),
    .A2(_0200_),
    .ZN(_0214_));
 NAND2_X1 _0772_ (.A1(\uart_rx_inst.data_reg[5] ),
    .A2(_0203_),
    .ZN(_0215_));
 AOI21_X1 _0773_ (.A(_0209_),
    .B1(_0214_),
    .B2(_0215_),
    .ZN(_0021_));
 NAND2_X1 _0774_ (.A1(net24),
    .A2(_0200_),
    .ZN(_0216_));
 NAND2_X1 _0775_ (.A1(\uart_rx_inst.data_reg[6] ),
    .A2(_0203_),
    .ZN(_0217_));
 AOI21_X1 _0776_ (.A(_0209_),
    .B1(_0216_),
    .B2(_0217_),
    .ZN(_0022_));
 NAND2_X1 _0777_ (.A1(net25),
    .A2(_0200_),
    .ZN(_0218_));
 NAND2_X1 _0778_ (.A1(\uart_rx_inst.data_reg[7] ),
    .A2(_0203_),
    .ZN(_0219_));
 AOI21_X1 _0779_ (.A(_0209_),
    .B1(_0218_),
    .B2(_0219_),
    .ZN(_0023_));
 INV_X1 _0780_ (.A(net1),
    .ZN(_0220_));
 NAND2_X1 _0781_ (.A1(net26),
    .A2(_0220_),
    .ZN(_0221_));
 CLKBUF_X3 _0782_ (.A(_0107_),
    .Z(_0222_));
 NAND4_X1 _0783_ (.A1(\uart_rx_inst.rxd_reg ),
    .A2(_0085_),
    .A3(_0222_),
    .A4(_0197_),
    .ZN(_0223_));
 AOI21_X1 _0784_ (.A(_0209_),
    .B1(_0221_),
    .B2(_0223_),
    .ZN(_0024_));
 NAND4_X1 _0785_ (.A1(\uart_rx_inst.rxd_reg ),
    .A2(net26),
    .A3(_0085_),
    .A4(_0197_),
    .ZN(_0224_));
 NOR3_X1 _0786_ (.A1(_0182_),
    .A2(_0185_),
    .A3(_0224_),
    .ZN(_0025_));
 OAI21_X4 _0787_ (.A(_0083_),
    .B1(_0094_),
    .B2(_0184_),
    .ZN(_0225_));
 CLKBUF_X3 _0788_ (.A(_0225_),
    .Z(_0226_));
 NOR2_X4 _0789_ (.A1(_0128_),
    .A2(_0172_),
    .ZN(_0227_));
 NAND2_X1 _0790_ (.A1(_0222_),
    .A2(_0227_),
    .ZN(_0228_));
 NAND2_X1 _0791_ (.A1(_0588_),
    .A2(_0185_),
    .ZN(_0229_));
 AOI21_X1 _0792_ (.A(_0226_),
    .B1(_0228_),
    .B2(_0229_),
    .ZN(_0026_));
 BUF_X4 _0793_ (.A(prescale[8]),
    .Z(_0230_));
 CLKBUF_X2 _0794_ (.A(_0594_),
    .Z(_0231_));
 BUF_X2 _0795_ (.A(prescale[2]),
    .Z(_0232_));
 CLKBUF_X2 _0796_ (.A(prescale[3]),
    .Z(_0233_));
 NOR2_X2 _0797_ (.A1(_0232_),
    .A2(_0233_),
    .ZN(_0234_));
 BUF_X1 _0798_ (.A(prescale[4]),
    .Z(_0235_));
 BUF_X1 _0799_ (.A(prescale[5]),
    .Z(_0236_));
 NOR2_X1 _0800_ (.A1(_0235_),
    .A2(_0236_),
    .ZN(_0237_));
 CLKBUF_X3 _0801_ (.A(prescale[6]),
    .Z(_0238_));
 BUF_X2 _0802_ (.A(prescale[7]),
    .Z(_0239_));
 NOR2_X1 _0803_ (.A1(_0238_),
    .A2(_0239_),
    .ZN(_0240_));
 NAND4_X2 _0804_ (.A1(_0231_),
    .A2(_0234_),
    .A3(_0237_),
    .A4(_0240_),
    .ZN(_0241_));
 XOR2_X2 _0805_ (.A(_0230_),
    .B(_0241_),
    .Z(_0242_));
 OR2_X1 _0806_ (.A1(_0232_),
    .A2(_0233_),
    .ZN(_0243_));
 OR4_X1 _0807_ (.A1(_0081_),
    .A2(net6),
    .A3(_0235_),
    .A4(_0236_),
    .ZN(_0244_));
 NOR3_X1 _0808_ (.A1(_0238_),
    .A2(_0243_),
    .A3(_0244_),
    .ZN(_0245_));
 XNOR2_X1 _0809_ (.A(_0239_),
    .B(_0245_),
    .ZN(_0246_));
 OAI221_X1 _0810_ (.A(_0107_),
    .B1(_0112_),
    .B2(_0242_),
    .C1(_0246_),
    .C2(_0173_),
    .ZN(_0247_));
 INV_X1 _0811_ (.A(_0096_),
    .ZN(_0248_));
 BUF_X1 _0812_ (.A(_0590_),
    .Z(_0249_));
 NAND4_X1 _0813_ (.A1(_0248_),
    .A2(_0249_),
    .A3(_0095_),
    .A4(_0099_),
    .ZN(_0250_));
 OAI21_X1 _0814_ (.A(\uart_rx_inst.prescale_reg[10] ),
    .B1(_0250_),
    .B2(\uart_rx_inst.prescale_reg[9] ),
    .ZN(_0251_));
 NAND2_X1 _0815_ (.A1(_0099_),
    .A2(_0100_),
    .ZN(_0252_));
 NAND3_X2 _0816_ (.A1(_0248_),
    .A2(_0249_),
    .A3(_0095_),
    .ZN(_0253_));
 OR2_X1 _0817_ (.A1(_0252_),
    .A2(_0253_),
    .ZN(_0254_));
 NAND2_X1 _0818_ (.A1(_0251_),
    .A2(_0254_),
    .ZN(_0255_));
 OAI21_X1 _0819_ (.A(_0247_),
    .B1(_0255_),
    .B2(_0222_),
    .ZN(_0256_));
 NOR2_X1 _0820_ (.A1(_0226_),
    .A2(_0256_),
    .ZN(_0027_));
 NOR4_X1 _0821_ (.A1(\uart_rx_inst.prescale_reg[15] ),
    .A2(_0102_),
    .A3(_0104_),
    .A4(_0105_),
    .ZN(_0257_));
 OR2_X1 _0822_ (.A1(_0101_),
    .A2(_0257_),
    .ZN(_0258_));
 NOR2_X1 _0823_ (.A1(_0103_),
    .A2(_0258_),
    .ZN(_0259_));
 AOI21_X1 _0824_ (.A(_0259_),
    .B1(_0101_),
    .B2(_0103_),
    .ZN(_0260_));
 NOR2_X1 _0825_ (.A1(_0173_),
    .A2(_0242_),
    .ZN(_0261_));
 OR2_X1 _0826_ (.A1(_0243_),
    .A2(_0244_),
    .ZN(_0262_));
 BUF_X8 _0827_ (.A(_0262_),
    .Z(_0263_));
 OR3_X1 _0828_ (.A1(_0238_),
    .A2(_0239_),
    .A3(_0230_),
    .ZN(_0264_));
 NOR2_X1 _0829_ (.A1(_0263_),
    .A2(_0264_),
    .ZN(_0265_));
 XOR2_X2 _0830_ (.A(net7),
    .B(_0265_),
    .Z(_0266_));
 AOI21_X1 _0831_ (.A(_0261_),
    .B1(_0266_),
    .B2(_0129_),
    .ZN(_0267_));
 NAND2_X1 _0832_ (.A1(_0090_),
    .A2(_0091_),
    .ZN(_0268_));
 AOI21_X1 _0833_ (.A(_0196_),
    .B1(_0268_),
    .B2(_0175_),
    .ZN(_0269_));
 AOI21_X2 _0834_ (.A(_0082_),
    .B1(_0269_),
    .B2(_0107_),
    .ZN(_0270_));
 NAND2_X1 _0835_ (.A1(_0222_),
    .A2(_0270_),
    .ZN(_0271_));
 OAI22_X1 _0836_ (.A1(_0226_),
    .A2(_0260_),
    .B1(_0267_),
    .B2(_0271_),
    .ZN(_0028_));
 BUF_X2 _0837_ (.A(prescale[10]),
    .Z(_0272_));
 NAND3_X1 _0838_ (.A1(_0231_),
    .A2(_0234_),
    .A3(_0237_),
    .ZN(_0273_));
 CLKBUF_X3 _0839_ (.A(_0273_),
    .Z(_0274_));
 OR4_X2 _0840_ (.A1(_0238_),
    .A2(_0239_),
    .A3(_0230_),
    .A4(net7),
    .ZN(_0275_));
 NOR2_X1 _0841_ (.A1(_0274_),
    .A2(_0275_),
    .ZN(_0276_));
 XOR2_X2 _0842_ (.A(_0272_),
    .B(_0276_),
    .Z(_0277_));
 AOI22_X1 _0843_ (.A1(_0227_),
    .A2(_0266_),
    .B1(_0277_),
    .B2(_0129_),
    .ZN(_0278_));
 NAND2_X1 _0844_ (.A1(_0083_),
    .A2(_0184_),
    .ZN(_0279_));
 NOR2_X1 _0845_ (.A1(_0103_),
    .A2(_0254_),
    .ZN(_0280_));
 XNOR2_X1 _0846_ (.A(\uart_rx_inst.prescale_reg[12] ),
    .B(_0280_),
    .ZN(_0281_));
 OAI22_X1 _0847_ (.A1(_0271_),
    .A2(_0278_),
    .B1(_0279_),
    .B2(_0281_),
    .ZN(_0029_));
 INV_X1 _0848_ (.A(\uart_rx_inst.prescale_reg[13] ),
    .ZN(_0282_));
 NOR3_X1 _0849_ (.A1(_0103_),
    .A2(\uart_rx_inst.prescale_reg[12] ),
    .A3(_0101_),
    .ZN(_0283_));
 NOR3_X1 _0850_ (.A1(_0082_),
    .A2(_0282_),
    .A3(_0283_),
    .ZN(_0284_));
 NOR4_X1 _0851_ (.A1(_0272_),
    .A2(_0243_),
    .A3(_0244_),
    .A4(_0275_),
    .ZN(_0285_));
 XNOR2_X1 _0852_ (.A(net2),
    .B(_0285_),
    .ZN(_0286_));
 NOR3_X1 _0853_ (.A1(_0184_),
    .A2(_0113_),
    .A3(_0286_),
    .ZN(_0287_));
 AOI21_X1 _0854_ (.A(_0284_),
    .B1(_0287_),
    .B2(_0270_),
    .ZN(_0288_));
 NOR2_X1 _0855_ (.A1(_0104_),
    .A2(_0258_),
    .ZN(_0289_));
 NOR2_X1 _0856_ (.A1(_0184_),
    .A2(_0173_),
    .ZN(_0290_));
 AOI21_X1 _0857_ (.A(_0289_),
    .B1(_0277_),
    .B2(_0290_),
    .ZN(_0291_));
 OAI21_X1 _0858_ (.A(_0288_),
    .B1(_0291_),
    .B2(_0226_),
    .ZN(_0030_));
 BUF_X2 _0859_ (.A(prescale[12]),
    .Z(_0292_));
 OR3_X1 _0860_ (.A1(_0272_),
    .A2(net2),
    .A3(_0275_),
    .ZN(_0293_));
 BUF_X8 _0861_ (.A(_0293_),
    .Z(_0294_));
 NOR2_X1 _0862_ (.A1(_0273_),
    .A2(_0294_),
    .ZN(_0295_));
 XOR2_X2 _0863_ (.A(_0292_),
    .B(_0295_),
    .Z(_0296_));
 OAI21_X1 _0864_ (.A(_0129_),
    .B1(_0296_),
    .B2(_0090_),
    .ZN(_0297_));
 NOR2_X1 _0865_ (.A1(_0173_),
    .A2(_0286_),
    .ZN(_0298_));
 OR2_X1 _0866_ (.A1(_0184_),
    .A2(_0197_),
    .ZN(_0299_));
 NOR2_X1 _0867_ (.A1(_0298_),
    .A2(_0299_),
    .ZN(_0300_));
 NOR2_X1 _0868_ (.A1(_0104_),
    .A2(_0254_),
    .ZN(_0301_));
 XNOR2_X1 _0869_ (.A(_0102_),
    .B(_0301_),
    .ZN(_0302_));
 AOI221_X1 _0870_ (.A(_0225_),
    .B1(_0297_),
    .B2(_0300_),
    .C1(_0302_),
    .C2(_0185_),
    .ZN(_0031_));
 INV_X1 _0871_ (.A(\uart_rx_inst.prescale_reg[15] ),
    .ZN(_0303_));
 AND2_X1 _0872_ (.A1(_0303_),
    .A2(_0105_),
    .ZN(_0304_));
 NOR3_X1 _0873_ (.A1(_0102_),
    .A2(_0101_),
    .A3(_0104_),
    .ZN(_0305_));
 MUX2_X1 _0874_ (.A(\uart_rx_inst.prescale_reg[15] ),
    .B(_0304_),
    .S(_0305_),
    .Z(_0306_));
 NOR3_X1 _0875_ (.A1(_0292_),
    .A2(_0263_),
    .A3(_0294_),
    .ZN(_0307_));
 XOR2_X2 _0876_ (.A(net3),
    .B(_0307_),
    .Z(_0308_));
 AOI221_X2 _0877_ (.A(_0306_),
    .B1(_0308_),
    .B2(_0194_),
    .C1(_0290_),
    .C2(_0296_),
    .ZN(_0309_));
 NOR2_X1 _0878_ (.A1(_0226_),
    .A2(_0309_),
    .ZN(_0032_));
 AOI21_X1 _0879_ (.A(_0299_),
    .B1(_0308_),
    .B2(_0227_),
    .ZN(_0310_));
 OR2_X1 _0880_ (.A1(_0292_),
    .A2(net3),
    .ZN(_0311_));
 OR3_X1 _0881_ (.A1(_0273_),
    .A2(_0294_),
    .A3(_0311_),
    .ZN(_0312_));
 XNOR2_X2 _0882_ (.A(net4),
    .B(_0312_),
    .ZN(_0313_));
 OAI21_X1 _0883_ (.A(_0129_),
    .B1(_0313_),
    .B2(_0090_),
    .ZN(_0314_));
 OR3_X1 _0884_ (.A1(\uart_rx_inst.prescale_reg[15] ),
    .A2(_0102_),
    .A3(_0104_),
    .ZN(_0315_));
 NOR2_X1 _0885_ (.A1(_0254_),
    .A2(_0315_),
    .ZN(_0316_));
 XNOR2_X1 _0886_ (.A(\uart_rx_inst.prescale_reg[16] ),
    .B(_0316_),
    .ZN(_0317_));
 AOI221_X1 _0887_ (.A(_0225_),
    .B1(_0310_),
    .B2(_0314_),
    .C1(_0317_),
    .C2(_0184_),
    .ZN(_0033_));
 NOR3_X1 _0888_ (.A1(\uart_rx_inst.prescale_reg[16] ),
    .A2(_0101_),
    .A3(_0315_),
    .ZN(_0318_));
 XNOR2_X1 _0889_ (.A(\uart_rx_inst.prescale_reg[17] ),
    .B(_0318_),
    .ZN(_0319_));
 OR2_X1 _0890_ (.A1(net4),
    .A2(_0311_),
    .ZN(_0320_));
 NOR3_X2 _0891_ (.A1(_0263_),
    .A2(_0294_),
    .A3(_0320_),
    .ZN(_0321_));
 XOR2_X2 _0892_ (.A(net5),
    .B(_0321_),
    .Z(_0322_));
 AOI221_X2 _0893_ (.A(_0184_),
    .B1(_0227_),
    .B2(_0313_),
    .C1(_0322_),
    .C2(_0129_),
    .ZN(_0323_));
 NOR3_X1 _0894_ (.A1(_0226_),
    .A2(_0319_),
    .A3(_0323_),
    .ZN(_0034_));
 OR4_X1 _0895_ (.A1(net5),
    .A2(_0274_),
    .A3(_0294_),
    .A4(_0320_),
    .ZN(_0324_));
 AOI21_X1 _0896_ (.A(_0112_),
    .B1(_0324_),
    .B2(_0089_),
    .ZN(_0325_));
 AOI21_X1 _0897_ (.A(_0325_),
    .B1(_0322_),
    .B2(_0227_),
    .ZN(_0326_));
 OR4_X1 _0898_ (.A1(\uart_rx_inst.prescale_reg[17] ),
    .A2(\uart_rx_inst.prescale_reg[16] ),
    .A3(_0252_),
    .A4(_0315_),
    .ZN(_0327_));
 NAND2_X1 _0899_ (.A1(_0095_),
    .A2(_0097_),
    .ZN(_0328_));
 AOI21_X1 _0900_ (.A(_0327_),
    .B1(_0253_),
    .B2(_0328_),
    .ZN(_0329_));
 NOR2_X1 _0901_ (.A1(\uart_rx_inst.prescale_reg[18] ),
    .A2(_0329_),
    .ZN(_0330_));
 INV_X1 _0902_ (.A(\uart_rx_inst.prescale_reg[18] ),
    .ZN(_0331_));
 NOR3_X1 _0903_ (.A1(_0331_),
    .A2(_0253_),
    .A3(_0327_),
    .ZN(_0332_));
 OAI33_X1 _0904_ (.A1(_0185_),
    .A2(_0225_),
    .A3(_0326_),
    .B1(_0330_),
    .B2(_0332_),
    .B3(_0279_),
    .ZN(_0035_));
 MUX2_X1 _0905_ (.A(_0591_),
    .B(_0172_),
    .S(_0107_),
    .Z(_0333_));
 NOR2_X1 _0906_ (.A1(_0226_),
    .A2(_0333_),
    .ZN(_0036_));
 AOI21_X1 _0907_ (.A(_0172_),
    .B1(_0129_),
    .B2(_0081_),
    .ZN(_0334_));
 NOR2_X1 _0908_ (.A1(_0185_),
    .A2(_0334_),
    .ZN(_0335_));
 XOR2_X1 _0909_ (.A(_0096_),
    .B(_0249_),
    .Z(_0336_));
 NOR2_X1 _0910_ (.A1(_0222_),
    .A2(_0336_),
    .ZN(_0337_));
 NOR3_X1 _0911_ (.A1(_0226_),
    .A2(_0335_),
    .A3(_0337_),
    .ZN(_0037_));
 NOR2_X1 _0912_ (.A1(_0595_),
    .A2(_0112_),
    .ZN(_0338_));
 NOR3_X1 _0913_ (.A1(_0081_),
    .A2(_0129_),
    .A3(_0172_),
    .ZN(_0339_));
 NOR3_X1 _0914_ (.A1(_0185_),
    .A2(_0338_),
    .A3(_0339_),
    .ZN(_0340_));
 XNOR2_X1 _0915_ (.A(\uart_rx_inst.prescale_reg[3] ),
    .B(_0097_),
    .ZN(_0341_));
 NOR3_X1 _0916_ (.A1(_0226_),
    .A2(_0340_),
    .A3(_0341_),
    .ZN(_0038_));
 XNOR2_X1 _0917_ (.A(_0232_),
    .B(_0231_),
    .ZN(_0342_));
 NOR2_X1 _0918_ (.A1(_0089_),
    .A2(_0087_),
    .ZN(_0343_));
 OR2_X1 _0919_ (.A1(_0595_),
    .A2(_0128_),
    .ZN(_0344_));
 OAI221_X1 _0920_ (.A(_0222_),
    .B1(_0113_),
    .B2(_0342_),
    .C1(_0343_),
    .C2(_0344_),
    .ZN(_0345_));
 NAND2_X1 _0921_ (.A1(_0248_),
    .A2(_0249_),
    .ZN(_0346_));
 OAI21_X1 _0922_ (.A(\uart_rx_inst.prescale_reg[4] ),
    .B1(\uart_rx_inst.prescale_reg[3] ),
    .B2(_0346_),
    .ZN(_0347_));
 NAND3_X1 _0923_ (.A1(_0185_),
    .A2(_0253_),
    .A3(_0347_),
    .ZN(_0348_));
 AND3_X1 _0924_ (.A1(_0270_),
    .A2(_0345_),
    .A3(_0348_),
    .ZN(_0039_));
 XNOR2_X1 _0925_ (.A(_0098_),
    .B(_0328_),
    .ZN(_0349_));
 NAND2_X1 _0926_ (.A1(_0299_),
    .A2(_0349_),
    .ZN(_0350_));
 OAI21_X1 _0927_ (.A(_0113_),
    .B1(_0342_),
    .B2(_0343_),
    .ZN(_0351_));
 NOR3_X2 _0928_ (.A1(_0081_),
    .A2(_0232_),
    .A3(net6),
    .ZN(_0352_));
 XNOR2_X1 _0929_ (.A(_0233_),
    .B(_0352_),
    .ZN(_0353_));
 NAND3_X1 _0930_ (.A1(_0089_),
    .A2(_0129_),
    .A3(_0353_),
    .ZN(_0354_));
 NAND3_X1 _0931_ (.A1(_0222_),
    .A2(_0351_),
    .A3(_0354_),
    .ZN(_0355_));
 AOI21_X1 _0932_ (.A(_0225_),
    .B1(_0350_),
    .B2(_0355_),
    .ZN(_0040_));
 INV_X1 _0933_ (.A(_0299_),
    .ZN(_0356_));
 OAI21_X1 _0934_ (.A(_0111_),
    .B1(_0343_),
    .B2(_0353_),
    .ZN(_0357_));
 NAND2_X1 _0935_ (.A1(_0231_),
    .A2(_0234_),
    .ZN(_0358_));
 XNOR2_X1 _0936_ (.A(_0235_),
    .B(_0358_),
    .ZN(_0359_));
 NAND2_X1 _0937_ (.A1(_0089_),
    .A2(_0128_),
    .ZN(_0360_));
 OAI21_X1 _0938_ (.A(_0357_),
    .B1(_0359_),
    .B2(_0360_),
    .ZN(_0361_));
 NOR2_X1 _0939_ (.A1(_0098_),
    .A2(_0253_),
    .ZN(_0362_));
 XNOR2_X1 _0940_ (.A(\uart_rx_inst.prescale_reg[6] ),
    .B(_0362_),
    .ZN(_0363_));
 AOI221_X1 _0941_ (.A(_0225_),
    .B1(_0356_),
    .B2(_0361_),
    .C1(_0363_),
    .C2(_0184_),
    .ZN(_0041_));
 NOR3_X1 _0942_ (.A1(\uart_rx_inst.prescale_reg[6] ),
    .A2(_0098_),
    .A3(_0328_),
    .ZN(_0364_));
 XOR2_X1 _0943_ (.A(\uart_rx_inst.prescale_reg[7] ),
    .B(_0364_),
    .Z(_0365_));
 NAND2_X1 _0944_ (.A1(_0270_),
    .A2(_0365_),
    .ZN(_0366_));
 NOR2_X1 _0945_ (.A1(_0233_),
    .A2(_0235_),
    .ZN(_0367_));
 NAND2_X1 _0946_ (.A1(_0352_),
    .A2(_0367_),
    .ZN(_0368_));
 XOR2_X1 _0947_ (.A(_0236_),
    .B(_0368_),
    .Z(_0369_));
 OAI21_X1 _0948_ (.A(_0359_),
    .B1(_0087_),
    .B2(_0089_),
    .ZN(_0370_));
 MUX2_X1 _0949_ (.A(_0369_),
    .B(_0370_),
    .S(_0112_),
    .Z(_0371_));
 AOI21_X1 _0950_ (.A(_0366_),
    .B1(_0371_),
    .B2(_0222_),
    .ZN(_0042_));
 INV_X1 _0951_ (.A(_0238_),
    .ZN(_0372_));
 XNOR2_X1 _0952_ (.A(_0372_),
    .B(_0274_),
    .ZN(_0373_));
 OAI221_X1 _0953_ (.A(_0107_),
    .B1(_0173_),
    .B2(_0369_),
    .C1(_0373_),
    .C2(_0112_),
    .ZN(_0374_));
 OR4_X1 _0954_ (.A1(\uart_rx_inst.prescale_reg[7] ),
    .A2(\uart_rx_inst.prescale_reg[6] ),
    .A3(_0098_),
    .A4(_0253_),
    .ZN(_0375_));
 XNOR2_X1 _0955_ (.A(\uart_rx_inst.prescale_reg[8] ),
    .B(_0375_),
    .ZN(_0376_));
 OAI21_X1 _0956_ (.A(_0374_),
    .B1(_0376_),
    .B2(_0222_),
    .ZN(_0377_));
 NOR2_X1 _0957_ (.A1(_0226_),
    .A2(_0377_),
    .ZN(_0043_));
 NAND3_X1 _0958_ (.A1(_0238_),
    .A2(_0227_),
    .A3(_0274_),
    .ZN(_0378_));
 AND2_X1 _0959_ (.A1(_0239_),
    .A2(_0128_),
    .ZN(_0379_));
 OAI21_X1 _0960_ (.A(_0379_),
    .B1(_0263_),
    .B2(_0238_),
    .ZN(_0380_));
 NOR3_X1 _0961_ (.A1(_0129_),
    .A2(_0172_),
    .A3(_0274_),
    .ZN(_0381_));
 NOR3_X1 _0962_ (.A1(_0239_),
    .A2(_0112_),
    .A3(_0263_),
    .ZN(_0382_));
 OAI21_X1 _0963_ (.A(_0372_),
    .B1(_0381_),
    .B2(_0382_),
    .ZN(_0383_));
 NAND4_X1 _0964_ (.A1(_0222_),
    .A2(_0378_),
    .A3(_0380_),
    .A4(_0383_),
    .ZN(_0384_));
 NOR2_X1 _0965_ (.A1(_0096_),
    .A2(\uart_rx_inst.prescale_reg[1] ),
    .ZN(_0385_));
 NAND4_X1 _0966_ (.A1(_0588_),
    .A2(_0095_),
    .A3(_0385_),
    .A4(_0099_),
    .ZN(_0386_));
 XOR2_X1 _0967_ (.A(\uart_rx_inst.prescale_reg[9] ),
    .B(_0386_),
    .Z(_0387_));
 AOI21_X1 _0968_ (.A(_0225_),
    .B1(_0387_),
    .B2(_0185_),
    .ZN(_0388_));
 AND2_X1 _0969_ (.A1(_0384_),
    .A2(_0388_),
    .ZN(_0044_));
 OR2_X1 _0970_ (.A1(_0209_),
    .A2(net8),
    .ZN(_0045_));
 AND2_X1 _0971_ (.A1(_0147_),
    .A2(_0134_),
    .ZN(_0389_));
 NAND3_X2 _0972_ (.A1(_0144_),
    .A2(_0146_),
    .A3(_0150_),
    .ZN(_0390_));
 BUF_X4 _0973_ (.A(_0390_),
    .Z(_0391_));
 NOR3_X1 _0974_ (.A1(_0133_),
    .A2(_0389_),
    .A3(_0391_),
    .ZN(_0392_));
 CLKBUF_X3 _0975_ (.A(_0391_),
    .Z(_0393_));
 AOI21_X1 _0976_ (.A(_0392_),
    .B1(_0393_),
    .B2(_0133_),
    .ZN(_0394_));
 NOR2_X1 _0977_ (.A1(_0182_),
    .A2(_0394_),
    .ZN(_0046_));
 OAI21_X1 _0978_ (.A(_0168_),
    .B1(_0393_),
    .B2(_0167_),
    .ZN(_0395_));
 NOR2_X1 _0979_ (.A1(_0133_),
    .A2(_0151_),
    .ZN(_0396_));
 XNOR2_X1 _0980_ (.A(_0132_),
    .B(_0396_),
    .ZN(_0397_));
 NOR2_X1 _0981_ (.A1(_0395_),
    .A2(_0397_),
    .ZN(_0047_));
 NOR3_X1 _0982_ (.A1(_0132_),
    .A2(_0133_),
    .A3(_0151_),
    .ZN(_0398_));
 XNOR2_X1 _0983_ (.A(_0131_),
    .B(_0398_),
    .ZN(_0399_));
 NOR2_X1 _0984_ (.A1(_0395_),
    .A2(_0399_),
    .ZN(_0048_));
 NOR4_X1 _0985_ (.A1(_0131_),
    .A2(_0132_),
    .A3(_0133_),
    .A4(_0391_),
    .ZN(_0400_));
 INV_X1 _0986_ (.A(\uart_tx_inst.bit_cnt[3] ),
    .ZN(_0401_));
 OAI22_X1 _0987_ (.A1(_0393_),
    .A2(_0167_),
    .B1(_0400_),
    .B2(_0401_),
    .ZN(_0402_));
 AND2_X1 _0988_ (.A1(_0168_),
    .A2(_0402_),
    .ZN(_0049_));
 OAI21_X4 _0989_ (.A(_0083_),
    .B1(_0148_),
    .B2(_0390_),
    .ZN(_0403_));
 AOI21_X1 _0990_ (.A(net31),
    .B1(_0135_),
    .B2(_0164_),
    .ZN(_0404_));
 NOR2_X1 _0991_ (.A1(_0403_),
    .A2(_0404_),
    .ZN(_0050_));
 NOR2_X1 _0992_ (.A1(_0604_),
    .A2(_0164_),
    .ZN(_0405_));
 NAND2_X2 _0993_ (.A1(_0133_),
    .A2(_0152_),
    .ZN(_0406_));
 NOR2_X1 _0994_ (.A1(_0406_),
    .A2(_0393_),
    .ZN(_0407_));
 NOR3_X1 _0995_ (.A1(_0403_),
    .A2(_0405_),
    .A3(_0407_),
    .ZN(_0060_));
 OR2_X1 _0996_ (.A1(\uart_tx_inst.prescale_reg[7] ),
    .A2(_0138_),
    .ZN(_0408_));
 BUF_X1 _0997_ (.A(_0606_),
    .Z(_0409_));
 NOR4_X4 _0998_ (.A1(\uart_tx_inst.prescale_reg[5] ),
    .A2(_0142_),
    .A3(\uart_tx_inst.prescale_reg[3] ),
    .A4(_0140_),
    .ZN(_0410_));
 NAND2_X1 _0999_ (.A1(_0409_),
    .A2(_0410_),
    .ZN(_0411_));
 OR4_X1 _1000_ (.A1(\uart_tx_inst.prescale_reg[9] ),
    .A2(\uart_tx_inst.prescale_reg[8] ),
    .A3(_0408_),
    .A4(_0411_),
    .ZN(_0412_));
 MUX2_X1 _1001_ (.A(_0389_),
    .B(_0412_),
    .S(_0391_),
    .Z(_0413_));
 AOI21_X1 _1002_ (.A(_0412_),
    .B1(_0164_),
    .B2(_0389_),
    .ZN(_0414_));
 MUX2_X1 _1003_ (.A(_0413_),
    .B(_0414_),
    .S(\uart_tx_inst.prescale_reg[10] ),
    .Z(_0415_));
 NOR3_X1 _1004_ (.A1(_0238_),
    .A2(_0154_),
    .A3(_0263_),
    .ZN(_0416_));
 XOR2_X1 _1005_ (.A(_0239_),
    .B(_0416_),
    .Z(_0417_));
 OAI21_X1 _1006_ (.A(_0168_),
    .B1(_0151_),
    .B2(_0417_),
    .ZN(_0418_));
 NOR2_X1 _1007_ (.A1(_0415_),
    .A2(_0418_),
    .ZN(_0061_));
 NOR4_X1 _1008_ (.A1(_0238_),
    .A2(_0239_),
    .A3(_0153_),
    .A4(_0274_),
    .ZN(_0419_));
 XOR2_X1 _1009_ (.A(_0230_),
    .B(_0419_),
    .Z(_0420_));
 OAI21_X1 _1010_ (.A(_0168_),
    .B1(_0151_),
    .B2(_0420_),
    .ZN(_0421_));
 OAI21_X1 _1011_ (.A(_0144_),
    .B1(_0148_),
    .B2(_0391_),
    .ZN(_0422_));
 XOR2_X1 _1012_ (.A(\uart_tx_inst.prescale_reg[11] ),
    .B(_0422_),
    .Z(_0423_));
 NOR2_X1 _1013_ (.A1(_0421_),
    .A2(_0423_),
    .ZN(_0062_));
 NAND4_X2 _1014_ (.A1(_0409_),
    .A2(_0137_),
    .A3(_0139_),
    .A4(_0410_),
    .ZN(_0424_));
 NOR2_X1 _1015_ (.A1(\uart_tx_inst.prescale_reg[11] ),
    .A2(_0424_),
    .ZN(_0425_));
 NAND2_X1 _1016_ (.A1(\uart_tx_inst.prescale_reg[12] ),
    .A2(_0425_),
    .ZN(_0426_));
 MUX2_X1 _1017_ (.A(_0148_),
    .B(_0425_),
    .S(_0391_),
    .Z(_0427_));
 OAI21_X1 _1018_ (.A(_0426_),
    .B1(_0427_),
    .B2(\uart_tx_inst.prescale_reg[12] ),
    .ZN(_0428_));
 OR3_X1 _1019_ (.A1(_0153_),
    .A2(_0263_),
    .A3(_0264_),
    .ZN(_0429_));
 XNOR2_X1 _1020_ (.A(net7),
    .B(_0429_),
    .ZN(_0430_));
 OAI21_X1 _1021_ (.A(_0168_),
    .B1(_0151_),
    .B2(_0430_),
    .ZN(_0431_));
 NOR2_X1 _1022_ (.A1(_0428_),
    .A2(_0431_),
    .ZN(_0063_));
 NOR3_X1 _1023_ (.A1(_0154_),
    .A2(_0274_),
    .A3(_0275_),
    .ZN(_0432_));
 XOR2_X1 _1024_ (.A(_0272_),
    .B(_0432_),
    .Z(_0433_));
 AOI21_X1 _1025_ (.A(_0393_),
    .B1(_0433_),
    .B2(_0148_),
    .ZN(_0434_));
 NOR2_X1 _1026_ (.A1(\uart_tx_inst.prescale_reg[12] ),
    .A2(\uart_tx_inst.prescale_reg[11] ),
    .ZN(_0435_));
 NAND2_X1 _1027_ (.A1(_0144_),
    .A2(_0435_),
    .ZN(_0436_));
 XOR2_X1 _1028_ (.A(\uart_tx_inst.prescale_reg[13] ),
    .B(_0436_),
    .Z(_0437_));
 NOR3_X1 _1029_ (.A1(_0182_),
    .A2(_0434_),
    .A3(_0437_),
    .ZN(_0064_));
 NOR4_X1 _1030_ (.A1(_0272_),
    .A2(_0153_),
    .A3(_0263_),
    .A4(_0275_),
    .ZN(_0438_));
 XNOR2_X1 _1031_ (.A(net2),
    .B(_0438_),
    .ZN(_0439_));
 NOR2_X1 _1032_ (.A1(_0145_),
    .A2(_0424_),
    .ZN(_0440_));
 XNOR2_X1 _1033_ (.A(\uart_tx_inst.prescale_reg[14] ),
    .B(_0440_),
    .ZN(_0441_));
 MUX2_X1 _1034_ (.A(_0439_),
    .B(_0441_),
    .S(_0391_),
    .Z(_0442_));
 NOR2_X1 _1035_ (.A1(_0403_),
    .A2(_0442_),
    .ZN(_0065_));
 OR2_X1 _1036_ (.A1(\uart_tx_inst.prescale_reg[14] ),
    .A2(\uart_tx_inst.prescale_reg[13] ),
    .ZN(_0443_));
 OAI21_X1 _1037_ (.A(\uart_tx_inst.prescale_reg[15] ),
    .B1(_0436_),
    .B2(_0443_),
    .ZN(_0444_));
 NAND2_X2 _1038_ (.A1(_0144_),
    .A2(_0146_),
    .ZN(_0445_));
 INV_X1 _1039_ (.A(_0445_),
    .ZN(_0446_));
 NAND2_X1 _1040_ (.A1(_0148_),
    .A2(_0150_),
    .ZN(_0447_));
 NOR3_X1 _1041_ (.A1(_0154_),
    .A2(_0274_),
    .A3(_0294_),
    .ZN(_0448_));
 XOR2_X1 _1042_ (.A(_0292_),
    .B(_0448_),
    .Z(_0449_));
 OAI21_X1 _1043_ (.A(_0446_),
    .B1(_0447_),
    .B2(_0449_),
    .ZN(_0450_));
 AOI21_X1 _1044_ (.A(_0403_),
    .B1(_0444_),
    .B2(_0450_),
    .ZN(_0066_));
 NOR4_X1 _1045_ (.A1(_0292_),
    .A2(_0153_),
    .A3(_0263_),
    .A4(_0294_),
    .ZN(_0451_));
 XNOR2_X1 _1046_ (.A(net3),
    .B(_0451_),
    .ZN(_0452_));
 OR4_X2 _1047_ (.A1(\uart_tx_inst.prescale_reg[15] ),
    .A2(\uart_tx_inst.prescale_reg[14] ),
    .A3(_0145_),
    .A4(_0424_),
    .ZN(_0453_));
 XOR2_X1 _1048_ (.A(\uart_tx_inst.prescale_reg[16] ),
    .B(_0453_),
    .Z(_0454_));
 MUX2_X1 _1049_ (.A(_0452_),
    .B(_0454_),
    .S(_0391_),
    .Z(_0455_));
 NOR2_X1 _1050_ (.A1(_0403_),
    .A2(_0455_),
    .ZN(_0067_));
 OAI21_X1 _1051_ (.A(\uart_tx_inst.prescale_reg[17] ),
    .B1(\uart_tx_inst.prescale_reg[16] ),
    .B2(_0445_),
    .ZN(_0456_));
 NOR2_X1 _1052_ (.A1(_0445_),
    .A2(_0149_),
    .ZN(_0457_));
 NOR4_X1 _1053_ (.A1(_0153_),
    .A2(_0274_),
    .A3(_0294_),
    .A4(_0311_),
    .ZN(_0458_));
 XOR2_X1 _1054_ (.A(net4),
    .B(_0458_),
    .Z(_0459_));
 OAI21_X1 _1055_ (.A(_0457_),
    .B1(_0459_),
    .B2(\uart_tx_inst.prescale_reg[18] ),
    .ZN(_0460_));
 AOI21_X1 _1056_ (.A(_0403_),
    .B1(_0456_),
    .B2(_0460_),
    .ZN(_0068_));
 NOR2_X1 _1057_ (.A1(\uart_tx_inst.prescale_reg[17] ),
    .A2(\uart_tx_inst.prescale_reg[16] ),
    .ZN(_0461_));
 NAND2_X1 _1058_ (.A1(\uart_tx_inst.prescale_reg[18] ),
    .A2(_0461_),
    .ZN(_0462_));
 OAI221_X1 _1059_ (.A(_0168_),
    .B1(_0148_),
    .B2(_0393_),
    .C1(_0453_),
    .C2(_0462_),
    .ZN(_0463_));
 AOI21_X1 _1060_ (.A(_0149_),
    .B1(_0453_),
    .B2(_0445_),
    .ZN(_0464_));
 NOR4_X1 _1061_ (.A1(_0154_),
    .A2(_0263_),
    .A3(_0294_),
    .A4(_0320_),
    .ZN(_0465_));
 XOR2_X1 _1062_ (.A(net5),
    .B(_0465_),
    .Z(_0466_));
 OAI21_X1 _1063_ (.A(_0464_),
    .B1(_0466_),
    .B2(_0445_),
    .ZN(_0467_));
 INV_X1 _1064_ (.A(\uart_tx_inst.prescale_reg[18] ),
    .ZN(_0468_));
 AOI21_X1 _1065_ (.A(_0463_),
    .B1(_0467_),
    .B2(_0468_),
    .ZN(_0069_));
 OR2_X1 _1066_ (.A1(_0607_),
    .A2(_0164_),
    .ZN(_0469_));
 NAND3_X1 _1067_ (.A1(_0148_),
    .A2(_0406_),
    .A3(_0164_),
    .ZN(_0470_));
 AOI21_X1 _1068_ (.A(_0209_),
    .B1(_0469_),
    .B2(_0470_),
    .ZN(_0070_));
 NOR2_X2 _1069_ (.A1(_0445_),
    .A2(_0447_),
    .ZN(_0471_));
 XOR2_X1 _1070_ (.A(_0140_),
    .B(_0409_),
    .Z(_0472_));
 AOI22_X1 _1071_ (.A1(_0471_),
    .A2(_0406_),
    .B1(_0393_),
    .B2(_0472_),
    .ZN(_0473_));
 NOR2_X1 _1072_ (.A1(_0182_),
    .A2(_0473_),
    .ZN(_0071_));
 XNOR2_X1 _1073_ (.A(_0081_),
    .B(_0154_),
    .ZN(_0474_));
 AOI22_X1 _1074_ (.A1(_0141_),
    .A2(_0393_),
    .B1(_0474_),
    .B2(_0471_),
    .ZN(_0475_));
 NOR2_X1 _1075_ (.A1(_0148_),
    .A2(_0393_),
    .ZN(_0476_));
 OR3_X1 _1076_ (.A1(\uart_tx_inst.prescale_reg[1] ),
    .A2(_0140_),
    .A3(\uart_tx_inst.prescale_reg[0] ),
    .ZN(_0477_));
 OAI21_X1 _1077_ (.A(\uart_tx_inst.prescale_reg[3] ),
    .B1(_0476_),
    .B2(_0477_),
    .ZN(_0478_));
 AOI21_X1 _1078_ (.A(_0209_),
    .B1(_0475_),
    .B2(_0478_),
    .ZN(_0072_));
 NOR2_X1 _1079_ (.A1(\uart_tx_inst.prescale_reg[3] ),
    .A2(_0140_),
    .ZN(_0479_));
 NAND2_X1 _1080_ (.A1(_0409_),
    .A2(_0479_),
    .ZN(_0480_));
 XOR2_X1 _1081_ (.A(_0142_),
    .B(_0480_),
    .Z(_0481_));
 MUX2_X1 _1082_ (.A(_0595_),
    .B(_0593_),
    .S(_0154_),
    .Z(_0482_));
 MUX2_X1 _1083_ (.A(_0481_),
    .B(_0482_),
    .S(_0164_),
    .Z(_0483_));
 NOR2_X1 _1084_ (.A1(_0403_),
    .A2(_0483_),
    .ZN(_0073_));
 INV_X1 _1085_ (.A(\uart_tx_inst.prescale_reg[1] ),
    .ZN(_0484_));
 INV_X1 _1086_ (.A(\uart_tx_inst.prescale_reg[0] ),
    .ZN(_0485_));
 NAND3_X1 _1087_ (.A1(_0484_),
    .A2(_0485_),
    .A3(_0479_),
    .ZN(_0486_));
 OAI21_X1 _1088_ (.A(\uart_tx_inst.prescale_reg[5] ),
    .B1(_0142_),
    .B2(_0486_),
    .ZN(_0487_));
 NAND2_X1 _1089_ (.A1(_0141_),
    .A2(_0143_),
    .ZN(_0488_));
 NAND2_X1 _1090_ (.A1(_0231_),
    .A2(_0406_),
    .ZN(_0489_));
 XOR2_X1 _1091_ (.A(_0232_),
    .B(_0489_),
    .Z(_0490_));
 AOI221_X1 _1092_ (.A(_0403_),
    .B1(_0487_),
    .B2(_0488_),
    .C1(_0490_),
    .C2(_0471_),
    .ZN(_0074_));
 AND2_X1 _1093_ (.A1(_0391_),
    .A2(_0411_),
    .ZN(_0491_));
 OAI21_X1 _1094_ (.A(_0138_),
    .B1(_0476_),
    .B2(_0491_),
    .ZN(_0492_));
 NOR3_X1 _1095_ (.A1(_0138_),
    .A2(_0164_),
    .A3(_0411_),
    .ZN(_0493_));
 NAND2_X1 _1096_ (.A1(_0406_),
    .A2(_0352_),
    .ZN(_0494_));
 XNOR2_X1 _1097_ (.A(_0233_),
    .B(_0494_),
    .ZN(_0495_));
 AOI21_X1 _1098_ (.A(_0493_),
    .B1(_0495_),
    .B2(_0471_),
    .ZN(_0496_));
 AOI21_X1 _1099_ (.A(_0209_),
    .B1(_0492_),
    .B2(_0496_),
    .ZN(_0075_));
 NOR2_X1 _1100_ (.A1(_0138_),
    .A2(_0488_),
    .ZN(_0497_));
 XNOR2_X1 _1101_ (.A(\uart_tx_inst.prescale_reg[7] ),
    .B(_0497_),
    .ZN(_0498_));
 NOR2_X1 _1102_ (.A1(_0154_),
    .A2(_0358_),
    .ZN(_0499_));
 XOR2_X1 _1103_ (.A(_0235_),
    .B(_0499_),
    .Z(_0500_));
 AOI21_X1 _1104_ (.A(_0393_),
    .B1(_0500_),
    .B2(_0148_),
    .ZN(_0501_));
 NOR3_X1 _1105_ (.A1(_0182_),
    .A2(_0498_),
    .A3(_0501_),
    .ZN(_0076_));
 NOR2_X1 _1106_ (.A1(_0408_),
    .A2(_0411_),
    .ZN(_0502_));
 XNOR2_X1 _1107_ (.A(\uart_tx_inst.prescale_reg[8] ),
    .B(_0502_),
    .ZN(_0503_));
 NOR2_X1 _1108_ (.A1(_0154_),
    .A2(_0368_),
    .ZN(_0504_));
 XNOR2_X1 _1109_ (.A(_0236_),
    .B(_0504_),
    .ZN(_0505_));
 MUX2_X1 _1110_ (.A(_0503_),
    .B(_0505_),
    .S(_0164_),
    .Z(_0506_));
 NOR2_X1 _1111_ (.A1(_0403_),
    .A2(_0506_),
    .ZN(_0077_));
 NOR2_X1 _1112_ (.A1(_0154_),
    .A2(_0274_),
    .ZN(_0507_));
 XNOR2_X1 _1113_ (.A(_0238_),
    .B(_0507_),
    .ZN(_0508_));
 NAND4_X1 _1114_ (.A1(_0484_),
    .A2(_0604_),
    .A3(_0139_),
    .A4(_0410_),
    .ZN(_0509_));
 XOR2_X1 _1115_ (.A(\uart_tx_inst.prescale_reg[9] ),
    .B(_0509_),
    .Z(_0510_));
 MUX2_X1 _1116_ (.A(_0508_),
    .B(_0510_),
    .S(_0391_),
    .Z(_0511_));
 NOR2_X1 _1117_ (.A1(_0403_),
    .A2(_0511_),
    .ZN(_0078_));
 NAND3_X1 _1118_ (.A1(net17),
    .A2(net30),
    .A3(_0135_),
    .ZN(_0512_));
 OAI21_X1 _1119_ (.A(_0512_),
    .B1(_0135_),
    .B2(net30),
    .ZN(_0513_));
 NOR2_X1 _1120_ (.A1(_0165_),
    .A2(_0513_),
    .ZN(_0079_));
 INV_X1 _1121_ (.A(\uart_tx_inst.data_reg[0] ),
    .ZN(_0514_));
 OAI21_X1 _1122_ (.A(_0406_),
    .B1(_0152_),
    .B2(_0514_),
    .ZN(_0515_));
 AOI221_X1 _1123_ (.A(_0082_),
    .B1(net32),
    .B2(_0151_),
    .C1(_0164_),
    .C2(_0515_),
    .ZN(_0516_));
 INV_X1 _1124_ (.A(_0516_),
    .ZN(_0080_));
 HA_X1 _1125_ (.A(_0588_),
    .B(_0589_),
    .CO(_0590_),
    .S(_0591_));
 HA_X1 _1126_ (.A(_0592_),
    .B(_0593_),
    .CO(_0594_),
    .S(_0595_));
 HA_X1 _1127_ (.A(_0596_),
    .B(_0597_),
    .CO(_0598_),
    .S(_0599_));
 HA_X1 _1128_ (.A(_0596_),
    .B(_0597_),
    .CO(_0600_),
    .S(_0601_));
 HA_X1 _1129_ (.A(\uart_rx_inst.bit_cnt[0] ),
    .B(_0597_),
    .CO(_0602_),
    .S(_0603_));
 HA_X1 _1130_ (.A(_0604_),
    .B(_0605_),
    .CO(_0606_),
    .S(_0607_));
 DFF_X2 \uart_rx_inst.bit_cnt[0]$_SDFFE_PP0P_  (.D(_0002_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\uart_rx_inst.bit_cnt[0] ),
    .QN(_0596_));
 DFF_X2 \uart_rx_inst.bit_cnt[1]$_SDFFE_PP0P_  (.D(_0003_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\uart_rx_inst.bit_cnt[1] ),
    .QN(_0597_));
 DFF_X1 \uart_rx_inst.bit_cnt[2]$_SDFFE_PP0P_  (.D(_0004_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\uart_rx_inst.bit_cnt[2] ),
    .QN(_0587_));
 DFF_X2 \uart_rx_inst.bit_cnt[3]$_SDFFE_PP0P_  (.D(_0005_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\uart_rx_inst.bit_cnt[3] ),
    .QN(_0001_));
 DFF_X1 \uart_rx_inst.busy_reg$_SDFFE_PP0P_  (.D(_0006_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net27),
    .QN(_0586_));
 DFF_X1 \uart_rx_inst.data_reg[0]$_SDFFCE_PP0P_  (.D(_0007_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\uart_rx_inst.data_reg[0] ),
    .QN(_0585_));
 DFF_X1 \uart_rx_inst.data_reg[1]$_SDFFCE_PP0P_  (.D(_0008_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\uart_rx_inst.data_reg[1] ),
    .QN(_0584_));
 DFF_X1 \uart_rx_inst.data_reg[2]$_SDFFCE_PP0P_  (.D(_0009_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\uart_rx_inst.data_reg[2] ),
    .QN(_0583_));
 DFF_X1 \uart_rx_inst.data_reg[3]$_SDFFCE_PP0P_  (.D(_0010_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\uart_rx_inst.data_reg[3] ),
    .QN(_0582_));
 DFF_X1 \uart_rx_inst.data_reg[4]$_SDFFCE_PP0P_  (.D(_0011_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\uart_rx_inst.data_reg[4] ),
    .QN(_0581_));
 DFF_X1 \uart_rx_inst.data_reg[5]$_SDFFCE_PP0P_  (.D(_0012_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\uart_rx_inst.data_reg[5] ),
    .QN(_0580_));
 DFF_X1 \uart_rx_inst.data_reg[6]$_SDFFCE_PP0P_  (.D(_0013_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\uart_rx_inst.data_reg[6] ),
    .QN(_0579_));
 DFF_X1 \uart_rx_inst.data_reg[7]$_SDFFCE_PP0P_  (.D(_0014_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\uart_rx_inst.data_reg[7] ),
    .QN(_0578_));
 DFF_X1 \uart_rx_inst.frame_error_reg$_SDFF_PP0_  (.D(_0015_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net28),
    .QN(_0577_));
 DFF_X1 \uart_rx_inst.m_axis_tdata_reg[0]$_SDFFE_PP0P_  (.D(_0016_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net18),
    .QN(_0576_));
 DFF_X1 \uart_rx_inst.m_axis_tdata_reg[1]$_SDFFE_PP0P_  (.D(_0017_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net19),
    .QN(_0575_));
 DFF_X1 \uart_rx_inst.m_axis_tdata_reg[2]$_SDFFE_PP0P_  (.D(_0018_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net20),
    .QN(_0574_));
 DFF_X1 \uart_rx_inst.m_axis_tdata_reg[3]$_SDFFE_PP0P_  (.D(_0019_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net21),
    .QN(_0573_));
 DFF_X1 \uart_rx_inst.m_axis_tdata_reg[4]$_SDFFE_PP0P_  (.D(_0020_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net22),
    .QN(_0572_));
 DFF_X1 \uart_rx_inst.m_axis_tdata_reg[5]$_SDFFE_PP0P_  (.D(_0021_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net23),
    .QN(_0571_));
 DFF_X1 \uart_rx_inst.m_axis_tdata_reg[6]$_SDFFE_PP0P_  (.D(_0022_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net24),
    .QN(_0570_));
 DFF_X1 \uart_rx_inst.m_axis_tdata_reg[7]$_SDFFE_PP0P_  (.D(_0023_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net25),
    .QN(_0569_));
 DFF_X1 \uart_rx_inst.m_axis_tvalid_reg$_SDFF_PP0_  (.D(_0024_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net26),
    .QN(_0568_));
 DFF_X1 \uart_rx_inst.overrun_error_reg$_SDFF_PP0_  (.D(_0025_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net29),
    .QN(_0567_));
 DFF_X1 \uart_rx_inst.prescale_reg[0]$_SDFFE_PP0P_  (.D(_0026_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[0] ),
    .QN(_0588_));
 DFF_X1 \uart_rx_inst.prescale_reg[10]$_SDFFE_PP0P_  (.D(_0027_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[10] ),
    .QN(_0566_));
 DFF_X1 \uart_rx_inst.prescale_reg[11]$_SDFFE_PP0P_  (.D(_0028_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[11] ),
    .QN(_0565_));
 DFF_X1 \uart_rx_inst.prescale_reg[12]$_SDFFE_PP0P_  (.D(_0029_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[12] ),
    .QN(_0564_));
 DFF_X1 \uart_rx_inst.prescale_reg[13]$_SDFFE_PP0P_  (.D(_0030_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[13] ),
    .QN(_0563_));
 DFF_X1 \uart_rx_inst.prescale_reg[14]$_SDFFE_PP0P_  (.D(_0031_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[14] ),
    .QN(_0562_));
 DFF_X1 \uart_rx_inst.prescale_reg[15]$_SDFFE_PP0P_  (.D(_0032_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[15] ),
    .QN(_0561_));
 DFF_X1 \uart_rx_inst.prescale_reg[16]$_SDFFE_PP0P_  (.D(_0033_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[16] ),
    .QN(_0560_));
 DFF_X1 \uart_rx_inst.prescale_reg[17]$_SDFFE_PP0P_  (.D(_0034_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[17] ),
    .QN(_0559_));
 DFF_X1 \uart_rx_inst.prescale_reg[18]$_SDFFE_PP0P_  (.D(_0035_),
    .CK(clknet_3_7__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[18] ),
    .QN(_0558_));
 DFF_X1 \uart_rx_inst.prescale_reg[1]$_SDFFE_PP0P_  (.D(_0036_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[1] ),
    .QN(_0589_));
 DFF_X1 \uart_rx_inst.prescale_reg[2]$_SDFFE_PP0P_  (.D(_0037_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[2] ),
    .QN(_0557_));
 DFF_X2 \uart_rx_inst.prescale_reg[3]$_SDFFE_PP0P_  (.D(_0038_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[3] ),
    .QN(_0556_));
 DFF_X2 \uart_rx_inst.prescale_reg[4]$_SDFFE_PP0P_  (.D(_0039_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[4] ),
    .QN(_0555_));
 DFF_X1 \uart_rx_inst.prescale_reg[5]$_SDFFE_PP0P_  (.D(_0040_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[5] ),
    .QN(_0554_));
 DFF_X2 \uart_rx_inst.prescale_reg[6]$_SDFFE_PP0P_  (.D(_0041_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[6] ),
    .QN(_0553_));
 DFF_X2 \uart_rx_inst.prescale_reg[7]$_SDFFE_PP0P_  (.D(_0042_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[7] ),
    .QN(_0552_));
 DFF_X2 \uart_rx_inst.prescale_reg[8]$_SDFFE_PP0P_  (.D(_0043_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[8] ),
    .QN(_0551_));
 DFF_X1 \uart_rx_inst.prescale_reg[9]$_SDFFE_PP0P_  (.D(_0044_),
    .CK(clknet_3_6__leaf_clk),
    .Q(\uart_rx_inst.prescale_reg[9] ),
    .QN(_0550_));
 DFF_X1 \uart_rx_inst.rxd_reg$_SDFF_PP1_  (.D(_0045_),
    .CK(clknet_3_3__leaf_clk),
    .Q(\uart_rx_inst.rxd_reg ),
    .QN(_0000_));
 DFF_X1 \uart_tx_inst.bit_cnt[0]$_SDFFE_PP0P_  (.D(_0046_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\uart_tx_inst.bit_cnt[0] ),
    .QN(_0549_));
 DFF_X1 \uart_tx_inst.bit_cnt[1]$_SDFFE_PP0P_  (.D(_0047_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\uart_tx_inst.bit_cnt[1] ),
    .QN(_0548_));
 DFF_X1 \uart_tx_inst.bit_cnt[2]$_SDFFE_PP0P_  (.D(_0048_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\uart_tx_inst.bit_cnt[2] ),
    .QN(_0547_));
 DFF_X2 \uart_tx_inst.bit_cnt[3]$_SDFFE_PP0P_  (.D(_0049_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\uart_tx_inst.bit_cnt[3] ),
    .QN(_0546_));
 DFF_X1 \uart_tx_inst.busy_reg$_SDFFE_PP0P_  (.D(_0050_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net31),
    .QN(_0545_));
 DFF_X1 \uart_tx_inst.data_reg[0]$_DFFE_PP_  (.D(_0051_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\uart_tx_inst.data_reg[0] ),
    .QN(_0544_));
 DFF_X1 \uart_tx_inst.data_reg[1]$_DFFE_PP_  (.D(_0052_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\uart_tx_inst.data_reg[1] ),
    .QN(_0543_));
 DFF_X1 \uart_tx_inst.data_reg[2]$_DFFE_PP_  (.D(_0053_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\uart_tx_inst.data_reg[2] ),
    .QN(_0542_));
 DFF_X1 \uart_tx_inst.data_reg[3]$_DFFE_PP_  (.D(_0054_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\uart_tx_inst.data_reg[3] ),
    .QN(_0541_));
 DFF_X1 \uart_tx_inst.data_reg[4]$_DFFE_PP_  (.D(_0055_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\uart_tx_inst.data_reg[4] ),
    .QN(_0540_));
 DFF_X1 \uart_tx_inst.data_reg[5]$_DFFE_PP_  (.D(_0056_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\uart_tx_inst.data_reg[5] ),
    .QN(_0539_));
 DFF_X1 \uart_tx_inst.data_reg[6]$_DFFE_PP_  (.D(_0057_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\uart_tx_inst.data_reg[6] ),
    .QN(_0538_));
 DFF_X1 \uart_tx_inst.data_reg[7]$_DFFE_PP_  (.D(_0058_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\uart_tx_inst.data_reg[7] ),
    .QN(_0537_));
 DFF_X1 \uart_tx_inst.data_reg[8]$_DFFE_PP_  (.D(_0059_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\uart_tx_inst.data_reg[8] ),
    .QN(_0536_));
 DFF_X1 \uart_tx_inst.prescale_reg[0]$_SDFFE_PP0P_  (.D(_0060_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[0] ),
    .QN(_0604_));
 DFF_X1 \uart_tx_inst.prescale_reg[10]$_SDFFE_PP0P_  (.D(_0061_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[10] ),
    .QN(_0535_));
 DFF_X1 \uart_tx_inst.prescale_reg[11]$_SDFFE_PP0P_  (.D(_0062_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[11] ),
    .QN(_0534_));
 DFF_X1 \uart_tx_inst.prescale_reg[12]$_SDFFE_PP0P_  (.D(_0063_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[12] ),
    .QN(_0533_));
 DFF_X1 \uart_tx_inst.prescale_reg[13]$_SDFFE_PP0P_  (.D(_0064_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[13] ),
    .QN(_0532_));
 DFF_X2 \uart_tx_inst.prescale_reg[14]$_SDFFE_PP0P_  (.D(_0065_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[14] ),
    .QN(_0531_));
 DFF_X2 \uart_tx_inst.prescale_reg[15]$_SDFFE_PP0P_  (.D(_0066_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[15] ),
    .QN(_0530_));
 DFF_X1 \uart_tx_inst.prescale_reg[16]$_SDFFE_PP0P_  (.D(_0067_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[16] ),
    .QN(_0529_));
 DFF_X1 \uart_tx_inst.prescale_reg[17]$_SDFFE_PP0P_  (.D(_0068_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[17] ),
    .QN(_0528_));
 DFF_X1 \uart_tx_inst.prescale_reg[18]$_SDFFE_PP0P_  (.D(_0069_),
    .CK(clknet_3_5__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[18] ),
    .QN(_0527_));
 DFF_X1 \uart_tx_inst.prescale_reg[1]$_SDFFE_PP0P_  (.D(_0070_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[1] ),
    .QN(_0605_));
 DFF_X1 \uart_tx_inst.prescale_reg[2]$_SDFFE_PP0P_  (.D(_0071_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[2] ),
    .QN(_0526_));
 DFF_X2 \uart_tx_inst.prescale_reg[3]$_SDFFE_PP0P_  (.D(_0072_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[3] ),
    .QN(_0525_));
 DFF_X1 \uart_tx_inst.prescale_reg[4]$_SDFFE_PP0P_  (.D(_0073_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[4] ),
    .QN(_0524_));
 DFF_X2 \uart_tx_inst.prescale_reg[5]$_SDFFE_PP0P_  (.D(_0074_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[5] ),
    .QN(_0523_));
 DFF_X1 \uart_tx_inst.prescale_reg[6]$_SDFFE_PP0P_  (.D(_0075_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[6] ),
    .QN(_0522_));
 DFF_X1 \uart_tx_inst.prescale_reg[7]$_SDFFE_PP0P_  (.D(_0076_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[7] ),
    .QN(_0521_));
 DFF_X1 \uart_tx_inst.prescale_reg[8]$_SDFFE_PP0P_  (.D(_0077_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[8] ),
    .QN(_0520_));
 DFF_X1 \uart_tx_inst.prescale_reg[9]$_SDFFE_PP0P_  (.D(_0078_),
    .CK(clknet_3_4__leaf_clk),
    .Q(\uart_tx_inst.prescale_reg[9] ),
    .QN(_0519_));
 DFF_X1 \uart_tx_inst.s_axis_tready_reg$_SDFFE_PP0P_  (.D(_0079_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net30),
    .QN(_0518_));
 DFF_X1 \uart_tx_inst.txd_reg$_SDFFE_PP1P_  (.D(_0080_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net32),
    .QN(_0517_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_69 ();
 BUF_X1 input1 (.A(m_axis_tready),
    .Z(net1));
 BUF_X1 input2 (.A(prescale[11]),
    .Z(net2));
 BUF_X1 input3 (.A(prescale[13]),
    .Z(net3));
 BUF_X1 input4 (.A(prescale[14]),
    .Z(net4));
 BUF_X1 input5 (.A(prescale[15]),
    .Z(net5));
 BUF_X1 input6 (.A(prescale[1]),
    .Z(net6));
 BUF_X1 input7 (.A(prescale[9]),
    .Z(net7));
 BUF_X1 input8 (.A(rxd),
    .Z(net8));
 BUF_X1 input9 (.A(s_axis_tdata[0]),
    .Z(net9));
 BUF_X1 input10 (.A(s_axis_tdata[1]),
    .Z(net10));
 BUF_X1 input11 (.A(s_axis_tdata[2]),
    .Z(net11));
 BUF_X1 input12 (.A(s_axis_tdata[3]),
    .Z(net12));
 BUF_X1 input13 (.A(s_axis_tdata[4]),
    .Z(net13));
 BUF_X1 input14 (.A(s_axis_tdata[5]),
    .Z(net14));
 BUF_X1 input15 (.A(s_axis_tdata[6]),
    .Z(net15));
 BUF_X1 input16 (.A(s_axis_tdata[7]),
    .Z(net16));
 BUF_X1 input17 (.A(s_axis_tvalid),
    .Z(net17));
 BUF_X1 output18 (.A(net18),
    .Z(m_axis_tdata[0]));
 BUF_X1 output19 (.A(net19),
    .Z(m_axis_tdata[1]));
 BUF_X1 output20 (.A(net20),
    .Z(m_axis_tdata[2]));
 BUF_X1 output21 (.A(net21),
    .Z(m_axis_tdata[3]));
 BUF_X1 output22 (.A(net22),
    .Z(m_axis_tdata[4]));
 BUF_X1 output23 (.A(net23),
    .Z(m_axis_tdata[5]));
 BUF_X1 output24 (.A(net24),
    .Z(m_axis_tdata[6]));
 BUF_X1 output25 (.A(net25),
    .Z(m_axis_tdata[7]));
 BUF_X1 output26 (.A(net26),
    .Z(m_axis_tvalid));
 BUF_X1 output27 (.A(net27),
    .Z(rx_busy));
 BUF_X1 output28 (.A(net28),
    .Z(rx_frame_error));
 BUF_X1 output29 (.A(net29),
    .Z(rx_overrun_error));
 BUF_X1 output30 (.A(net30),
    .Z(s_axis_tready));
 BUF_X1 output31 (.A(net31),
    .Z(tx_busy));
 BUF_X1 output32 (.A(net32),
    .Z(txd));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 CLKBUF_X3 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 CLKBUF_X3 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 CLKBUF_X3 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 CLKBUF_X3 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 CLKBUF_X3 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 CLKBUF_X3 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 CLKBUF_X3 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 INV_X4 clkload0 (.A(clknet_3_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_3_1__leaf_clk));
 INV_X4 clkload2 (.A(clknet_3_3__leaf_clk));
 INV_X4 clkload3 (.A(clknet_3_4__leaf_clk));
 INV_X4 clkload4 (.A(clknet_3_5__leaf_clk));
 INV_X4 clkload5 (.A(clknet_3_6__leaf_clk));
 INV_X4 clkload6 (.A(clknet_3_7__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_33 ();
 FILLCELL_X4 FILLER_0_41 ();
 FILLCELL_X1 FILLER_0_64 ();
 FILLCELL_X8 FILLER_0_68 ();
 FILLCELL_X8 FILLER_0_89 ();
 FILLCELL_X2 FILLER_0_103 ();
 FILLCELL_X1 FILLER_0_105 ();
 FILLCELL_X1 FILLER_0_109 ();
 FILLCELL_X16 FILLER_0_116 ();
 FILLCELL_X4 FILLER_0_132 ();
 FILLCELL_X2 FILLER_0_136 ();
 FILLCELL_X32 FILLER_0_155 ();
 FILLCELL_X32 FILLER_0_187 ();
 FILLCELL_X32 FILLER_0_219 ();
 FILLCELL_X8 FILLER_0_251 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_17 ();
 FILLCELL_X1 FILLER_1_19 ();
 FILLCELL_X2 FILLER_1_61 ();
 FILLCELL_X1 FILLER_1_87 ();
 FILLCELL_X1 FILLER_1_95 ();
 FILLCELL_X1 FILLER_1_100 ();
 FILLCELL_X1 FILLER_1_105 ();
 FILLCELL_X16 FILLER_1_120 ();
 FILLCELL_X1 FILLER_1_136 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X2 FILLER_1_257 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X1 FILLER_2_33 ();
 FILLCELL_X8 FILLER_2_55 ();
 FILLCELL_X1 FILLER_2_63 ();
 FILLCELL_X4 FILLER_2_81 ();
 FILLCELL_X2 FILLER_2_105 ();
 FILLCELL_X1 FILLER_2_107 ();
 FILLCELL_X1 FILLER_2_149 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X2 FILLER_2_257 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X4 FILLER_3_33 ();
 FILLCELL_X1 FILLER_3_37 ();
 FILLCELL_X16 FILLER_3_59 ();
 FILLCELL_X4 FILLER_3_75 ();
 FILLCELL_X2 FILLER_3_79 ();
 FILLCELL_X1 FILLER_3_81 ();
 FILLCELL_X1 FILLER_3_103 ();
 FILLCELL_X2 FILLER_3_111 ();
 FILLCELL_X1 FILLER_3_113 ();
 FILLCELL_X32 FILLER_3_159 ();
 FILLCELL_X32 FILLER_3_191 ();
 FILLCELL_X32 FILLER_3_223 ();
 FILLCELL_X4 FILLER_3_255 ();
 FILLCELL_X16 FILLER_4_1 ();
 FILLCELL_X8 FILLER_4_17 ();
 FILLCELL_X4 FILLER_4_25 ();
 FILLCELL_X2 FILLER_4_29 ();
 FILLCELL_X1 FILLER_4_31 ();
 FILLCELL_X1 FILLER_4_49 ();
 FILLCELL_X4 FILLER_4_81 ();
 FILLCELL_X2 FILLER_4_85 ();
 FILLCELL_X1 FILLER_4_87 ();
 FILLCELL_X8 FILLER_4_92 ();
 FILLCELL_X4 FILLER_4_100 ();
 FILLCELL_X1 FILLER_4_104 ();
 FILLCELL_X4 FILLER_4_110 ();
 FILLCELL_X1 FILLER_4_114 ();
 FILLCELL_X8 FILLER_4_117 ();
 FILLCELL_X1 FILLER_4_125 ();
 FILLCELL_X4 FILLER_4_130 ();
 FILLCELL_X4 FILLER_4_148 ();
 FILLCELL_X8 FILLER_4_159 ();
 FILLCELL_X4 FILLER_4_167 ();
 FILLCELL_X4 FILLER_4_176 ();
 FILLCELL_X1 FILLER_4_197 ();
 FILLCELL_X32 FILLER_4_215 ();
 FILLCELL_X8 FILLER_4_247 ();
 FILLCELL_X4 FILLER_4_255 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X4 FILLER_5_33 ();
 FILLCELL_X16 FILLER_5_54 ();
 FILLCELL_X2 FILLER_5_70 ();
 FILLCELL_X1 FILLER_5_72 ();
 FILLCELL_X1 FILLER_5_95 ();
 FILLCELL_X4 FILLER_5_113 ();
 FILLCELL_X1 FILLER_5_117 ();
 FILLCELL_X16 FILLER_5_131 ();
 FILLCELL_X2 FILLER_5_147 ();
 FILLCELL_X1 FILLER_5_149 ();
 FILLCELL_X1 FILLER_5_167 ();
 FILLCELL_X8 FILLER_5_173 ();
 FILLCELL_X2 FILLER_5_184 ();
 FILLCELL_X1 FILLER_5_192 ();
 FILLCELL_X1 FILLER_5_200 ();
 FILLCELL_X1 FILLER_5_208 ();
 FILLCELL_X32 FILLER_5_212 ();
 FILLCELL_X8 FILLER_5_244 ();
 FILLCELL_X4 FILLER_5_252 ();
 FILLCELL_X2 FILLER_5_256 ();
 FILLCELL_X1 FILLER_5_258 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X2 FILLER_6_97 ();
 FILLCELL_X16 FILLER_6_111 ();
 FILLCELL_X8 FILLER_6_127 ();
 FILLCELL_X4 FILLER_6_144 ();
 FILLCELL_X2 FILLER_6_155 ();
 FILLCELL_X1 FILLER_6_157 ();
 FILLCELL_X16 FILLER_6_163 ();
 FILLCELL_X1 FILLER_6_179 ();
 FILLCELL_X4 FILLER_6_184 ();
 FILLCELL_X1 FILLER_6_188 ();
 FILLCELL_X2 FILLER_6_203 ();
 FILLCELL_X32 FILLER_6_211 ();
 FILLCELL_X16 FILLER_6_243 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X4 FILLER_7_65 ();
 FILLCELL_X2 FILLER_7_69 ();
 FILLCELL_X1 FILLER_7_71 ();
 FILLCELL_X2 FILLER_7_96 ();
 FILLCELL_X2 FILLER_7_101 ();
 FILLCELL_X2 FILLER_7_144 ();
 FILLCELL_X16 FILLER_7_149 ();
 FILLCELL_X2 FILLER_7_165 ();
 FILLCELL_X4 FILLER_7_222 ();
 FILLCELL_X2 FILLER_7_245 ();
 FILLCELL_X4 FILLER_7_254 ();
 FILLCELL_X1 FILLER_7_258 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X16 FILLER_8_33 ();
 FILLCELL_X8 FILLER_8_49 ();
 FILLCELL_X2 FILLER_8_57 ();
 FILLCELL_X2 FILLER_8_86 ();
 FILLCELL_X4 FILLER_8_99 ();
 FILLCELL_X4 FILLER_8_107 ();
 FILLCELL_X2 FILLER_8_111 ();
 FILLCELL_X1 FILLER_8_113 ();
 FILLCELL_X1 FILLER_8_131 ();
 FILLCELL_X4 FILLER_8_143 ();
 FILLCELL_X1 FILLER_8_147 ();
 FILLCELL_X2 FILLER_8_188 ();
 FILLCELL_X2 FILLER_8_213 ();
 FILLCELL_X1 FILLER_8_215 ();
 FILLCELL_X1 FILLER_8_219 ();
 FILLCELL_X2 FILLER_8_226 ();
 FILLCELL_X16 FILLER_8_231 ();
 FILLCELL_X8 FILLER_8_247 ();
 FILLCELL_X4 FILLER_8_255 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X8 FILLER_9_49 ();
 FILLCELL_X4 FILLER_9_57 ();
 FILLCELL_X1 FILLER_9_61 ();
 FILLCELL_X2 FILLER_9_84 ();
 FILLCELL_X1 FILLER_9_102 ();
 FILLCELL_X2 FILLER_9_123 ();
 FILLCELL_X2 FILLER_9_131 ();
 FILLCELL_X1 FILLER_9_133 ();
 FILLCELL_X1 FILLER_9_137 ();
 FILLCELL_X2 FILLER_9_155 ();
 FILLCELL_X2 FILLER_9_181 ();
 FILLCELL_X1 FILLER_9_183 ();
 FILLCELL_X4 FILLER_9_197 ();
 FILLCELL_X1 FILLER_9_201 ();
 FILLCELL_X2 FILLER_9_219 ();
 FILLCELL_X1 FILLER_9_221 ();
 FILLCELL_X16 FILLER_9_229 ();
 FILLCELL_X8 FILLER_9_245 ();
 FILLCELL_X4 FILLER_9_253 ();
 FILLCELL_X2 FILLER_9_257 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X8 FILLER_10_33 ();
 FILLCELL_X4 FILLER_10_41 ();
 FILLCELL_X2 FILLER_10_45 ();
 FILLCELL_X1 FILLER_10_47 ();
 FILLCELL_X2 FILLER_10_70 ();
 FILLCELL_X1 FILLER_10_85 ();
 FILLCELL_X2 FILLER_10_100 ();
 FILLCELL_X2 FILLER_10_105 ();
 FILLCELL_X1 FILLER_10_107 ();
 FILLCELL_X1 FILLER_10_114 ();
 FILLCELL_X1 FILLER_10_118 ();
 FILLCELL_X2 FILLER_10_140 ();
 FILLCELL_X1 FILLER_10_148 ();
 FILLCELL_X8 FILLER_10_164 ();
 FILLCELL_X4 FILLER_10_172 ();
 FILLCELL_X2 FILLER_10_209 ();
 FILLCELL_X32 FILLER_10_217 ();
 FILLCELL_X8 FILLER_10_249 ();
 FILLCELL_X2 FILLER_10_257 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X16 FILLER_11_33 ();
 FILLCELL_X4 FILLER_11_49 ();
 FILLCELL_X2 FILLER_11_53 ();
 FILLCELL_X4 FILLER_11_77 ();
 FILLCELL_X2 FILLER_11_124 ();
 FILLCELL_X2 FILLER_11_130 ();
 FILLCELL_X16 FILLER_11_158 ();
 FILLCELL_X8 FILLER_11_174 ();
 FILLCELL_X4 FILLER_11_182 ();
 FILLCELL_X2 FILLER_11_186 ();
 FILLCELL_X1 FILLER_11_188 ();
 FILLCELL_X32 FILLER_11_224 ();
 FILLCELL_X2 FILLER_11_256 ();
 FILLCELL_X1 FILLER_11_258 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X8 FILLER_12_65 ();
 FILLCELL_X4 FILLER_12_73 ();
 FILLCELL_X2 FILLER_12_77 ();
 FILLCELL_X1 FILLER_12_79 ();
 FILLCELL_X2 FILLER_12_89 ();
 FILLCELL_X1 FILLER_12_95 ();
 FILLCELL_X2 FILLER_12_102 ();
 FILLCELL_X2 FILLER_12_121 ();
 FILLCELL_X2 FILLER_12_127 ();
 FILLCELL_X4 FILLER_12_132 ();
 FILLCELL_X2 FILLER_12_136 ();
 FILLCELL_X1 FILLER_12_138 ();
 FILLCELL_X16 FILLER_12_149 ();
 FILLCELL_X2 FILLER_12_165 ();
 FILLCELL_X1 FILLER_12_167 ();
 FILLCELL_X1 FILLER_12_205 ();
 FILLCELL_X8 FILLER_12_209 ();
 FILLCELL_X16 FILLER_12_234 ();
 FILLCELL_X8 FILLER_12_250 ();
 FILLCELL_X1 FILLER_12_258 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X4 FILLER_13_65 ();
 FILLCELL_X2 FILLER_13_69 ();
 FILLCELL_X1 FILLER_13_71 ();
 FILLCELL_X8 FILLER_13_98 ();
 FILLCELL_X4 FILLER_13_106 ();
 FILLCELL_X2 FILLER_13_110 ();
 FILLCELL_X1 FILLER_13_112 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X16 FILLER_13_193 ();
 FILLCELL_X2 FILLER_13_209 ();
 FILLCELL_X32 FILLER_13_217 ();
 FILLCELL_X8 FILLER_13_249 ();
 FILLCELL_X2 FILLER_13_257 ();
 FILLCELL_X32 FILLER_14_18 ();
 FILLCELL_X8 FILLER_14_50 ();
 FILLCELL_X1 FILLER_14_58 ();
 FILLCELL_X1 FILLER_14_76 ();
 FILLCELL_X8 FILLER_14_81 ();
 FILLCELL_X2 FILLER_14_89 ();
 FILLCELL_X1 FILLER_14_91 ();
 FILLCELL_X2 FILLER_14_95 ();
 FILLCELL_X2 FILLER_14_103 ();
 FILLCELL_X1 FILLER_14_105 ();
 FILLCELL_X4 FILLER_14_109 ();
 FILLCELL_X2 FILLER_14_113 ();
 FILLCELL_X4 FILLER_14_118 ();
 FILLCELL_X16 FILLER_14_125 ();
 FILLCELL_X8 FILLER_14_141 ();
 FILLCELL_X4 FILLER_14_149 ();
 FILLCELL_X2 FILLER_14_153 ();
 FILLCELL_X16 FILLER_14_164 ();
 FILLCELL_X2 FILLER_14_180 ();
 FILLCELL_X1 FILLER_14_182 ();
 FILLCELL_X4 FILLER_14_189 ();
 FILLCELL_X2 FILLER_14_209 ();
 FILLCELL_X2 FILLER_14_216 ();
 FILLCELL_X1 FILLER_14_218 ();
 FILLCELL_X1 FILLER_14_225 ();
 FILLCELL_X4 FILLER_14_232 ();
 FILLCELL_X2 FILLER_14_236 ();
 FILLCELL_X1 FILLER_14_238 ();
 FILLCELL_X1 FILLER_14_242 ();
 FILLCELL_X8 FILLER_14_246 ();
 FILLCELL_X4 FILLER_14_254 ();
 FILLCELL_X1 FILLER_14_258 ();
 FILLCELL_X2 FILLER_15_29 ();
 FILLCELL_X32 FILLER_15_34 ();
 FILLCELL_X16 FILLER_15_66 ();
 FILLCELL_X8 FILLER_15_82 ();
 FILLCELL_X4 FILLER_15_90 ();
 FILLCELL_X2 FILLER_15_94 ();
 FILLCELL_X1 FILLER_15_96 ();
 FILLCELL_X2 FILLER_15_99 ();
 FILLCELL_X1 FILLER_15_101 ();
 FILLCELL_X8 FILLER_15_113 ();
 FILLCELL_X4 FILLER_15_121 ();
 FILLCELL_X2 FILLER_15_147 ();
 FILLCELL_X1 FILLER_15_172 ();
 FILLCELL_X2 FILLER_15_188 ();
 FILLCELL_X1 FILLER_15_196 ();
 FILLCELL_X2 FILLER_15_202 ();
 FILLCELL_X1 FILLER_15_207 ();
 FILLCELL_X2 FILLER_15_212 ();
 FILLCELL_X8 FILLER_15_245 ();
 FILLCELL_X2 FILLER_15_253 ();
 FILLCELL_X1 FILLER_16_4 ();
 FILLCELL_X2 FILLER_16_35 ();
 FILLCELL_X8 FILLER_16_40 ();
 FILLCELL_X4 FILLER_16_48 ();
 FILLCELL_X8 FILLER_16_81 ();
 FILLCELL_X4 FILLER_16_89 ();
 FILLCELL_X1 FILLER_16_93 ();
 FILLCELL_X4 FILLER_16_110 ();
 FILLCELL_X1 FILLER_16_114 ();
 FILLCELL_X2 FILLER_16_131 ();
 FILLCELL_X4 FILLER_16_155 ();
 FILLCELL_X8 FILLER_16_162 ();
 FILLCELL_X2 FILLER_16_170 ();
 FILLCELL_X1 FILLER_16_176 ();
 FILLCELL_X1 FILLER_16_193 ();
 FILLCELL_X2 FILLER_16_198 ();
 FILLCELL_X2 FILLER_16_206 ();
 FILLCELL_X2 FILLER_16_217 ();
 FILLCELL_X1 FILLER_16_219 ();
 FILLCELL_X8 FILLER_16_240 ();
 FILLCELL_X1 FILLER_16_248 ();
 FILLCELL_X2 FILLER_16_252 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_9 ();
 FILLCELL_X4 FILLER_17_16 ();
 FILLCELL_X2 FILLER_17_20 ();
 FILLCELL_X1 FILLER_17_22 ();
 FILLCELL_X8 FILLER_17_46 ();
 FILLCELL_X2 FILLER_17_54 ();
 FILLCELL_X2 FILLER_17_85 ();
 FILLCELL_X2 FILLER_17_91 ();
 FILLCELL_X1 FILLER_17_93 ();
 FILLCELL_X4 FILLER_17_101 ();
 FILLCELL_X2 FILLER_17_111 ();
 FILLCELL_X1 FILLER_17_126 ();
 FILLCELL_X8 FILLER_17_142 ();
 FILLCELL_X2 FILLER_17_150 ();
 FILLCELL_X4 FILLER_17_170 ();
 FILLCELL_X2 FILLER_17_183 ();
 FILLCELL_X1 FILLER_17_185 ();
 FILLCELL_X1 FILLER_17_192 ();
 FILLCELL_X4 FILLER_17_201 ();
 FILLCELL_X2 FILLER_17_227 ();
 FILLCELL_X1 FILLER_17_229 ();
 FILLCELL_X4 FILLER_17_233 ();
 FILLCELL_X4 FILLER_17_240 ();
 FILLCELL_X2 FILLER_17_244 ();
 FILLCELL_X4 FILLER_17_253 ();
 FILLCELL_X2 FILLER_17_257 ();
 FILLCELL_X2 FILLER_18_1 ();
 FILLCELL_X8 FILLER_18_6 ();
 FILLCELL_X4 FILLER_18_14 ();
 FILLCELL_X4 FILLER_18_21 ();
 FILLCELL_X1 FILLER_18_25 ();
 FILLCELL_X8 FILLER_18_40 ();
 FILLCELL_X4 FILLER_18_48 ();
 FILLCELL_X2 FILLER_18_52 ();
 FILLCELL_X1 FILLER_18_54 ();
 FILLCELL_X1 FILLER_18_59 ();
 FILLCELL_X2 FILLER_18_81 ();
 FILLCELL_X1 FILLER_18_83 ();
 FILLCELL_X1 FILLER_18_87 ();
 FILLCELL_X4 FILLER_18_92 ();
 FILLCELL_X2 FILLER_18_96 ();
 FILLCELL_X8 FILLER_18_105 ();
 FILLCELL_X2 FILLER_18_113 ();
 FILLCELL_X1 FILLER_18_115 ();
 FILLCELL_X8 FILLER_18_124 ();
 FILLCELL_X4 FILLER_18_132 ();
 FILLCELL_X1 FILLER_18_136 ();
 FILLCELL_X8 FILLER_18_142 ();
 FILLCELL_X4 FILLER_18_150 ();
 FILLCELL_X1 FILLER_18_154 ();
 FILLCELL_X4 FILLER_18_171 ();
 FILLCELL_X2 FILLER_18_175 ();
 FILLCELL_X4 FILLER_18_181 ();
 FILLCELL_X1 FILLER_18_202 ();
 FILLCELL_X8 FILLER_18_212 ();
 FILLCELL_X32 FILLER_18_223 ();
 FILLCELL_X4 FILLER_18_255 ();
 FILLCELL_X2 FILLER_19_1 ();
 FILLCELL_X1 FILLER_19_24 ();
 FILLCELL_X16 FILLER_19_42 ();
 FILLCELL_X1 FILLER_19_58 ();
 FILLCELL_X1 FILLER_19_70 ();
 FILLCELL_X2 FILLER_19_74 ();
 FILLCELL_X1 FILLER_19_76 ();
 FILLCELL_X4 FILLER_19_80 ();
 FILLCELL_X8 FILLER_19_89 ();
 FILLCELL_X1 FILLER_19_97 ();
 FILLCELL_X1 FILLER_19_130 ();
 FILLCELL_X2 FILLER_19_138 ();
 FILLCELL_X8 FILLER_19_151 ();
 FILLCELL_X2 FILLER_19_159 ();
 FILLCELL_X2 FILLER_19_165 ();
 FILLCELL_X1 FILLER_19_176 ();
 FILLCELL_X1 FILLER_19_183 ();
 FILLCELL_X2 FILLER_19_193 ();
 FILLCELL_X1 FILLER_19_195 ();
 FILLCELL_X8 FILLER_19_199 ();
 FILLCELL_X4 FILLER_19_207 ();
 FILLCELL_X2 FILLER_19_211 ();
 FILLCELL_X1 FILLER_19_213 ();
 FILLCELL_X8 FILLER_19_218 ();
 FILLCELL_X4 FILLER_19_226 ();
 FILLCELL_X1 FILLER_19_230 ();
 FILLCELL_X8 FILLER_19_248 ();
 FILLCELL_X2 FILLER_19_256 ();
 FILLCELL_X1 FILLER_19_258 ();
 FILLCELL_X2 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_27 ();
 FILLCELL_X1 FILLER_20_29 ();
 FILLCELL_X16 FILLER_20_36 ();
 FILLCELL_X8 FILLER_20_52 ();
 FILLCELL_X4 FILLER_20_60 ();
 FILLCELL_X1 FILLER_20_74 ();
 FILLCELL_X1 FILLER_20_115 ();
 FILLCELL_X8 FILLER_20_123 ();
 FILLCELL_X8 FILLER_20_150 ();
 FILLCELL_X1 FILLER_20_158 ();
 FILLCELL_X4 FILLER_20_168 ();
 FILLCELL_X2 FILLER_20_172 ();
 FILLCELL_X1 FILLER_20_174 ();
 FILLCELL_X4 FILLER_20_179 ();
 FILLCELL_X8 FILLER_20_197 ();
 FILLCELL_X1 FILLER_20_209 ();
 FILLCELL_X1 FILLER_20_219 ();
 FILLCELL_X1 FILLER_20_225 ();
 FILLCELL_X1 FILLER_20_230 ();
 FILLCELL_X4 FILLER_20_252 ();
 FILLCELL_X2 FILLER_20_256 ();
 FILLCELL_X1 FILLER_20_258 ();
 FILLCELL_X2 FILLER_21_1 ();
 FILLCELL_X1 FILLER_21_3 ();
 FILLCELL_X8 FILLER_21_7 ();
 FILLCELL_X2 FILLER_21_15 ();
 FILLCELL_X1 FILLER_21_20 ();
 FILLCELL_X4 FILLER_21_38 ();
 FILLCELL_X2 FILLER_21_42 ();
 FILLCELL_X1 FILLER_21_44 ();
 FILLCELL_X1 FILLER_21_69 ();
 FILLCELL_X4 FILLER_21_110 ();
 FILLCELL_X2 FILLER_21_118 ();
 FILLCELL_X4 FILLER_21_125 ();
 FILLCELL_X2 FILLER_21_129 ();
 FILLCELL_X2 FILLER_21_144 ();
 FILLCELL_X8 FILLER_21_153 ();
 FILLCELL_X4 FILLER_21_161 ();
 FILLCELL_X1 FILLER_21_165 ();
 FILLCELL_X16 FILLER_21_169 ();
 FILLCELL_X2 FILLER_21_185 ();
 FILLCELL_X1 FILLER_21_187 ();
 FILLCELL_X1 FILLER_21_192 ();
 FILLCELL_X4 FILLER_21_197 ();
 FILLCELL_X2 FILLER_21_201 ();
 FILLCELL_X1 FILLER_21_203 ();
 FILLCELL_X1 FILLER_21_219 ();
 FILLCELL_X1 FILLER_21_224 ();
 FILLCELL_X1 FILLER_21_229 ();
 FILLCELL_X4 FILLER_21_253 ();
 FILLCELL_X2 FILLER_21_257 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_17 ();
 FILLCELL_X1 FILLER_22_21 ();
 FILLCELL_X2 FILLER_22_25 ();
 FILLCELL_X8 FILLER_22_37 ();
 FILLCELL_X4 FILLER_22_45 ();
 FILLCELL_X2 FILLER_22_49 ();
 FILLCELL_X1 FILLER_22_51 ();
 FILLCELL_X1 FILLER_22_65 ();
 FILLCELL_X1 FILLER_22_71 ();
 FILLCELL_X1 FILLER_22_123 ();
 FILLCELL_X4 FILLER_22_132 ();
 FILLCELL_X2 FILLER_22_140 ();
 FILLCELL_X1 FILLER_22_142 ();
 FILLCELL_X8 FILLER_22_161 ();
 FILLCELL_X2 FILLER_22_169 ();
 FILLCELL_X2 FILLER_22_228 ();
 FILLCELL_X2 FILLER_22_233 ();
 FILLCELL_X2 FILLER_22_239 ();
 FILLCELL_X8 FILLER_22_247 ();
 FILLCELL_X4 FILLER_22_255 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X1 FILLER_23_5 ();
 FILLCELL_X4 FILLER_23_34 ();
 FILLCELL_X1 FILLER_23_38 ();
 FILLCELL_X2 FILLER_23_43 ();
 FILLCELL_X4 FILLER_23_48 ();
 FILLCELL_X8 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_94 ();
 FILLCELL_X1 FILLER_23_110 ();
 FILLCELL_X2 FILLER_23_119 ();
 FILLCELL_X2 FILLER_23_152 ();
 FILLCELL_X2 FILLER_23_164 ();
 FILLCELL_X2 FILLER_23_189 ();
 FILLCELL_X8 FILLER_23_211 ();
 FILLCELL_X1 FILLER_23_219 ();
 FILLCELL_X2 FILLER_23_223 ();
 FILLCELL_X1 FILLER_23_225 ();
 FILLCELL_X16 FILLER_23_233 ();
 FILLCELL_X8 FILLER_23_249 ();
 FILLCELL_X2 FILLER_23_257 ();
 FILLCELL_X4 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_5 ();
 FILLCELL_X1 FILLER_24_7 ();
 FILLCELL_X1 FILLER_24_32 ();
 FILLCELL_X2 FILLER_24_67 ();
 FILLCELL_X16 FILLER_24_86 ();
 FILLCELL_X4 FILLER_24_102 ();
 FILLCELL_X1 FILLER_24_106 ();
 FILLCELL_X1 FILLER_24_143 ();
 FILLCELL_X8 FILLER_24_209 ();
 FILLCELL_X1 FILLER_24_217 ();
 FILLCELL_X16 FILLER_24_235 ();
 FILLCELL_X8 FILLER_24_251 ();
 FILLCELL_X4 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_5 ();
 FILLCELL_X1 FILLER_25_17 ();
 FILLCELL_X8 FILLER_25_30 ();
 FILLCELL_X2 FILLER_25_38 ();
 FILLCELL_X8 FILLER_25_46 ();
 FILLCELL_X4 FILLER_25_61 ();
 FILLCELL_X1 FILLER_25_65 ();
 FILLCELL_X2 FILLER_25_90 ();
 FILLCELL_X1 FILLER_25_96 ();
 FILLCELL_X8 FILLER_25_101 ();
 FILLCELL_X2 FILLER_25_109 ();
 FILLCELL_X8 FILLER_25_120 ();
 FILLCELL_X4 FILLER_25_132 ();
 FILLCELL_X1 FILLER_25_136 ();
 FILLCELL_X4 FILLER_25_140 ();
 FILLCELL_X8 FILLER_25_149 ();
 FILLCELL_X4 FILLER_25_157 ();
 FILLCELL_X1 FILLER_25_173 ();
 FILLCELL_X1 FILLER_25_178 ();
 FILLCELL_X16 FILLER_25_183 ();
 FILLCELL_X8 FILLER_25_199 ();
 FILLCELL_X2 FILLER_25_207 ();
 FILLCELL_X1 FILLER_25_209 ();
 FILLCELL_X16 FILLER_25_236 ();
 FILLCELL_X4 FILLER_25_252 ();
 FILLCELL_X2 FILLER_25_256 ();
 FILLCELL_X1 FILLER_25_258 ();
 FILLCELL_X1 FILLER_26_24 ();
 FILLCELL_X8 FILLER_26_32 ();
 FILLCELL_X1 FILLER_26_40 ();
 FILLCELL_X32 FILLER_26_48 ();
 FILLCELL_X8 FILLER_26_80 ();
 FILLCELL_X2 FILLER_26_119 ();
 FILLCELL_X16 FILLER_26_131 ();
 FILLCELL_X2 FILLER_26_147 ();
 FILLCELL_X16 FILLER_26_177 ();
 FILLCELL_X2 FILLER_26_202 ();
 FILLCELL_X2 FILLER_26_224 ();
 FILLCELL_X1 FILLER_26_226 ();
 FILLCELL_X16 FILLER_26_231 ();
 FILLCELL_X8 FILLER_26_247 ();
 FILLCELL_X4 FILLER_26_255 ();
 FILLCELL_X2 FILLER_27_1 ();
 FILLCELL_X1 FILLER_27_3 ();
 FILLCELL_X2 FILLER_27_7 ();
 FILLCELL_X8 FILLER_27_33 ();
 FILLCELL_X2 FILLER_27_41 ();
 FILLCELL_X16 FILLER_27_60 ();
 FILLCELL_X2 FILLER_27_76 ();
 FILLCELL_X1 FILLER_27_78 ();
 FILLCELL_X16 FILLER_27_90 ();
 FILLCELL_X2 FILLER_27_151 ();
 FILLCELL_X4 FILLER_27_158 ();
 FILLCELL_X2 FILLER_27_168 ();
 FILLCELL_X16 FILLER_27_186 ();
 FILLCELL_X32 FILLER_27_206 ();
 FILLCELL_X16 FILLER_27_238 ();
 FILLCELL_X4 FILLER_27_254 ();
 FILLCELL_X1 FILLER_27_258 ();
 FILLCELL_X4 FILLER_28_1 ();
 FILLCELL_X1 FILLER_28_5 ();
 FILLCELL_X32 FILLER_28_23 ();
 FILLCELL_X8 FILLER_28_55 ();
 FILLCELL_X4 FILLER_28_63 ();
 FILLCELL_X16 FILLER_28_97 ();
 FILLCELL_X2 FILLER_28_113 ();
 FILLCELL_X1 FILLER_28_115 ();
 FILLCELL_X1 FILLER_28_160 ();
 FILLCELL_X2 FILLER_28_182 ();
 FILLCELL_X16 FILLER_28_187 ();
 FILLCELL_X32 FILLER_28_223 ();
 FILLCELL_X4 FILLER_28_255 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X8 FILLER_29_69 ();
 FILLCELL_X4 FILLER_29_77 ();
 FILLCELL_X1 FILLER_29_81 ();
 FILLCELL_X8 FILLER_29_90 ();
 FILLCELL_X4 FILLER_29_98 ();
 FILLCELL_X2 FILLER_29_102 ();
 FILLCELL_X1 FILLER_29_104 ();
 FILLCELL_X1 FILLER_29_122 ();
 FILLCELL_X8 FILLER_29_127 ();
 FILLCELL_X1 FILLER_29_135 ();
 FILLCELL_X2 FILLER_29_138 ();
 FILLCELL_X1 FILLER_29_153 ();
 FILLCELL_X32 FILLER_29_199 ();
 FILLCELL_X16 FILLER_29_231 ();
 FILLCELL_X8 FILLER_29_247 ();
 FILLCELL_X4 FILLER_29_255 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X16 FILLER_30_33 ();
 FILLCELL_X8 FILLER_30_49 ();
 FILLCELL_X4 FILLER_30_57 ();
 FILLCELL_X2 FILLER_30_61 ();
 FILLCELL_X1 FILLER_30_63 ();
 FILLCELL_X4 FILLER_30_81 ();
 FILLCELL_X2 FILLER_30_85 ();
 FILLCELL_X1 FILLER_30_87 ();
 FILLCELL_X32 FILLER_30_105 ();
 FILLCELL_X16 FILLER_30_151 ();
 FILLCELL_X4 FILLER_30_167 ();
 FILLCELL_X1 FILLER_30_171 ();
 FILLCELL_X32 FILLER_30_189 ();
 FILLCELL_X32 FILLER_30_221 ();
 FILLCELL_X4 FILLER_30_253 ();
 FILLCELL_X2 FILLER_30_257 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X8 FILLER_31_65 ();
 FILLCELL_X2 FILLER_31_73 ();
 FILLCELL_X1 FILLER_31_75 ();
 FILLCELL_X1 FILLER_31_78 ();
 FILLCELL_X1 FILLER_31_82 ();
 FILLCELL_X32 FILLER_31_100 ();
 FILLCELL_X32 FILLER_31_132 ();
 FILLCELL_X32 FILLER_31_164 ();
 FILLCELL_X32 FILLER_31_196 ();
 FILLCELL_X16 FILLER_31_228 ();
 FILLCELL_X8 FILLER_31_244 ();
 FILLCELL_X4 FILLER_31_252 ();
 FILLCELL_X2 FILLER_31_256 ();
 FILLCELL_X1 FILLER_31_258 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X2 FILLER_32_257 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X2 FILLER_33_257 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X16 FILLER_34_33 ();
 FILLCELL_X8 FILLER_34_49 ();
 FILLCELL_X4 FILLER_34_57 ();
 FILLCELL_X2 FILLER_34_61 ();
 FILLCELL_X1 FILLER_34_63 ();
 FILLCELL_X4 FILLER_34_67 ();
 FILLCELL_X2 FILLER_34_71 ();
 FILLCELL_X1 FILLER_34_73 ();
 FILLCELL_X2 FILLER_34_77 ();
 FILLCELL_X1 FILLER_34_79 ();
 FILLCELL_X8 FILLER_34_83 ();
 FILLCELL_X4 FILLER_34_91 ();
 FILLCELL_X4 FILLER_34_98 ();
 FILLCELL_X1 FILLER_34_102 ();
 FILLCELL_X32 FILLER_34_106 ();
 FILLCELL_X16 FILLER_34_138 ();
 FILLCELL_X8 FILLER_34_154 ();
 FILLCELL_X4 FILLER_34_162 ();
 FILLCELL_X32 FILLER_34_169 ();
 FILLCELL_X32 FILLER_34_201 ();
 FILLCELL_X16 FILLER_34_233 ();
 FILLCELL_X8 FILLER_34_249 ();
 FILLCELL_X2 FILLER_34_257 ();
endmodule
