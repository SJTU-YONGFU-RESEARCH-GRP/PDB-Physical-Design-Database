module configurable_priority_encoder (valid,
    grant_index,
    request);
 output valid;
 output [2:0] grant_index;
 input [7:0] request;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;

 INV_X1 _12_ (.A(net1),
    .ZN(_00_));
 NAND2_X1 _13_ (.A1(_00_),
    .A2(net2),
    .ZN(_01_));
 NAND2_X1 _14_ (.A1(_00_),
    .A2(net4),
    .ZN(_02_));
 INV_X1 _15_ (.A(net7),
    .ZN(_03_));
 AOI21_X1 _16_ (.A(net6),
    .B1(net8),
    .B2(_03_),
    .ZN(_04_));
 OR3_X1 _17_ (.A1(net1),
    .A2(net5),
    .A3(net3),
    .ZN(_05_));
 OAI221_X2 _18_ (.A(_01_),
    .B1(_02_),
    .B2(net3),
    .C1(_04_),
    .C2(_05_),
    .ZN(net9));
 OR2_X1 _19_ (.A1(net1),
    .A2(net2),
    .ZN(_06_));
 NOR2_X1 _20_ (.A1(net4),
    .A2(net3),
    .ZN(_07_));
 NOR2_X1 _21_ (.A1(net6),
    .A2(net5),
    .ZN(_08_));
 OAI21_X1 _22_ (.A(_08_),
    .B1(net8),
    .B2(net7),
    .ZN(_09_));
 AOI21_X1 _23_ (.A(_06_),
    .B1(_07_),
    .B2(_09_),
    .ZN(net10));
 NOR4_X2 _24_ (.A1(net7),
    .A2(net8),
    .A3(net6),
    .A4(net5),
    .ZN(_10_));
 NOR4_X2 _25_ (.A1(net4),
    .A2(net3),
    .A3(_06_),
    .A4(_10_),
    .ZN(net11));
 NOR2_X1 _26_ (.A1(net1),
    .A2(net2),
    .ZN(_11_));
 NAND3_X1 _27_ (.A1(_11_),
    .A2(_07_),
    .A3(_10_),
    .ZN(net12));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_83 ();
 BUF_X1 input1 (.A(request[0]),
    .Z(net1));
 BUF_X1 input2 (.A(request[1]),
    .Z(net2));
 CLKBUF_X2 input3 (.A(request[2]),
    .Z(net3));
 BUF_X1 input4 (.A(request[3]),
    .Z(net4));
 BUF_X1 input5 (.A(request[4]),
    .Z(net5));
 BUF_X1 input6 (.A(request[5]),
    .Z(net6));
 BUF_X1 input7 (.A(request[6]),
    .Z(net7));
 BUF_X1 input8 (.A(request[7]),
    .Z(net8));
 BUF_X1 output9 (.A(net9),
    .Z(grant_index[0]));
 BUF_X1 output10 (.A(net10),
    .Z(grant_index[1]));
 BUF_X1 output11 (.A(net11),
    .Z(grant_index[2]));
 BUF_X1 output12 (.A(net12),
    .Z(valid));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X16 FILLER_0_289 ();
 FILLCELL_X8 FILLER_0_305 ();
 FILLCELL_X1 FILLER_0_313 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X16 FILLER_1_289 ();
 FILLCELL_X8 FILLER_1_305 ();
 FILLCELL_X1 FILLER_1_313 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X16 FILLER_2_289 ();
 FILLCELL_X8 FILLER_2_305 ();
 FILLCELL_X1 FILLER_2_313 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X16 FILLER_3_289 ();
 FILLCELL_X8 FILLER_3_305 ();
 FILLCELL_X1 FILLER_3_313 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X16 FILLER_4_289 ();
 FILLCELL_X8 FILLER_4_305 ();
 FILLCELL_X1 FILLER_4_313 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X16 FILLER_5_289 ();
 FILLCELL_X8 FILLER_5_305 ();
 FILLCELL_X1 FILLER_5_313 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X16 FILLER_6_289 ();
 FILLCELL_X8 FILLER_6_305 ();
 FILLCELL_X1 FILLER_6_313 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X16 FILLER_7_289 ();
 FILLCELL_X8 FILLER_7_305 ();
 FILLCELL_X1 FILLER_7_313 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X16 FILLER_8_289 ();
 FILLCELL_X8 FILLER_8_305 ();
 FILLCELL_X1 FILLER_8_313 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X16 FILLER_9_289 ();
 FILLCELL_X8 FILLER_9_305 ();
 FILLCELL_X1 FILLER_9_313 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X16 FILLER_10_289 ();
 FILLCELL_X8 FILLER_10_305 ();
 FILLCELL_X1 FILLER_10_313 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X16 FILLER_11_289 ();
 FILLCELL_X8 FILLER_11_305 ();
 FILLCELL_X1 FILLER_11_313 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X16 FILLER_12_289 ();
 FILLCELL_X8 FILLER_12_305 ();
 FILLCELL_X1 FILLER_12_313 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X16 FILLER_13_289 ();
 FILLCELL_X8 FILLER_13_305 ();
 FILLCELL_X1 FILLER_13_313 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X16 FILLER_14_289 ();
 FILLCELL_X8 FILLER_14_305 ();
 FILLCELL_X1 FILLER_14_313 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X16 FILLER_15_289 ();
 FILLCELL_X8 FILLER_15_305 ();
 FILLCELL_X1 FILLER_15_313 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X16 FILLER_16_289 ();
 FILLCELL_X8 FILLER_16_305 ();
 FILLCELL_X1 FILLER_16_313 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X16 FILLER_17_289 ();
 FILLCELL_X8 FILLER_17_305 ();
 FILLCELL_X1 FILLER_17_313 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X16 FILLER_18_289 ();
 FILLCELL_X8 FILLER_18_305 ();
 FILLCELL_X1 FILLER_18_313 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X16 FILLER_19_289 ();
 FILLCELL_X8 FILLER_19_305 ();
 FILLCELL_X1 FILLER_19_313 ();
 FILLCELL_X16 FILLER_20_4 ();
 FILLCELL_X8 FILLER_20_20 ();
 FILLCELL_X4 FILLER_20_28 ();
 FILLCELL_X32 FILLER_20_35 ();
 FILLCELL_X32 FILLER_20_67 ();
 FILLCELL_X16 FILLER_20_99 ();
 FILLCELL_X8 FILLER_20_115 ();
 FILLCELL_X4 FILLER_20_123 ();
 FILLCELL_X1 FILLER_20_127 ();
 FILLCELL_X16 FILLER_20_131 ();
 FILLCELL_X8 FILLER_20_147 ();
 FILLCELL_X4 FILLER_20_159 ();
 FILLCELL_X32 FILLER_20_171 ();
 FILLCELL_X32 FILLER_20_203 ();
 FILLCELL_X32 FILLER_20_235 ();
 FILLCELL_X8 FILLER_20_267 ();
 FILLCELL_X2 FILLER_20_275 ();
 FILLCELL_X1 FILLER_20_277 ();
 FILLCELL_X1 FILLER_20_281 ();
 FILLCELL_X16 FILLER_20_285 ();
 FILLCELL_X8 FILLER_20_301 ();
 FILLCELL_X4 FILLER_20_309 ();
 FILLCELL_X1 FILLER_20_313 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X1 FILLER_21_9 ();
 FILLCELL_X2 FILLER_21_13 ();
 FILLCELL_X16 FILLER_21_18 ();
 FILLCELL_X1 FILLER_21_34 ();
 FILLCELL_X32 FILLER_21_38 ();
 FILLCELL_X32 FILLER_21_70 ();
 FILLCELL_X16 FILLER_21_102 ();
 FILLCELL_X1 FILLER_21_118 ();
 FILLCELL_X2 FILLER_21_138 ();
 FILLCELL_X1 FILLER_21_140 ();
 FILLCELL_X32 FILLER_21_173 ();
 FILLCELL_X32 FILLER_21_205 ();
 FILLCELL_X32 FILLER_21_237 ();
 FILLCELL_X8 FILLER_21_269 ();
 FILLCELL_X1 FILLER_21_280 ();
 FILLCELL_X16 FILLER_21_284 ();
 FILLCELL_X8 FILLER_21_300 ();
 FILLCELL_X4 FILLER_21_308 ();
 FILLCELL_X2 FILLER_21_312 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X16 FILLER_22_129 ();
 FILLCELL_X4 FILLER_22_145 ();
 FILLCELL_X2 FILLER_22_149 ();
 FILLCELL_X32 FILLER_22_158 ();
 FILLCELL_X32 FILLER_22_190 ();
 FILLCELL_X32 FILLER_22_222 ();
 FILLCELL_X32 FILLER_22_254 ();
 FILLCELL_X16 FILLER_22_286 ();
 FILLCELL_X8 FILLER_22_302 ();
 FILLCELL_X4 FILLER_22_310 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X16 FILLER_23_289 ();
 FILLCELL_X8 FILLER_23_305 ();
 FILLCELL_X1 FILLER_23_313 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X16 FILLER_24_289 ();
 FILLCELL_X8 FILLER_24_305 ();
 FILLCELL_X1 FILLER_24_313 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X16 FILLER_25_289 ();
 FILLCELL_X8 FILLER_25_305 ();
 FILLCELL_X1 FILLER_25_313 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X16 FILLER_26_289 ();
 FILLCELL_X8 FILLER_26_305 ();
 FILLCELL_X1 FILLER_26_313 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X16 FILLER_27_289 ();
 FILLCELL_X8 FILLER_27_305 ();
 FILLCELL_X1 FILLER_27_313 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X16 FILLER_28_289 ();
 FILLCELL_X8 FILLER_28_305 ();
 FILLCELL_X1 FILLER_28_313 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X16 FILLER_29_289 ();
 FILLCELL_X8 FILLER_29_305 ();
 FILLCELL_X1 FILLER_29_313 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X16 FILLER_30_289 ();
 FILLCELL_X8 FILLER_30_305 ();
 FILLCELL_X1 FILLER_30_313 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X16 FILLER_31_289 ();
 FILLCELL_X8 FILLER_31_305 ();
 FILLCELL_X1 FILLER_31_313 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X16 FILLER_32_289 ();
 FILLCELL_X8 FILLER_32_305 ();
 FILLCELL_X1 FILLER_32_313 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X16 FILLER_33_289 ();
 FILLCELL_X8 FILLER_33_305 ();
 FILLCELL_X1 FILLER_33_313 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X16 FILLER_34_289 ();
 FILLCELL_X8 FILLER_34_305 ();
 FILLCELL_X1 FILLER_34_313 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X16 FILLER_35_289 ();
 FILLCELL_X8 FILLER_35_305 ();
 FILLCELL_X1 FILLER_35_313 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X16 FILLER_36_289 ();
 FILLCELL_X8 FILLER_36_305 ();
 FILLCELL_X1 FILLER_36_313 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X16 FILLER_37_289 ();
 FILLCELL_X8 FILLER_37_305 ();
 FILLCELL_X1 FILLER_37_313 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X16 FILLER_38_289 ();
 FILLCELL_X8 FILLER_38_305 ();
 FILLCELL_X1 FILLER_38_313 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X16 FILLER_39_289 ();
 FILLCELL_X8 FILLER_39_305 ();
 FILLCELL_X1 FILLER_39_313 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X16 FILLER_40_289 ();
 FILLCELL_X8 FILLER_40_305 ();
 FILLCELL_X1 FILLER_40_313 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X16 FILLER_41_129 ();
 FILLCELL_X8 FILLER_41_145 ();
 FILLCELL_X1 FILLER_41_153 ();
 FILLCELL_X2 FILLER_41_160 ();
 FILLCELL_X32 FILLER_41_166 ();
 FILLCELL_X32 FILLER_41_198 ();
 FILLCELL_X32 FILLER_41_230 ();
 FILLCELL_X32 FILLER_41_262 ();
 FILLCELL_X16 FILLER_41_294 ();
 FILLCELL_X4 FILLER_41_310 ();
endmodule
