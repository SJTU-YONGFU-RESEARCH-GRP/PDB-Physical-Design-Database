module scan_register (clk,
    rst_n,
    scan_en,
    scan_in,
    scan_out,
    data_in,
    data_out);
 input clk;
 input rst_n;
 input scan_en;
 input scan_in;
 output scan_out;
 input [7:0] data_in;
 output [7:0] data_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire _37_;
 wire _38_;
 wire _39_;
 wire _40_;
 wire _41_;
 wire _42_;
 wire _43_;
 wire _44_;
 wire _45_;
 wire _46_;
 wire _47_;
 wire _48_;
 wire _49_;
 wire _50_;
 wire _51_;
 wire \scan_reg[0] ;
 wire \scan_reg[1] ;
 wire \scan_reg[2] ;
 wire \scan_reg[3] ;
 wire \scan_reg[4] ;
 wire \scan_reg[5] ;
 wire \scan_reg[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X1 _52_ (.A(rst_n),
    .Z(_16_));
 BUF_X2 _53_ (.A(_16_),
    .Z(_17_));
 BUF_X4 _54_ (.A(scan_en),
    .Z(_18_));
 BUF_X8 _55_ (.A(_18_),
    .Z(_19_));
 MUX2_X1 _56_ (.A(\scan_reg[0] ),
    .B(net9),
    .S(_19_),
    .Z(_20_));
 AND2_X1 _57_ (.A1(_17_),
    .A2(_20_),
    .ZN(_00_));
 MUX2_X1 _58_ (.A(\scan_reg[1] ),
    .B(\scan_reg[0] ),
    .S(_19_),
    .Z(_21_));
 AND2_X1 _59_ (.A1(_17_),
    .A2(_21_),
    .ZN(_01_));
 MUX2_X1 _60_ (.A(\scan_reg[2] ),
    .B(\scan_reg[1] ),
    .S(_19_),
    .Z(_22_));
 AND2_X1 _61_ (.A1(_17_),
    .A2(_22_),
    .ZN(_02_));
 MUX2_X1 _62_ (.A(\scan_reg[3] ),
    .B(\scan_reg[2] ),
    .S(_19_),
    .Z(_23_));
 AND2_X1 _63_ (.A1(_17_),
    .A2(_23_),
    .ZN(_03_));
 MUX2_X1 _64_ (.A(\scan_reg[4] ),
    .B(\scan_reg[3] ),
    .S(_19_),
    .Z(_24_));
 AND2_X1 _65_ (.A1(_17_),
    .A2(_24_),
    .ZN(_04_));
 MUX2_X1 _66_ (.A(\scan_reg[5] ),
    .B(\scan_reg[4] ),
    .S(_19_),
    .Z(_25_));
 AND2_X1 _67_ (.A1(_17_),
    .A2(_25_),
    .ZN(_05_));
 MUX2_X1 _68_ (.A(\scan_reg[6] ),
    .B(\scan_reg[5] ),
    .S(_19_),
    .Z(_26_));
 AND2_X1 _69_ (.A1(_17_),
    .A2(_26_),
    .ZN(_06_));
 MUX2_X1 _70_ (.A(net18),
    .B(\scan_reg[6] ),
    .S(_19_),
    .Z(_27_));
 AND2_X1 _71_ (.A1(_17_),
    .A2(_27_),
    .ZN(_07_));
 MUX2_X1 _72_ (.A(net1),
    .B(net9),
    .S(_19_),
    .Z(_28_));
 AND2_X1 _73_ (.A1(_17_),
    .A2(_28_),
    .ZN(_08_));
 MUX2_X1 _74_ (.A(net2),
    .B(\scan_reg[0] ),
    .S(_19_),
    .Z(_29_));
 AND2_X1 _75_ (.A1(_17_),
    .A2(_29_),
    .ZN(_09_));
 MUX2_X1 _76_ (.A(net3),
    .B(\scan_reg[1] ),
    .S(_18_),
    .Z(_30_));
 AND2_X1 _77_ (.A1(_16_),
    .A2(_30_),
    .ZN(_10_));
 MUX2_X1 _78_ (.A(net4),
    .B(\scan_reg[2] ),
    .S(_18_),
    .Z(_31_));
 AND2_X1 _79_ (.A1(_16_),
    .A2(_31_),
    .ZN(_11_));
 MUX2_X1 _80_ (.A(net5),
    .B(\scan_reg[3] ),
    .S(_18_),
    .Z(_32_));
 AND2_X1 _81_ (.A1(_16_),
    .A2(_32_),
    .ZN(_12_));
 MUX2_X1 _82_ (.A(net6),
    .B(\scan_reg[4] ),
    .S(_18_),
    .Z(_33_));
 AND2_X1 _83_ (.A1(_16_),
    .A2(_33_),
    .ZN(_13_));
 MUX2_X1 _84_ (.A(net7),
    .B(\scan_reg[5] ),
    .S(_18_),
    .Z(_34_));
 AND2_X1 _85_ (.A1(_16_),
    .A2(_34_),
    .ZN(_14_));
 MUX2_X1 _86_ (.A(net8),
    .B(\scan_reg[6] ),
    .S(_18_),
    .Z(_35_));
 AND2_X1 _87_ (.A1(_16_),
    .A2(_35_),
    .ZN(_15_));
 DFF_X1 \data_out[0]$_SDFF_PN0_  (.D(_00_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net10),
    .QN(_51_));
 DFF_X1 \data_out[1]$_SDFF_PN0_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net11),
    .QN(_50_));
 DFF_X1 \data_out[2]$_SDFF_PN0_  (.D(_02_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net12),
    .QN(_49_));
 DFF_X1 \data_out[3]$_SDFF_PN0_  (.D(_03_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net13),
    .QN(_48_));
 DFF_X1 \data_out[4]$_SDFF_PN0_  (.D(_04_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net14),
    .QN(_47_));
 DFF_X1 \data_out[5]$_SDFF_PN0_  (.D(_05_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net15),
    .QN(_46_));
 DFF_X1 \data_out[6]$_SDFF_PN0_  (.D(_06_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net16),
    .QN(_45_));
 DFF_X1 \data_out[7]$_SDFF_PN0_  (.D(_07_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net17),
    .QN(_44_));
 DFF_X1 \scan_reg[0]$_SDFF_PN0_  (.D(_08_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\scan_reg[0] ),
    .QN(_43_));
 DFF_X1 \scan_reg[1]$_SDFF_PN0_  (.D(_09_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\scan_reg[1] ),
    .QN(_42_));
 DFF_X1 \scan_reg[2]$_SDFF_PN0_  (.D(_10_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\scan_reg[2] ),
    .QN(_41_));
 DFF_X1 \scan_reg[3]$_SDFF_PN0_  (.D(_11_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\scan_reg[3] ),
    .QN(_40_));
 DFF_X1 \scan_reg[4]$_SDFF_PN0_  (.D(_12_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\scan_reg[4] ),
    .QN(_39_));
 DFF_X1 \scan_reg[5]$_SDFF_PN0_  (.D(_13_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\scan_reg[5] ),
    .QN(_38_));
 DFF_X1 \scan_reg[6]$_SDFF_PN0_  (.D(_14_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\scan_reg[6] ),
    .QN(_37_));
 DFF_X1 \scan_reg[7]$_SDFF_PN0_  (.D(_15_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net18),
    .QN(_36_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_71 ();
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[2]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[3]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[5]),
    .Z(net6));
 BUF_X1 input7 (.A(data_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[7]),
    .Z(net8));
 BUF_X1 input9 (.A(scan_in),
    .Z(net9));
 BUF_X1 output10 (.A(net10),
    .Z(data_out[0]));
 BUF_X1 output11 (.A(net11),
    .Z(data_out[1]));
 BUF_X1 output12 (.A(net12),
    .Z(data_out[2]));
 BUF_X1 output13 (.A(net13),
    .Z(data_out[3]));
 BUF_X1 output14 (.A(net14),
    .Z(data_out[4]));
 BUF_X1 output15 (.A(net15),
    .Z(data_out[5]));
 BUF_X1 output16 (.A(net16),
    .Z(data_out[6]));
 BUF_X1 output17 (.A(net17),
    .Z(data_out[7]));
 BUF_X1 output18 (.A(net18),
    .Z(scan_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 INV_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X16 FILLER_0_97 ();
 FILLCELL_X1 FILLER_0_113 ();
 FILLCELL_X4 FILLER_0_117 ();
 FILLCELL_X2 FILLER_0_121 ();
 FILLCELL_X1 FILLER_0_123 ();
 FILLCELL_X8 FILLER_0_127 ();
 FILLCELL_X4 FILLER_0_135 ();
 FILLCELL_X2 FILLER_0_139 ();
 FILLCELL_X1 FILLER_0_144 ();
 FILLCELL_X16 FILLER_0_148 ();
 FILLCELL_X8 FILLER_0_164 ();
 FILLCELL_X2 FILLER_0_172 ();
 FILLCELL_X32 FILLER_0_177 ();
 FILLCELL_X32 FILLER_0_209 ();
 FILLCELL_X16 FILLER_0_241 ();
 FILLCELL_X8 FILLER_0_257 ();
 FILLCELL_X2 FILLER_0_265 ();
 FILLCELL_X1 FILLER_0_267 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X8 FILLER_1_257 ();
 FILLCELL_X2 FILLER_1_265 ();
 FILLCELL_X1 FILLER_1_267 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X8 FILLER_2_257 ();
 FILLCELL_X2 FILLER_2_265 ();
 FILLCELL_X1 FILLER_2_267 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X8 FILLER_3_257 ();
 FILLCELL_X2 FILLER_3_265 ();
 FILLCELL_X1 FILLER_3_267 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X8 FILLER_4_257 ();
 FILLCELL_X2 FILLER_4_265 ();
 FILLCELL_X1 FILLER_4_267 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X8 FILLER_5_257 ();
 FILLCELL_X2 FILLER_5_265 ();
 FILLCELL_X1 FILLER_5_267 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X8 FILLER_6_257 ();
 FILLCELL_X2 FILLER_6_265 ();
 FILLCELL_X1 FILLER_6_267 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X8 FILLER_7_257 ();
 FILLCELL_X2 FILLER_7_265 ();
 FILLCELL_X1 FILLER_7_267 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X8 FILLER_8_129 ();
 FILLCELL_X4 FILLER_8_137 ();
 FILLCELL_X2 FILLER_8_141 ();
 FILLCELL_X8 FILLER_8_150 ();
 FILLCELL_X32 FILLER_8_175 ();
 FILLCELL_X32 FILLER_8_207 ();
 FILLCELL_X16 FILLER_8_239 ();
 FILLCELL_X8 FILLER_8_255 ();
 FILLCELL_X4 FILLER_8_263 ();
 FILLCELL_X1 FILLER_8_267 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X16 FILLER_9_97 ();
 FILLCELL_X8 FILLER_9_113 ();
 FILLCELL_X2 FILLER_9_121 ();
 FILLCELL_X1 FILLER_9_123 ();
 FILLCELL_X32 FILLER_9_156 ();
 FILLCELL_X32 FILLER_9_188 ();
 FILLCELL_X32 FILLER_9_220 ();
 FILLCELL_X16 FILLER_9_252 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X16 FILLER_10_97 ();
 FILLCELL_X8 FILLER_10_113 ();
 FILLCELL_X4 FILLER_10_121 ();
 FILLCELL_X32 FILLER_10_132 ();
 FILLCELL_X32 FILLER_10_164 ();
 FILLCELL_X32 FILLER_10_196 ();
 FILLCELL_X32 FILLER_10_228 ();
 FILLCELL_X8 FILLER_10_260 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X16 FILLER_11_97 ();
 FILLCELL_X8 FILLER_11_113 ();
 FILLCELL_X2 FILLER_11_121 ();
 FILLCELL_X1 FILLER_11_123 ();
 FILLCELL_X8 FILLER_11_128 ();
 FILLCELL_X4 FILLER_11_136 ();
 FILLCELL_X1 FILLER_11_140 ();
 FILLCELL_X32 FILLER_11_148 ();
 FILLCELL_X32 FILLER_11_180 ();
 FILLCELL_X32 FILLER_11_212 ();
 FILLCELL_X16 FILLER_11_244 ();
 FILLCELL_X8 FILLER_11_260 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X8 FILLER_12_113 ();
 FILLCELL_X1 FILLER_12_121 ();
 FILLCELL_X8 FILLER_12_139 ();
 FILLCELL_X4 FILLER_12_147 ();
 FILLCELL_X32 FILLER_12_155 ();
 FILLCELL_X32 FILLER_12_187 ();
 FILLCELL_X32 FILLER_12_219 ();
 FILLCELL_X16 FILLER_12_251 ();
 FILLCELL_X1 FILLER_12_267 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X16 FILLER_13_129 ();
 FILLCELL_X8 FILLER_13_145 ();
 FILLCELL_X4 FILLER_13_153 ();
 FILLCELL_X32 FILLER_13_174 ();
 FILLCELL_X32 FILLER_13_206 ();
 FILLCELL_X16 FILLER_13_238 ();
 FILLCELL_X8 FILLER_13_254 ();
 FILLCELL_X2 FILLER_13_265 ();
 FILLCELL_X1 FILLER_13_267 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X8 FILLER_14_33 ();
 FILLCELL_X4 FILLER_14_41 ();
 FILLCELL_X32 FILLER_14_52 ();
 FILLCELL_X16 FILLER_14_84 ();
 FILLCELL_X8 FILLER_14_100 ();
 FILLCELL_X4 FILLER_14_108 ();
 FILLCELL_X2 FILLER_14_112 ();
 FILLCELL_X16 FILLER_14_121 ();
 FILLCELL_X8 FILLER_14_137 ();
 FILLCELL_X2 FILLER_14_145 ();
 FILLCELL_X32 FILLER_14_154 ();
 FILLCELL_X32 FILLER_14_186 ();
 FILLCELL_X32 FILLER_14_218 ();
 FILLCELL_X16 FILLER_14_250 ();
 FILLCELL_X2 FILLER_14_266 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X16 FILLER_15_97 ();
 FILLCELL_X8 FILLER_15_113 ();
 FILLCELL_X4 FILLER_15_121 ();
 FILLCELL_X2 FILLER_15_125 ();
 FILLCELL_X1 FILLER_15_127 ();
 FILLCELL_X4 FILLER_15_133 ();
 FILLCELL_X1 FILLER_15_137 ();
 FILLCELL_X2 FILLER_15_145 ();
 FILLCELL_X32 FILLER_15_151 ();
 FILLCELL_X32 FILLER_15_183 ();
 FILLCELL_X32 FILLER_15_215 ();
 FILLCELL_X16 FILLER_15_247 ();
 FILLCELL_X4 FILLER_15_263 ();
 FILLCELL_X1 FILLER_15_267 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_17 ();
 FILLCELL_X1 FILLER_16_19 ();
 FILLCELL_X32 FILLER_16_23 ();
 FILLCELL_X16 FILLER_16_55 ();
 FILLCELL_X2 FILLER_16_71 ();
 FILLCELL_X32 FILLER_16_84 ();
 FILLCELL_X2 FILLER_16_116 ();
 FILLCELL_X1 FILLER_16_118 ();
 FILLCELL_X16 FILLER_16_140 ();
 FILLCELL_X4 FILLER_16_156 ();
 FILLCELL_X32 FILLER_16_177 ();
 FILLCELL_X16 FILLER_16_209 ();
 FILLCELL_X8 FILLER_16_225 ();
 FILLCELL_X2 FILLER_16_233 ();
 FILLCELL_X16 FILLER_16_238 ();
 FILLCELL_X8 FILLER_16_254 ();
 FILLCELL_X4 FILLER_16_262 ();
 FILLCELL_X2 FILLER_16_266 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X8 FILLER_17_33 ();
 FILLCELL_X4 FILLER_17_41 ();
 FILLCELL_X2 FILLER_17_45 ();
 FILLCELL_X1 FILLER_17_47 ();
 FILLCELL_X16 FILLER_17_51 ();
 FILLCELL_X8 FILLER_17_67 ();
 FILLCELL_X4 FILLER_17_75 ();
 FILLCELL_X32 FILLER_17_96 ();
 FILLCELL_X8 FILLER_17_128 ();
 FILLCELL_X1 FILLER_17_136 ();
 FILLCELL_X4 FILLER_17_144 ();
 FILLCELL_X2 FILLER_17_148 ();
 FILLCELL_X1 FILLER_17_150 ();
 FILLCELL_X4 FILLER_17_155 ();
 FILLCELL_X32 FILLER_17_176 ();
 FILLCELL_X16 FILLER_17_208 ();
 FILLCELL_X8 FILLER_17_224 ();
 FILLCELL_X2 FILLER_17_232 ();
 FILLCELL_X1 FILLER_17_234 ();
 FILLCELL_X16 FILLER_17_238 ();
 FILLCELL_X8 FILLER_17_254 ();
 FILLCELL_X4 FILLER_17_262 ();
 FILLCELL_X2 FILLER_17_266 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X8 FILLER_18_65 ();
 FILLCELL_X1 FILLER_18_73 ();
 FILLCELL_X32 FILLER_18_78 ();
 FILLCELL_X4 FILLER_18_110 ();
 FILLCELL_X1 FILLER_18_114 ();
 FILLCELL_X32 FILLER_18_128 ();
 FILLCELL_X32 FILLER_18_160 ();
 FILLCELL_X32 FILLER_18_192 ();
 FILLCELL_X32 FILLER_18_224 ();
 FILLCELL_X8 FILLER_18_256 ();
 FILLCELL_X4 FILLER_18_264 ();
 FILLCELL_X16 FILLER_19_1 ();
 FILLCELL_X8 FILLER_19_17 ();
 FILLCELL_X2 FILLER_19_25 ();
 FILLCELL_X1 FILLER_19_27 ();
 FILLCELL_X32 FILLER_19_31 ();
 FILLCELL_X4 FILLER_19_63 ();
 FILLCELL_X1 FILLER_19_67 ();
 FILLCELL_X1 FILLER_19_75 ();
 FILLCELL_X16 FILLER_19_93 ();
 FILLCELL_X8 FILLER_19_109 ();
 FILLCELL_X4 FILLER_19_117 ();
 FILLCELL_X32 FILLER_19_125 ();
 FILLCELL_X32 FILLER_19_157 ();
 FILLCELL_X32 FILLER_19_189 ();
 FILLCELL_X32 FILLER_19_221 ();
 FILLCELL_X8 FILLER_19_253 ();
 FILLCELL_X4 FILLER_19_261 ();
 FILLCELL_X2 FILLER_19_265 ();
 FILLCELL_X1 FILLER_19_267 ();
 FILLCELL_X16 FILLER_20_1 ();
 FILLCELL_X8 FILLER_20_17 ();
 FILLCELL_X2 FILLER_20_25 ();
 FILLCELL_X32 FILLER_20_30 ();
 FILLCELL_X8 FILLER_20_62 ();
 FILLCELL_X2 FILLER_20_70 ();
 FILLCELL_X1 FILLER_20_72 ();
 FILLCELL_X2 FILLER_20_80 ();
 FILLCELL_X1 FILLER_20_82 ();
 FILLCELL_X8 FILLER_20_87 ();
 FILLCELL_X2 FILLER_20_95 ();
 FILLCELL_X16 FILLER_20_108 ();
 FILLCELL_X4 FILLER_20_124 ();
 FILLCELL_X2 FILLER_20_128 ();
 FILLCELL_X4 FILLER_20_144 ();
 FILLCELL_X2 FILLER_20_148 ();
 FILLCELL_X8 FILLER_20_154 ();
 FILLCELL_X32 FILLER_20_179 ();
 FILLCELL_X16 FILLER_20_211 ();
 FILLCELL_X4 FILLER_20_227 ();
 FILLCELL_X32 FILLER_20_234 ();
 FILLCELL_X2 FILLER_20_266 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X16 FILLER_21_65 ();
 FILLCELL_X4 FILLER_21_81 ();
 FILLCELL_X2 FILLER_21_85 ();
 FILLCELL_X4 FILLER_21_121 ();
 FILLCELL_X2 FILLER_21_125 ();
 FILLCELL_X4 FILLER_21_132 ();
 FILLCELL_X2 FILLER_21_136 ();
 FILLCELL_X1 FILLER_21_138 ();
 FILLCELL_X32 FILLER_21_146 ();
 FILLCELL_X32 FILLER_21_178 ();
 FILLCELL_X32 FILLER_21_210 ();
 FILLCELL_X16 FILLER_21_242 ();
 FILLCELL_X8 FILLER_21_258 ();
 FILLCELL_X2 FILLER_21_266 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X16 FILLER_22_97 ();
 FILLCELL_X8 FILLER_22_124 ();
 FILLCELL_X2 FILLER_22_143 ();
 FILLCELL_X1 FILLER_22_145 ();
 FILLCELL_X1 FILLER_22_150 ();
 FILLCELL_X32 FILLER_22_155 ();
 FILLCELL_X32 FILLER_22_187 ();
 FILLCELL_X32 FILLER_22_219 ();
 FILLCELL_X16 FILLER_22_251 ();
 FILLCELL_X1 FILLER_22_267 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_97 ();
 FILLCELL_X4 FILLER_23_113 ();
 FILLCELL_X2 FILLER_23_117 ();
 FILLCELL_X16 FILLER_23_136 ();
 FILLCELL_X2 FILLER_23_152 ();
 FILLCELL_X1 FILLER_23_154 ();
 FILLCELL_X32 FILLER_23_172 ();
 FILLCELL_X32 FILLER_23_204 ();
 FILLCELL_X32 FILLER_23_236 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X1 FILLER_24_129 ();
 FILLCELL_X4 FILLER_24_147 ();
 FILLCELL_X32 FILLER_24_168 ();
 FILLCELL_X32 FILLER_24_200 ();
 FILLCELL_X32 FILLER_24_232 ();
 FILLCELL_X4 FILLER_24_264 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X8 FILLER_25_257 ();
 FILLCELL_X2 FILLER_25_265 ();
 FILLCELL_X1 FILLER_25_267 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X8 FILLER_26_257 ();
 FILLCELL_X2 FILLER_26_265 ();
 FILLCELL_X1 FILLER_26_267 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X8 FILLER_27_257 ();
 FILLCELL_X2 FILLER_27_265 ();
 FILLCELL_X1 FILLER_27_267 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X8 FILLER_28_257 ();
 FILLCELL_X2 FILLER_28_265 ();
 FILLCELL_X1 FILLER_28_267 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X8 FILLER_29_257 ();
 FILLCELL_X2 FILLER_29_265 ();
 FILLCELL_X1 FILLER_29_267 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X8 FILLER_30_257 ();
 FILLCELL_X2 FILLER_30_265 ();
 FILLCELL_X1 FILLER_30_267 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X8 FILLER_31_257 ();
 FILLCELL_X2 FILLER_31_265 ();
 FILLCELL_X1 FILLER_31_267 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X8 FILLER_32_257 ();
 FILLCELL_X2 FILLER_32_265 ();
 FILLCELL_X1 FILLER_32_267 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X8 FILLER_33_257 ();
 FILLCELL_X2 FILLER_33_265 ();
 FILLCELL_X1 FILLER_33_267 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X16 FILLER_34_65 ();
 FILLCELL_X8 FILLER_34_81 ();
 FILLCELL_X4 FILLER_34_89 ();
 FILLCELL_X2 FILLER_34_93 ();
 FILLCELL_X1 FILLER_34_95 ();
 FILLCELL_X32 FILLER_34_99 ();
 FILLCELL_X32 FILLER_34_131 ();
 FILLCELL_X32 FILLER_34_163 ();
 FILLCELL_X32 FILLER_34_195 ();
 FILLCELL_X32 FILLER_34_227 ();
 FILLCELL_X8 FILLER_34_259 ();
 FILLCELL_X1 FILLER_34_267 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X16 FILLER_35_97 ();
 FILLCELL_X2 FILLER_35_113 ();
 FILLCELL_X16 FILLER_35_118 ();
 FILLCELL_X2 FILLER_35_134 ();
 FILLCELL_X4 FILLER_35_139 ();
 FILLCELL_X2 FILLER_35_143 ();
 FILLCELL_X1 FILLER_35_145 ();
 FILLCELL_X16 FILLER_35_149 ();
 FILLCELL_X2 FILLER_35_165 ();
 FILLCELL_X1 FILLER_35_170 ();
 FILLCELL_X32 FILLER_35_174 ();
 FILLCELL_X32 FILLER_35_206 ();
 FILLCELL_X16 FILLER_35_238 ();
 FILLCELL_X8 FILLER_35_254 ();
 FILLCELL_X4 FILLER_35_262 ();
 FILLCELL_X2 FILLER_35_266 ();
endmodule
