module uart_rx (busy,
    clk,
    frame_error,
    m_axis_tready,
    m_axis_tvalid,
    overrun_error,
    rst,
    rxd,
    m_axis_tdata,
    prescale);
 output busy;
 input clk;
 output frame_error;
 input m_axis_tready;
 output m_axis_tvalid;
 output overrun_error;
 input rst;
 input rxd;
 output [7:0] m_axis_tdata;
 input [15:0] prescale;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire net16;
 wire _045_;
 wire net15;
 wire _047_;
 wire net14;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire net13;
 wire _065_;
 wire _066_;
 wire _067_;
 wire net12;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire net11;
 wire net10;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire net9;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire net8;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire net7;
 wire net6;
 wire net5;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire net4;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire net3;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire net2;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire net1;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire \bit_cnt[0] ;
 wire \bit_cnt[1] ;
 wire \bit_cnt[2] ;
 wire \bit_cnt[3] ;
 wire net20;
 wire \data_reg[0] ;
 wire \data_reg[1] ;
 wire \data_reg[2] ;
 wire \data_reg[3] ;
 wire \data_reg[4] ;
 wire \data_reg[5] ;
 wire \data_reg[6] ;
 wire \data_reg[7] ;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire \prescale_reg[0] ;
 wire \prescale_reg[10] ;
 wire \prescale_reg[11] ;
 wire \prescale_reg[12] ;
 wire \prescale_reg[13] ;
 wire \prescale_reg[14] ;
 wire \prescale_reg[15] ;
 wire \prescale_reg[16] ;
 wire \prescale_reg[17] ;
 wire \prescale_reg[18] ;
 wire \prescale_reg[1] ;
 wire \prescale_reg[2] ;
 wire \prescale_reg[3] ;
 wire \prescale_reg[4] ;
 wire \prescale_reg[5] ;
 wire \prescale_reg[6] ;
 wire \prescale_reg[7] ;
 wire \prescale_reg[8] ;
 wire \prescale_reg[9] ;
 wire rxd_reg;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire [0:0] _298_;
 wire [0:0] _299_;
 wire [0:0] _300_;
 wire [0:0] _301_;
 wire [0:0] _302_;
 wire [0:0] _303_;
 wire [0:0] _304_;
 wire [0:0] _305_;
 wire [0:0] _306_;
 wire [0:0] _307_;
 wire [0:0] _308_;
 wire [0:0] _309_;
 wire [0:0] _310_;
 wire [0:0] _311_;
 wire [0:0] _312_;
 wire [0:0] _313_;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _314_ (.I(\prescale_reg[0] ),
    .ZN(_304_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _315_ (.I(net2),
    .ZN(_310_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _316_ (.I(\bit_cnt[0] ),
    .ZN(_298_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _317_ (.I(\bit_cnt[1] ),
    .ZN(_299_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _318_ (.I(\prescale_reg[1] ),
    .ZN(_305_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _319_ (.I(net9),
    .ZN(_311_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input16 (.I(prescale[8]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _321_ (.A1(\bit_cnt[3] ),
    .A2(\bit_cnt[2] ),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input15 (.I(prescale[7]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _323_ (.A1(_300_[0]),
    .A2(_045_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input14 (.I(prescale[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _325_ (.A1(\data_reg[1] ),
    .A2(_047_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _326_ (.I0(_302_[0]),
    .I1(rxd_reg),
    .S(_300_[0]),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _327_ (.A1(_045_),
    .A2(_050_),
    .B(net18),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _328_ (.A1(_300_[0]),
    .A2(_302_[0]),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _329_ (.A1(\bit_cnt[2] ),
    .A2(_052_),
    .B(\bit_cnt[3] ),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _330_ (.A1(\prescale_reg[13] ),
    .A2(\prescale_reg[15] ),
    .A3(\prescale_reg[14] ),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _331_ (.A1(\prescale_reg[16] ),
    .A2(_054_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _332_ (.A1(\prescale_reg[1] ),
    .A2(\prescale_reg[0] ),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _333_ (.A1(\prescale_reg[4] ),
    .A2(\prescale_reg[3] ),
    .A3(\prescale_reg[2] ),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _334_ (.A1(\prescale_reg[5] ),
    .A2(\prescale_reg[8] ),
    .A3(\prescale_reg[7] ),
    .A4(\prescale_reg[6] ),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _335_ (.A1(\prescale_reg[12] ),
    .A2(\prescale_reg[11] ),
    .A3(\prescale_reg[10] ),
    .A4(\prescale_reg[9] ),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _336_ (.A1(_056_),
    .A2(_057_),
    .A3(_058_),
    .A4(_059_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _337_ (.A1(_055_),
    .A2(_060_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _338_ (.A1(\prescale_reg[17] ),
    .A2(\prescale_reg[18] ),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _339_ (.A1(_051_),
    .A2(_053_),
    .A3(_061_),
    .A4(_062_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input13 (.I(prescale[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _341_ (.I0(\data_reg[0] ),
    .I1(_049_),
    .S(_063_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _342_ (.A1(\data_reg[2] ),
    .A2(_047_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _343_ (.I0(\data_reg[1] ),
    .I1(_065_),
    .S(_063_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _344_ (.A1(\data_reg[3] ),
    .A2(_047_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _345_ (.I0(\data_reg[2] ),
    .I1(_066_),
    .S(_063_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _346_ (.A1(\data_reg[4] ),
    .A2(_047_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _347_ (.I0(\data_reg[3] ),
    .I1(_067_),
    .S(_063_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input12 (.I(prescale[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _349_ (.A1(\data_reg[5] ),
    .A2(_047_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _350_ (.I0(\data_reg[4] ),
    .I1(_069_),
    .S(_063_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _351_ (.A1(\data_reg[6] ),
    .A2(_047_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _352_ (.I0(\data_reg[5] ),
    .I1(_070_),
    .S(_063_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _353_ (.A1(\data_reg[7] ),
    .A2(_047_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _354_ (.I0(\data_reg[6] ),
    .I1(_071_),
    .S(_063_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _355_ (.A1(rxd_reg),
    .A2(_047_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _356_ (.I0(\data_reg[7] ),
    .I1(_072_),
    .S(_063_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _357_ (.I(net18),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input11 (.I(prescale[3]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input10 (.I(prescale[2]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _360_ (.A1(\bit_cnt[2] ),
    .A2(_052_),
    .B(rxd_reg),
    .C(\bit_cnt[3] ),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _361_ (.A1(_298_[0]),
    .A2(_047_),
    .A3(_076_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _362_ (.A1(_300_[0]),
    .A2(_045_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _363_ (.A1(\prescale_reg[3] ),
    .A2(\prescale_reg[2] ),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _364_ (.A1(\prescale_reg[17] ),
    .A2(\prescale_reg[16] ),
    .A3(\prescale_reg[18] ),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _365_ (.A1(_306_[0]),
    .A2(_079_),
    .A3(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _366_ (.A1(\prescale_reg[4] ),
    .A2(_058_),
    .A3(_059_),
    .A4(_054_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _367_ (.A1(rxd_reg),
    .A2(_078_),
    .B(_081_),
    .C(_082_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _368_ (.I0(\bit_cnt[0] ),
    .I1(_077_),
    .S(_083_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _369_ (.A1(_073_),
    .A2(_084_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _370_ (.I(\bit_cnt[2] ),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _371_ (.A1(_300_[0]),
    .A2(_302_[0]),
    .Z(_086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _372_ (.A1(rxd_reg),
    .A2(\bit_cnt[3] ),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _373_ (.A1(_085_),
    .A2(_086_),
    .B(_087_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input9 (.I(prescale[1]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _375_ (.A1(_301_[0]),
    .A2(_088_),
    .B(_047_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _376_ (.I0(\bit_cnt[1] ),
    .I1(_090_),
    .S(_083_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _377_ (.A1(_073_),
    .A2(_091_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _378_ (.A1(_306_[0]),
    .A2(_079_),
    .A3(_080_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _379_ (.A1(\prescale_reg[4] ),
    .A2(_058_),
    .A3(_059_),
    .A4(_054_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _380_ (.A1(_092_),
    .A2(_093_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input8 (.I(prescale[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _382_ (.I(_300_[0]),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _383_ (.A1(_096_),
    .A2(_087_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _384_ (.A1(_094_),
    .A2(_097_),
    .B(\bit_cnt[2] ),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _385_ (.A1(\bit_cnt[3] ),
    .A2(_085_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _386_ (.A1(_096_),
    .A2(_094_),
    .A3(_099_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input7 (.I(prescale[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input6 (.I(prescale[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _389_ (.A1(_098_),
    .A2(_100_),
    .B(net18),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input5 (.I(prescale[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _391_ (.A1(\bit_cnt[0] ),
    .A2(\bit_cnt[1] ),
    .A3(_099_),
    .B(_076_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _392_ (.A1(\bit_cnt[2] ),
    .A2(\bit_cnt[0] ),
    .A3(\bit_cnt[1] ),
    .B(_047_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _393_ (.A1(_083_),
    .A2(_105_),
    .B(\bit_cnt[3] ),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _394_ (.A1(_083_),
    .A2(_104_),
    .B(_106_),
    .C(net18),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _395_ (.I(rxd_reg),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _396_ (.A1(_078_),
    .A2(_092_),
    .A3(_093_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _397_ (.I0(net20),
    .I1(_107_),
    .S(_108_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _398_ (.A1(_073_),
    .A2(_109_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _399_ (.A1(_096_),
    .A2(_302_[0]),
    .A3(_045_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _400_ (.A1(rxd_reg),
    .A2(net18),
    .A3(_094_),
    .A4(_110_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _401_ (.A1(rxd_reg),
    .A2(_096_),
    .A3(_302_[0]),
    .A4(_045_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _402_ (.A1(\bit_cnt[0] ),
    .A2(_299_[0]),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _403_ (.A1(_092_),
    .A2(_093_),
    .A3(_111_),
    .A4(_112_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input4 (.I(prescale[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _405_ (.I0(net22),
    .I1(\data_reg[0] ),
    .S(_113_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _406_ (.A1(_073_),
    .A2(_115_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _407_ (.I0(net23),
    .I1(\data_reg[1] ),
    .S(_113_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _408_ (.A1(_073_),
    .A2(_116_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _409_ (.I0(net24),
    .I1(\data_reg[2] ),
    .S(_113_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _410_ (.A1(_073_),
    .A2(_117_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _411_ (.I0(net25),
    .I1(\data_reg[3] ),
    .S(_113_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _412_ (.A1(_073_),
    .A2(_118_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _413_ (.I0(net26),
    .I1(\data_reg[4] ),
    .S(_113_),
    .Z(_119_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _414_ (.A1(_073_),
    .A2(_119_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _415_ (.I0(net27),
    .I1(\data_reg[5] ),
    .S(_113_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _416_ (.A1(_073_),
    .A2(_120_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _417_ (.I0(net28),
    .I1(\data_reg[6] ),
    .S(_113_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _418_ (.A1(_073_),
    .A2(_121_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _419_ (.I0(net29),
    .I1(\data_reg[7] ),
    .S(_113_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _420_ (.A1(_073_),
    .A2(_122_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _421_ (.I(net1),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _422_ (.A1(_092_),
    .A2(_093_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input3 (.I(prescale[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _424_ (.A1(net30),
    .A2(_123_),
    .B1(_124_),
    .B2(_111_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _425_ (.A1(net18),
    .A2(_126_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _426_ (.A1(_073_),
    .A2(net30),
    .A3(_124_),
    .A4(_111_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _427_ (.A1(\prescale_reg[0] ),
    .A2(_094_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _428_ (.A1(_045_),
    .A2(_050_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _429_ (.A1(_047_),
    .A2(_076_),
    .A3(_110_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _430_ (.A1(_304_[0]),
    .A2(_128_),
    .B(_124_),
    .C(_129_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _431_ (.A1(_073_),
    .A2(_127_),
    .A3(_130_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input2 (.I(prescale[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _433_ (.I(_312_[0]),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _434_ (.A1(net10),
    .A2(net11),
    .Z(_133_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _435_ (.A1(net12),
    .A2(net13),
    .A3(net14),
    .Z(_134_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _436_ (.A1(net15),
    .A2(_132_),
    .A3(_133_),
    .A4(_134_),
    .Z(_135_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _437_ (.A1(net16),
    .A2(_135_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _438_ (.A1(net2),
    .A2(net10),
    .A3(net9),
    .A4(net11),
    .Z(_137_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(m_axis_tready),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _440_ (.A1(_137_),
    .A2(_134_),
    .B(net15),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _441_ (.A1(net15),
    .A2(_137_),
    .A3(_134_),
    .Z(_140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _442_ (.A1(_139_),
    .A2(_140_),
    .B(_078_),
    .C(_088_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _443_ (.A1(_078_),
    .A2(_136_),
    .B(_141_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _444_ (.A1(_128_),
    .A2(_092_),
    .A3(_093_),
    .Z(_143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _445_ (.A1(_073_),
    .A2(_143_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _446_ (.A1(\prescale_reg[10] ),
    .A2(_073_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _447_ (.A1(\prescale_reg[10] ),
    .A2(net18),
    .Z(_146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _448_ (.I(_308_[0]),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _449_ (.A1(\prescale_reg[9] ),
    .A2(_147_),
    .A3(_057_),
    .A4(_058_),
    .Z(_148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _450_ (.A1(_092_),
    .A2(_093_),
    .B(_148_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _451_ (.I0(_145_),
    .I1(_146_),
    .S(_149_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _452_ (.A1(_142_),
    .A2(_144_),
    .B(_150_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _453_ (.A1(_056_),
    .A2(_057_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _454_ (.A1(\prescale_reg[10] ),
    .A2(\prescale_reg[9] ),
    .Z(_152_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _455_ (.A1(_151_),
    .A2(_058_),
    .A3(_152_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _456_ (.A1(\prescale_reg[11] ),
    .A2(_153_),
    .Z(_154_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _457_ (.A1(_047_),
    .A2(_076_),
    .Z(_155_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _458_ (.A1(net15),
    .A2(net16),
    .A3(_137_),
    .A4(_134_),
    .Z(_156_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _459_ (.A1(net17),
    .A2(_156_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _460_ (.A1(_155_),
    .A2(_136_),
    .B1(_157_),
    .B2(_078_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _461_ (.A1(net18),
    .A2(_124_),
    .A3(_154_),
    .B1(_158_),
    .B2(_144_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _462_ (.A1(_147_),
    .A2(_057_),
    .Z(_159_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _463_ (.A1(\prescale_reg[11] ),
    .A2(_058_),
    .A3(_152_),
    .A4(_159_),
    .Z(_160_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _464_ (.A1(\prescale_reg[12] ),
    .A2(_160_),
    .Z(_161_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _465_ (.A1(net15),
    .A2(net16),
    .A3(net17),
    .Z(_162_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _466_ (.A1(_132_),
    .A2(_133_),
    .A3(_134_),
    .A4(_162_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _467_ (.A1(net3),
    .A2(_163_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _468_ (.A1(_155_),
    .A2(_157_),
    .B1(_164_),
    .B2(_078_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _469_ (.A1(net18),
    .A2(_124_),
    .A3(_161_),
    .B1(_165_),
    .B2(_144_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _470_ (.A1(_137_),
    .A2(_134_),
    .A3(_162_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _471_ (.A1(net4),
    .A2(_078_),
    .A3(_166_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _472_ (.A1(net3),
    .A2(net4),
    .Z(_168_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _473_ (.A1(_047_),
    .A2(_166_),
    .A3(_168_),
    .Z(_169_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _474_ (.A1(net3),
    .A2(_078_),
    .A3(_088_),
    .A4(_163_),
    .Z(_170_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _475_ (.A1(_167_),
    .A2(_169_),
    .A3(_170_),
    .Z(_171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _476_ (.A1(_051_),
    .A2(_124_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _477_ (.A1(\prescale_reg[13] ),
    .A2(_060_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _478_ (.A1(net18),
    .A2(_124_),
    .A3(_173_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _479_ (.A1(net3),
    .A2(_047_),
    .A3(_076_),
    .A4(_163_),
    .Z(_175_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _480_ (.A1(net3),
    .A2(net4),
    .A3(_078_),
    .Z(_176_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _481_ (.A1(_175_),
    .A2(_176_),
    .B(_051_),
    .C(_124_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _482_ (.A1(_171_),
    .A2(_172_),
    .B(_174_),
    .C(_177_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _483_ (.A1(_058_),
    .A2(_059_),
    .Z(_178_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _484_ (.A1(\prescale_reg[13] ),
    .A2(_178_),
    .A3(_159_),
    .Z(_179_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _485_ (.A1(\prescale_reg[14] ),
    .A2(_179_),
    .Z(_180_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _486_ (.A1(_107_),
    .A2(_300_[0]),
    .A3(_045_),
    .Z(_181_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _487_ (.A1(_163_),
    .A2(_168_),
    .B(_181_),
    .C(net5),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _488_ (.A1(\bit_cnt[3] ),
    .A2(\bit_cnt[2] ),
    .Z(_183_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _489_ (.A1(rxd_reg),
    .A2(_096_),
    .A3(_183_),
    .Z(_184_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _490_ (.A1(net5),
    .A2(_163_),
    .A3(_168_),
    .A4(_184_),
    .Z(_185_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _491_ (.A1(_124_),
    .A2(_182_),
    .A3(_185_),
    .Z(_186_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _492_ (.A1(net3),
    .A2(_137_),
    .A3(_134_),
    .A4(_162_),
    .Z(_187_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _493_ (.A1(net4),
    .A2(_187_),
    .Z(_188_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _494_ (.A1(_129_),
    .A2(_188_),
    .Z(_189_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _495_ (.A1(_094_),
    .A2(_180_),
    .B1(_186_),
    .B2(_189_),
    .C(net18),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _496_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .Z(_190_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _497_ (.A1(_137_),
    .A2(_134_),
    .A3(_162_),
    .A4(_190_),
    .Z(_191_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _498_ (.A1(net6),
    .A2(_191_),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _499_ (.A1(_132_),
    .A2(_133_),
    .A3(_134_),
    .A4(_162_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _500_ (.A1(net3),
    .A2(net4),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _501_ (.A1(_300_[0]),
    .A2(_045_),
    .B(net5),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _502_ (.A1(_076_),
    .A2(_193_),
    .A3(_194_),
    .A4(_195_),
    .Z(_196_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _503_ (.A1(_096_),
    .A2(_183_),
    .B(net5),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _504_ (.A1(_193_),
    .A2(_194_),
    .B(_197_),
    .C(_088_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _505_ (.A1(_078_),
    .A2(_192_),
    .B(_196_),
    .C(_198_),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _506_ (.A1(\prescale_reg[13] ),
    .A2(\prescale_reg[14] ),
    .A3(\prescale_reg[1] ),
    .A4(\prescale_reg[0] ),
    .Z(_200_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _507_ (.A1(_057_),
    .A2(_058_),
    .A3(_059_),
    .A4(_200_),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _508_ (.A1(\prescale_reg[15] ),
    .A2(_201_),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _509_ (.A1(_073_),
    .A2(_202_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _510_ (.A1(_045_),
    .A2(_050_),
    .Z(_204_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _511_ (.A1(\prescale_reg[15] ),
    .A2(_201_),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _512_ (.I0(_204_),
    .I1(_205_),
    .S(_094_),
    .Z(_206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _513_ (.A1(_143_),
    .A2(_199_),
    .B(_203_),
    .C(_206_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _514_ (.A1(_155_),
    .A2(_110_),
    .A3(_192_),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _515_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .A4(net6),
    .Z(_208_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _516_ (.A1(_163_),
    .A2(_208_),
    .B(_181_),
    .C(net7),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _517_ (.A1(net7),
    .A2(_163_),
    .A3(_184_),
    .A4(_208_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _518_ (.A1(_124_),
    .A2(_209_),
    .A3(_210_),
    .Z(_211_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _519_ (.A1(_308_[0]),
    .A2(_079_),
    .Z(_212_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _520_ (.A1(\prescale_reg[16] ),
    .A2(_093_),
    .A3(_212_),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _521_ (.A1(_073_),
    .A2(_213_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _522_ (.A1(_092_),
    .A2(_212_),
    .Z(_215_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _523_ (.A1(_093_),
    .A2(_215_),
    .B(\prescale_reg[16] ),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _524_ (.A1(_207_),
    .A2(_211_),
    .B(_214_),
    .C(_216_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _525_ (.A1(_055_),
    .A2(_060_),
    .B(\prescale_reg[17] ),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _526_ (.A1(\prescale_reg[17] ),
    .A2(_055_),
    .A3(_060_),
    .Z(_218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _527_ (.A1(_217_),
    .A2(_218_),
    .B(net18),
    .C(_124_),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _528_ (.A1(net7),
    .A2(_208_),
    .Z(_220_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _529_ (.A1(_166_),
    .A2(_220_),
    .B(net8),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _530_ (.A1(net8),
    .A2(_166_),
    .A3(_220_),
    .Z(_222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _531_ (.A1(_051_),
    .A2(_078_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _532_ (.A1(_221_),
    .A2(_222_),
    .B(_223_),
    .C(_094_),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _533_ (.A1(_163_),
    .A2(_208_),
    .B(net7),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _534_ (.A1(_163_),
    .A2(_220_),
    .Z(_226_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _535_ (.A1(_051_),
    .A2(_047_),
    .A3(_076_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _536_ (.A1(_225_),
    .A2(_226_),
    .B(_227_),
    .C(_094_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _537_ (.A1(_219_),
    .A2(_224_),
    .A3(_228_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _538_ (.A1(\prescale_reg[17] ),
    .A2(_178_),
    .A3(_055_),
    .A4(_159_),
    .Z(_229_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _539_ (.A1(\prescale_reg[18] ),
    .A2(_229_),
    .Z(_230_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _540_ (.I(net8),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _541_ (.A1(_300_[0]),
    .A2(_045_),
    .B(_231_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _542_ (.A1(_166_),
    .A2(_220_),
    .B(_232_),
    .C(_076_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _543_ (.A1(_096_),
    .A2(_183_),
    .B(_231_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _544_ (.A1(_088_),
    .A2(_166_),
    .A3(_220_),
    .A4(_234_),
    .Z(_235_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _545_ (.A1(net8),
    .A2(_047_),
    .A3(_163_),
    .A4(_220_),
    .Z(_236_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _546_ (.A1(_233_),
    .A2(_235_),
    .A3(_236_),
    .Z(_237_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _547_ (.A1(net18),
    .A2(_124_),
    .A3(_230_),
    .B1(_237_),
    .B2(_172_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _548_ (.A1(\prescale_reg[1] ),
    .A2(_128_),
    .B(_076_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _549_ (.I0(_307_[0]),
    .I1(_238_),
    .S(_124_),
    .Z(_239_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _550_ (.A1(net18),
    .A2(_239_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _551_ (.A1(net2),
    .A2(_078_),
    .B(_088_),
    .C(_204_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _552_ (.A1(\prescale_reg[2] ),
    .A2(_308_[0]),
    .Z(_241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _553_ (.I0(_240_),
    .I1(_241_),
    .S(_094_),
    .Z(_242_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _554_ (.A1(_073_),
    .A2(_242_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _555_ (.A1(\prescale_reg[2] ),
    .A2(_056_),
    .Z(_243_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _556_ (.A1(\prescale_reg[3] ),
    .A2(_243_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _557_ (.A1(_094_),
    .A2(_244_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _558_ (.A1(_313_[0]),
    .A2(_047_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _559_ (.A1(_310_[0]),
    .A2(_047_),
    .A3(_076_),
    .Z(_247_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _560_ (.A1(_246_),
    .A2(_247_),
    .B(_128_),
    .C(_124_),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _561_ (.A1(_245_),
    .A2(_248_),
    .B(net18),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _562_ (.A1(_313_[0]),
    .A2(_078_),
    .A3(_088_),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _563_ (.A1(net10),
    .A2(_312_[0]),
    .Z(_250_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _564_ (.A1(_078_),
    .A2(_250_),
    .Z(_251_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _565_ (.A1(_249_),
    .A2(_251_),
    .B(_128_),
    .C(_124_),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _566_ (.A1(_094_),
    .A2(_212_),
    .B(\prescale_reg[4] ),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _567_ (.A1(\prescale_reg[4] ),
    .A2(_212_),
    .B1(_252_),
    .B2(_253_),
    .C(net18),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _568_ (.A1(net2),
    .A2(net10),
    .A3(net9),
    .Z(_254_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _569_ (.A1(_300_[0]),
    .A2(net11),
    .A3(_045_),
    .A4(_254_),
    .ZN(_255_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _570_ (.A1(_047_),
    .A2(_137_),
    .B(_255_),
    .ZN(_256_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _571_ (.A1(_047_),
    .A2(_076_),
    .A3(_250_),
    .Z(_257_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _572_ (.A1(_256_),
    .A2(_257_),
    .B(_128_),
    .C(_124_),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _573_ (.A1(_092_),
    .A2(_093_),
    .B(_151_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _574_ (.A1(\prescale_reg[5] ),
    .A2(_259_),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _575_ (.A1(\prescale_reg[5] ),
    .A2(_259_),
    .Z(_261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _576_ (.A1(_258_),
    .A2(_260_),
    .B(_261_),
    .C(net18),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _577_ (.A1(\prescale_reg[5] ),
    .A2(_147_),
    .A3(_057_),
    .Z(_262_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _578_ (.A1(\prescale_reg[6] ),
    .A2(_262_),
    .ZN(_263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _579_ (.A1(_094_),
    .A2(_263_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _580_ (.A1(net11),
    .A2(_254_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _581_ (.A1(_137_),
    .A2(_265_),
    .B(_078_),
    .C(_088_),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _582_ (.A1(_132_),
    .A2(_133_),
    .B(net12),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _583_ (.A1(net12),
    .A2(_132_),
    .A3(_133_),
    .Z(_268_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _584_ (.A1(_267_),
    .A2(_268_),
    .B(_047_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _585_ (.A1(_266_),
    .A2(_269_),
    .B(_128_),
    .C(_124_),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _586_ (.A1(_264_),
    .A2(_270_),
    .B(net18),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _587_ (.I(net13),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _588_ (.A1(_096_),
    .A2(_183_),
    .B1(_133_),
    .B2(_132_),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _589_ (.A1(_271_),
    .A2(_047_),
    .B1(_088_),
    .B2(_272_),
    .ZN(_273_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _590_ (.A1(net12),
    .A2(net13),
    .Z(_274_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _591_ (.A1(_300_[0]),
    .A2(net13),
    .A3(_045_),
    .A4(_137_),
    .ZN(_275_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _592_ (.A1(_047_),
    .A2(_137_),
    .A3(_274_),
    .B(_275_),
    .ZN(_276_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _593_ (.A1(_078_),
    .A2(_088_),
    .A3(_268_),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _594_ (.A1(net12),
    .A2(_273_),
    .B(_276_),
    .C(_277_),
    .ZN(_278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _595_ (.A1(\prescale_reg[7] ),
    .A2(_073_),
    .ZN(_279_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _596_ (.A1(\prescale_reg[7] ),
    .A2(net18),
    .Z(_280_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _597_ (.A1(\prescale_reg[5] ),
    .A2(\prescale_reg[6] ),
    .A3(_056_),
    .A4(_057_),
    .Z(_281_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _598_ (.A1(_092_),
    .A2(_093_),
    .B(_281_),
    .ZN(_282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _599_ (.I0(_279_),
    .I1(_280_),
    .S(_282_),
    .Z(_283_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _600_ (.A1(_144_),
    .A2(_278_),
    .B(_283_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _601_ (.A1(\prescale_reg[5] ),
    .A2(\prescale_reg[7] ),
    .A3(\prescale_reg[6] ),
    .A4(_159_),
    .ZN(_284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _602_ (.A1(\prescale_reg[8] ),
    .A2(_284_),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _603_ (.A1(_132_),
    .A2(_133_),
    .A3(_134_),
    .Z(_286_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _604_ (.A1(_132_),
    .A2(_133_),
    .A3(_274_),
    .B(net14),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _605_ (.A1(_286_),
    .A2(_287_),
    .Z(_288_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _606_ (.A1(net12),
    .A2(_137_),
    .ZN(_289_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _607_ (.A1(net13),
    .A2(_289_),
    .ZN(_290_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _608_ (.A1(_184_),
    .A2(_288_),
    .B1(_290_),
    .B2(_129_),
    .C(_124_),
    .ZN(_291_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _609_ (.A1(\prescale_reg[8] ),
    .A2(_124_),
    .A3(_284_),
    .Z(_292_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _610_ (.A1(_073_),
    .A2(_285_),
    .A3(_291_),
    .A4(_292_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _611_ (.A1(_151_),
    .A2(_058_),
    .ZN(_293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _612_ (.A1(_286_),
    .A2(_287_),
    .B(_078_),
    .C(_088_),
    .ZN(_294_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _613_ (.A1(_139_),
    .A2(_140_),
    .B(_047_),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _614_ (.A1(_294_),
    .A2(_295_),
    .B(_143_),
    .ZN(_296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _615_ (.A1(_094_),
    .A2(_293_),
    .B(\prescale_reg[9] ),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _616_ (.A1(\prescale_reg[9] ),
    .A2(_293_),
    .B1(_296_),
    .B2(_297_),
    .C(net18),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _617_ (.A1(net18),
    .A2(net19),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _618_ (.A(_298_[0]),
    .B(_299_[0]),
    .CO(_300_[0]),
    .S(_301_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _619_ (.A(\bit_cnt[0] ),
    .B(_299_[0]),
    .CO(_302_[0]),
    .S(_303_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _620_ (.A(_304_[0]),
    .B(_305_[0]),
    .CO(_306_[0]),
    .S(_307_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _621_ (.A(_304_[0]),
    .B(_305_[0]),
    .CO(_308_[0]),
    .S(_309_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _622_ (.A(_310_[0]),
    .B(_311_[0]),
    .CO(_312_[0]),
    .S(_313_[0]));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bit_cnt[0]$_SDFFE_PP0P_  (.D(_000_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_cnt[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bit_cnt[1]$_SDFFE_PP0P_  (.D(_001_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_cnt[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bit_cnt[2]$_SDFFE_PP0P_  (.D(_002_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_cnt[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \bit_cnt[3]$_SDFFE_PP0P_  (.D(_003_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_cnt[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \busy_reg$_SDFFE_PP0P_  (.D(_004_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \data_reg[0]$_SDFFCE_PP0P_  (.D(_005_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\data_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \data_reg[1]$_SDFFCE_PP0P_  (.D(_006_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\data_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \data_reg[2]$_SDFFCE_PP0P_  (.D(_007_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\data_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \data_reg[3]$_SDFFCE_PP0P_  (.D(_008_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\data_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \data_reg[4]$_SDFFCE_PP0P_  (.D(_009_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\data_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \data_reg[5]$_SDFFCE_PP0P_  (.D(_010_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\data_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \data_reg[6]$_SDFFCE_PP0P_  (.D(_011_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\data_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \data_reg[7]$_SDFFCE_PP0P_  (.D(_012_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\data_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \frame_error_reg$_SDFF_PP0_  (.D(_013_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \m_axis_tdata_reg[0]$_SDFFE_PP0P_  (.D(_014_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \m_axis_tdata_reg[1]$_SDFFE_PP0P_  (.D(_015_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \m_axis_tdata_reg[2]$_SDFFE_PP0P_  (.D(_016_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \m_axis_tdata_reg[3]$_SDFFE_PP0P_  (.D(_017_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \m_axis_tdata_reg[4]$_SDFFE_PP0P_  (.D(_018_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \m_axis_tdata_reg[5]$_SDFFE_PP0P_  (.D(_019_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \m_axis_tdata_reg[6]$_SDFFE_PP0P_  (.D(_020_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \m_axis_tdata_reg[7]$_SDFFE_PP0P_  (.D(_021_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \m_axis_tvalid_reg$_SDFF_PP0_  (.D(_022_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \overrun_error_reg$_SDFF_PP0_  (.D(_023_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[0]$_SDFFE_PP0P_  (.D(_024_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\prescale_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[10]$_SDFFE_PP0P_  (.D(_025_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\prescale_reg[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[11]$_SDFFE_PP0P_  (.D(_026_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\prescale_reg[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[12]$_SDFFE_PP0P_  (.D(_027_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\prescale_reg[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[13]$_SDFFE_PP0P_  (.D(_028_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\prescale_reg[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[14]$_SDFFE_PP0P_  (.D(_029_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\prescale_reg[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[15]$_SDFFE_PP0P_  (.D(_030_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\prescale_reg[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[16]$_SDFFE_PP0P_  (.D(_031_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\prescale_reg[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[17]$_SDFFE_PP0P_  (.D(_032_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\prescale_reg[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[18]$_SDFFE_PP0P_  (.D(_033_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\prescale_reg[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[1]$_SDFFE_PP0P_  (.D(_034_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\prescale_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[2]$_SDFFE_PP0P_  (.D(_035_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\prescale_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[3]$_SDFFE_PP0P_  (.D(_036_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\prescale_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[4]$_SDFFE_PP0P_  (.D(_037_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\prescale_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[5]$_SDFFE_PP0P_  (.D(_038_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\prescale_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[6]$_SDFFE_PP0P_  (.D(_039_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\prescale_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[7]$_SDFFE_PP0P_  (.D(_040_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\prescale_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[8]$_SDFFE_PP0P_  (.D(_041_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\prescale_reg[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \prescale_reg[9]$_SDFFE_PP0P_  (.D(_042_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\prescale_reg[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \rxd_reg$_SDFF_PP1_  (.D(_043_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(rxd_reg));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_85 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_86 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_87 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_88 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_89 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_90 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_91 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_92 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_93 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_94 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_95 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_96 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_97 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_98 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_99 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input17 (.I(prescale[9]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 input18 (.I(rst),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input19 (.I(rxd),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output20 (.I(net20),
    .Z(busy));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output21 (.I(net21),
    .Z(frame_error));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output22 (.I(net22),
    .Z(m_axis_tdata[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output23 (.I(net23),
    .Z(m_axis_tdata[1]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output24 (.I(net24),
    .Z(m_axis_tdata[2]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output25 (.I(net25),
    .Z(m_axis_tdata[3]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output26 (.I(net26),
    .Z(m_axis_tdata[4]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output27 (.I(net27),
    .Z(m_axis_tdata[5]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output28 (.I(net28),
    .Z(m_axis_tdata[6]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output29 (.I(net29),
    .Z(m_axis_tdata[7]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output30 (.I(net30),
    .Z(m_axis_tvalid));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output31 (.I(net31),
    .Z(overrun_error));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload1 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload2 (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_11 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_396 ();
endmodule
