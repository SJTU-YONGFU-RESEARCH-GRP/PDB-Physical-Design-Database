module parameterized_spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire \bit_count[0] ;
 wire \bit_count[1] ;
 wire \bit_count[2] ;
 wire \bit_count[3] ;
 wire \clk_divider[0] ;
 wire \clk_divider[1] ;
 wire \clk_divider[2] ;
 wire \rx_shift[0] ;
 wire \rx_shift[1] ;
 wire \rx_shift[2] ;
 wire \rx_shift[3] ;
 wire \rx_shift[4] ;
 wire \rx_shift[5] ;
 wire \rx_shift[6] ;
 wire \rx_shift[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \tx_shift[0] ;
 wire \tx_shift[1] ;
 wire \tx_shift[2] ;
 wire \tx_shift[3] ;
 wire \tx_shift[4] ;
 wire \tx_shift[5] ;
 wire \tx_shift[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net26;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _139_ (.I(\bit_count[3] ),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _140_ (.A1(_122_),
    .A2(\bit_count[2] ),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _141_ (.A1(_120_),
    .A2(_037_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _142_ (.I(_126_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _143_ (.I(\state[0] ),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _144_ (.A1(\state[1] ),
    .A2(_038_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _145_ (.I(_039_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _146_ (.I(\bit_count[0] ),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _147_ (.I(\bit_count[1] ),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _148_ (.I(\bit_count[2] ),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _149_ (.A1(_040_),
    .A2(_116_),
    .A3(_117_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _150_ (.A1(\bit_count[3] ),
    .A2(_123_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _151_ (.I(\state[1] ),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _152_ (.I(_041_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _153_ (.A1(_042_),
    .A2(_116_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _154_ (.I(\clk_divider[2] ),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _155_ (.A1(_120_),
    .A2(net22),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _156_ (.A1(_129_),
    .A2(net22),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _157_ (.A1(\bit_count[3] ),
    .A2(_040_),
    .A3(_045_),
    .B(_046_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _158_ (.A1(_114_),
    .A2(_044_),
    .A3(_047_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _159_ (.I0(_116_),
    .I1(_043_),
    .S(_048_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _160_ (.A1(\state[0] ),
    .A2(net12),
    .B(_042_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _161_ (.A1(\bit_count[0] ),
    .A2(_050_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _162_ (.A1(_038_),
    .A2(_049_),
    .B(_051_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _163_ (.A1(\state[0] ),
    .A2(_114_),
    .A3(_044_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _164_ (.A1(_047_),
    .A2(_052_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _165_ (.A1(_042_),
    .A2(_119_),
    .A3(_053_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _166_ (.A1(_038_),
    .A2(net12),
    .B(_117_),
    .C(_053_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _167_ (.A1(\state[1] ),
    .A2(\bit_count[1] ),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _168_ (.A1(_054_),
    .A2(_055_),
    .A3(_056_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _169_ (.A1(_038_),
    .A2(net12),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _170_ (.A1(_129_),
    .A2(net22),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _171_ (.A1(_041_),
    .A2(\state[0] ),
    .A3(_114_),
    .A4(_044_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _172_ (.A1(_058_),
    .A2(_059_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _173_ (.A1(_053_),
    .A2(_057_),
    .B1(_060_),
    .B2(_120_),
    .C(_042_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _174_ (.A1(_120_),
    .A2(_058_),
    .A3(_059_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _175_ (.I0(_061_),
    .I1(_062_),
    .S(_040_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _176_ (.A1(_042_),
    .A2(_125_),
    .A3(_053_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _177_ (.A1(_038_),
    .A2(net12),
    .B(_053_),
    .C(_122_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _178_ (.A1(\state[1] ),
    .A2(\bit_count[3] ),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _179_ (.A1(_063_),
    .A2(_064_),
    .A3(_065_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _180_ (.A1(_114_),
    .A2(_044_),
    .B(\clk_divider[0] ),
    .C(_038_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _181_ (.I0(\clk_divider[0] ),
    .I1(_066_),
    .S(_042_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _182_ (.A1(_114_),
    .A2(_044_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _183_ (.A1(\state[0] ),
    .A2(_115_),
    .A3(_067_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _184_ (.I0(\clk_divider[1] ),
    .I1(_068_),
    .S(_042_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _185_ (.A1(_038_),
    .A2(_114_),
    .B(_042_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _186_ (.A1(\clk_divider[2] ),
    .A2(_069_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _187_ (.I0(\rx_shift[0] ),
    .I1(net13),
    .S(_039_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _188_ (.I0(\rx_shift[1] ),
    .I1(net14),
    .S(_039_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _189_ (.I0(\rx_shift[2] ),
    .I1(net15),
    .S(_039_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _190_ (.I0(\rx_shift[3] ),
    .I1(net16),
    .S(_039_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _191_ (.I0(\rx_shift[4] ),
    .I1(net17),
    .S(_039_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _192_ (.I0(\rx_shift[5] ),
    .I1(net18),
    .S(_039_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _193_ (.I0(\rx_shift[6] ),
    .I1(net19),
    .S(_039_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _194_ (.I0(\rx_shift[7] ),
    .I1(net20),
    .S(_039_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _195_ (.I(net22),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _196_ (.A1(_128_),
    .A2(_138_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _197_ (.A1(_128_),
    .A2(_138_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _198_ (.A1(_124_),
    .A2(_137_),
    .A3(_072_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _199_ (.A1(_124_),
    .A2(_137_),
    .A3(_071_),
    .B(_073_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _200_ (.I(_119_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _201_ (.A1(\bit_count[0] ),
    .A2(_075_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _202_ (.A1(\bit_count[2] ),
    .A2(_120_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _203_ (.A1(_134_),
    .A2(_131_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _204_ (.A1(_128_),
    .A2(_125_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _205_ (.A1(_076_),
    .A2(_077_),
    .A3(_078_),
    .A4(_079_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _206_ (.A1(_070_),
    .A2(_059_),
    .A3(_074_),
    .A4(_080_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _207_ (.I0(\rx_shift[0] ),
    .I1(net3),
    .S(_081_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _208_ (.I(_077_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _209_ (.A1(net22),
    .A2(_125_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _210_ (.A1(_059_),
    .A2(_082_),
    .A3(_083_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _211_ (.A1(_124_),
    .A2(_137_),
    .A3(_072_),
    .A4(_078_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _212_ (.A1(_116_),
    .A2(_119_),
    .A3(_085_),
    .Z(_086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _213_ (.A1(_084_),
    .A2(_086_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _214_ (.I0(net3),
    .I1(\rx_shift[1] ),
    .S(_087_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _215_ (.A1(\bit_count[0] ),
    .A2(_119_),
    .A3(_084_),
    .A4(_085_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _216_ (.I0(\rx_shift[2] ),
    .I1(net3),
    .S(_088_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _217_ (.A1(_116_),
    .A2(_075_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _218_ (.A1(_084_),
    .A2(_085_),
    .A3(_089_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _219_ (.I0(\rx_shift[3] ),
    .I1(net3),
    .S(_090_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _220_ (.A1(_076_),
    .A2(_084_),
    .A3(_085_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _221_ (.I0(\rx_shift[4] ),
    .I1(net3),
    .S(_091_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _222_ (.A1(_059_),
    .A2(_077_),
    .A3(_083_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _223_ (.A1(_086_),
    .A2(_092_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _224_ (.I0(net3),
    .I1(\rx_shift[5] ),
    .S(_093_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _225_ (.A1(\bit_count[0] ),
    .A2(_119_),
    .A3(_085_),
    .A4(_092_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _226_ (.I0(\rx_shift[6] ),
    .I1(net3),
    .S(_094_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _227_ (.A1(_085_),
    .A2(_089_),
    .A3(_092_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _228_ (.I0(\rx_shift[7] ),
    .I1(net3),
    .S(_095_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _229_ (.A1(\state[1] ),
    .A2(_067_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _230_ (.A1(net22),
    .A2(_096_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _231_ (.A1(\state[0] ),
    .A2(_097_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _232_ (.A1(_042_),
    .A2(net12),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _233_ (.I0(net23),
    .I1(_098_),
    .S(_038_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _234_ (.A1(_041_),
    .A2(\state[0] ),
    .Z(_099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _235_ (.I0(net11),
    .I1(\tx_shift[6] ),
    .S(_099_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _236_ (.A1(_058_),
    .A2(_052_),
    .B(_057_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _237_ (.A1(\state[1] ),
    .A2(_101_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _238_ (.I0(net24),
    .I1(_100_),
    .S(_102_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _239_ (.A1(\bit_count[3] ),
    .A2(_040_),
    .A3(_070_),
    .A4(_118_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _240_ (.A1(_052_),
    .A2(_103_),
    .B(_050_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _241_ (.A1(_059_),
    .A2(_103_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _242_ (.I(net12),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _243_ (.A1(_042_),
    .A2(_038_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _244_ (.I0(_104_),
    .I1(net25),
    .S(_105_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _245_ (.I(\tx_shift[0] ),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _246_ (.A1(_038_),
    .A2(net4),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _247_ (.A1(_106_),
    .A2(_102_),
    .B1(_107_),
    .B2(_098_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _248_ (.I0(net5),
    .I1(\tx_shift[0] ),
    .S(_099_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _249_ (.I0(\tx_shift[1] ),
    .I1(_108_),
    .S(_102_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _250_ (.I0(net6),
    .I1(\tx_shift[1] ),
    .S(_099_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _251_ (.I0(\tx_shift[2] ),
    .I1(_109_),
    .S(_102_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _252_ (.I0(net7),
    .I1(\tx_shift[2] ),
    .S(_099_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _253_ (.I0(\tx_shift[3] ),
    .I1(_110_),
    .S(_102_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _254_ (.I0(net8),
    .I1(\tx_shift[3] ),
    .S(_099_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _255_ (.I0(\tx_shift[4] ),
    .I1(_111_),
    .S(_102_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _256_ (.I0(net9),
    .I1(\tx_shift[4] ),
    .S(_099_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _257_ (.I0(\tx_shift[5] ),
    .I1(_112_),
    .S(_102_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _258_ (.I0(net10),
    .I1(\tx_shift[5] ),
    .S(_099_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _259_ (.I0(\tx_shift[6] ),
    .I1(_113_),
    .S(_102_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _260_ (.A(\clk_divider[0] ),
    .B(\clk_divider[1] ),
    .CO(_114_),
    .S(_115_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _261_ (.A(_116_),
    .B(_117_),
    .CO(_118_),
    .S(_119_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _262_ (.A(\bit_count[0] ),
    .B(\bit_count[1] ),
    .CO(_120_),
    .S(_121_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _263_ (.A(_122_),
    .B(_123_),
    .CO(_124_),
    .S(_125_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _264_ (.A(_122_),
    .B(_126_),
    .CO(_127_),
    .S(_128_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _265_ (.A(_122_),
    .B(_126_),
    .CO(_129_),
    .S(_130_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _266_ (.A(\bit_count[3] ),
    .B(_126_),
    .CO(_131_),
    .S(_132_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _267_ (.A(\bit_count[3] ),
    .B(_133_),
    .CO(_134_),
    .S(_135_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _268_ (.A(_122_),
    .B(_136_),
    .CO(_137_),
    .S(_138_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[0]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[1]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\bit_count[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[2]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[3]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_divider[0]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\clk_divider[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_divider[1]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\clk_divider[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_divider[2]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\clk_divider[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[0]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[1]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[2]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[3]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[4]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[5]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[6]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[7]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift[0]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rx_shift[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift[1]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\rx_shift[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift[2]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rx_shift[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift[3]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rx_shift[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift[4]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rx_shift[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift[5]$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift[6]$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift[7]$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rx_shift[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_valid$_DFF_PN0_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_clk$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \spi_cs_n$_DFFE_PN1P_  (.D(_025_),
    .SETN(net2),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_mosi$_DFFE_PN0P_  (.D(_026_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[0]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[1]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \tx_ready$_DFFE_PN1P_  (.D(_029_),
    .SETN(net2),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[0]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[1]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[2]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[3]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[4]$_DFFE_PN0P_  (.D(_034_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[5]$_DFFE_PN0P_  (.D(_035_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[6]$_DFFE_PN0P_  (.D(_036_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift[6] ));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 hold1 (.I(net2),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_67 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(net26),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input2 (.I(spi_miso),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(tx_data[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(tx_data[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(tx_data[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(tx_data[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(tx_data[4]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(tx_data[5]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(tx_data[6]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(tx_data[7]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input11 (.I(tx_valid),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(rx_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(rx_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(rx_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(rx_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(rx_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(rx_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(rx_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(rx_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(rx_valid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(spi_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(spi_cs_n));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(spi_mosi));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net25),
    .Z(tx_ready));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload1 (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload2 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_250 ();
endmodule
