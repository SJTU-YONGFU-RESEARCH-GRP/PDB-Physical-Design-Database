module gpio_controller (clk,
    int_out,
    rst_n,
    gpio_dir,
    gpio_in,
    gpio_out,
    gpio_pins,
    int_clear,
    int_enable,
    int_polarity,
    int_status,
    int_type);
 input clk;
 output int_out;
 input rst_n;
 input [31:0] gpio_dir;
 output [31:0] gpio_in;
 input [31:0] gpio_out;
 inout [31:0] gpio_pins;
 input [31:0] int_clear;
 input [31:0] int_enable;
 input [31:0] int_polarity;
 output [31:0] int_status;
 input [31:0] int_type;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire _486_;
 wire _487_;
 wire _488_;
 wire _489_;
 wire _490_;
 wire _491_;
 wire _492_;
 wire _493_;
 wire _494_;
 wire _495_;
 wire _496_;
 wire _497_;
 wire _498_;
 wire _499_;
 wire _500_;
 wire _501_;
 wire _502_;
 wire _503_;
 wire _504_;
 wire _505_;
 wire _506_;
 wire _507_;
 wire _508_;
 wire _509_;
 wire _510_;
 wire _511_;
 wire _512_;
 wire _513_;
 wire _514_;
 wire _515_;
 wire _516_;
 wire _517_;
 wire _518_;
 wire _519_;
 wire _520_;
 wire _521_;
 wire _522_;
 wire _523_;
 wire _524_;
 wire _525_;
 wire _526_;
 wire _527_;
 wire \gpio_in_prev[0] ;
 wire \gpio_in_prev[10] ;
 wire \gpio_in_prev[11] ;
 wire \gpio_in_prev[12] ;
 wire \gpio_in_prev[13] ;
 wire \gpio_in_prev[14] ;
 wire \gpio_in_prev[15] ;
 wire \gpio_in_prev[16] ;
 wire \gpio_in_prev[17] ;
 wire \gpio_in_prev[18] ;
 wire \gpio_in_prev[19] ;
 wire \gpio_in_prev[1] ;
 wire \gpio_in_prev[20] ;
 wire \gpio_in_prev[21] ;
 wire \gpio_in_prev[22] ;
 wire \gpio_in_prev[23] ;
 wire \gpio_in_prev[24] ;
 wire \gpio_in_prev[25] ;
 wire \gpio_in_prev[26] ;
 wire \gpio_in_prev[27] ;
 wire \gpio_in_prev[28] ;
 wire \gpio_in_prev[29] ;
 wire \gpio_in_prev[2] ;
 wire \gpio_in_prev[30] ;
 wire \gpio_in_prev[31] ;
 wire \gpio_in_prev[3] ;
 wire \gpio_in_prev[4] ;
 wire \gpio_in_prev[5] ;
 wire \gpio_in_prev[6] ;
 wire \gpio_in_prev[7] ;
 wire \gpio_in_prev[8] ;
 wire \gpio_in_prev[9] ;
 wire \gpio_in_sync1[0] ;
 wire \gpio_in_sync1[10] ;
 wire \gpio_in_sync1[11] ;
 wire \gpio_in_sync1[12] ;
 wire \gpio_in_sync1[13] ;
 wire \gpio_in_sync1[14] ;
 wire \gpio_in_sync1[15] ;
 wire \gpio_in_sync1[16] ;
 wire \gpio_in_sync1[17] ;
 wire \gpio_in_sync1[18] ;
 wire \gpio_in_sync1[19] ;
 wire \gpio_in_sync1[1] ;
 wire \gpio_in_sync1[20] ;
 wire \gpio_in_sync1[21] ;
 wire \gpio_in_sync1[22] ;
 wire \gpio_in_sync1[23] ;
 wire \gpio_in_sync1[24] ;
 wire \gpio_in_sync1[25] ;
 wire \gpio_in_sync1[26] ;
 wire \gpio_in_sync1[27] ;
 wire \gpio_in_sync1[28] ;
 wire \gpio_in_sync1[29] ;
 wire \gpio_in_sync1[2] ;
 wire \gpio_in_sync1[30] ;
 wire \gpio_in_sync1[31] ;
 wire \gpio_in_sync1[3] ;
 wire \gpio_in_sync1[4] ;
 wire \gpio_in_sync1[5] ;
 wire \gpio_in_sync1[6] ;
 wire \gpio_in_sync1[7] ;
 wire \gpio_in_sync1[8] ;
 wire \gpio_in_sync1[9] ;
 wire \gpio_in_sync2[0] ;
 wire \gpio_in_sync2[10] ;
 wire \gpio_in_sync2[11] ;
 wire \gpio_in_sync2[12] ;
 wire \gpio_in_sync2[13] ;
 wire \gpio_in_sync2[14] ;
 wire \gpio_in_sync2[15] ;
 wire \gpio_in_sync2[16] ;
 wire \gpio_in_sync2[17] ;
 wire \gpio_in_sync2[18] ;
 wire \gpio_in_sync2[19] ;
 wire \gpio_in_sync2[1] ;
 wire \gpio_in_sync2[20] ;
 wire \gpio_in_sync2[21] ;
 wire \gpio_in_sync2[22] ;
 wire \gpio_in_sync2[23] ;
 wire \gpio_in_sync2[24] ;
 wire \gpio_in_sync2[25] ;
 wire \gpio_in_sync2[26] ;
 wire \gpio_in_sync2[27] ;
 wire \gpio_in_sync2[28] ;
 wire \gpio_in_sync2[29] ;
 wire \gpio_in_sync2[2] ;
 wire \gpio_in_sync2[30] ;
 wire \gpio_in_sync2[31] ;
 wire \gpio_in_sync2[3] ;
 wire \gpio_in_sync2[4] ;
 wire \gpio_in_sync2[5] ;
 wire \gpio_in_sync2[6] ;
 wire \gpio_in_sync2[7] ;
 wire \gpio_in_sync2[8] ;
 wire \gpio_in_sync2[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 BUF_X4 _528_ (.A(rst_n),
    .Z(_128_));
 INV_X2 _529_ (.A(_128_),
    .ZN(_129_));
 BUF_X4 _530_ (.A(_129_),
    .Z(_130_));
 XNOR2_X1 _531_ (.A(\gpio_in_sync2[0] ),
    .B(\gpio_in_prev[0] ),
    .ZN(_131_));
 NAND2_X1 _532_ (.A1(net129),
    .A2(_131_),
    .ZN(_132_));
 XNOR2_X1 _533_ (.A(\gpio_in_sync2[0] ),
    .B(net97),
    .ZN(_133_));
 AND2_X1 _534_ (.A1(net65),
    .A2(_133_),
    .ZN(_134_));
 AOI21_X1 _535_ (.A(net194),
    .B1(_132_),
    .B2(_134_),
    .ZN(_135_));
 NOR3_X1 _536_ (.A1(net33),
    .A2(_130_),
    .A3(_135_),
    .ZN(_096_));
 OR2_X1 _537_ (.A1(_130_),
    .A2(net34),
    .ZN(_136_));
 NAND2_X1 _538_ (.A1(\gpio_in_sync2[10] ),
    .A2(net98),
    .ZN(_137_));
 AOI21_X1 _539_ (.A(_137_),
    .B1(\gpio_in_prev[10] ),
    .B2(net130),
    .ZN(_138_));
 OR2_X1 _540_ (.A1(\gpio_in_sync2[10] ),
    .A2(net98),
    .ZN(_139_));
 INV_X1 _541_ (.A(\gpio_in_prev[10] ),
    .ZN(_140_));
 AOI21_X1 _542_ (.A(_139_),
    .B1(_140_),
    .B2(net130),
    .ZN(_141_));
 OAI21_X1 _543_ (.A(net66),
    .B1(_138_),
    .B2(_141_),
    .ZN(_142_));
 INV_X1 _544_ (.A(net195),
    .ZN(_143_));
 AOI21_X1 _545_ (.A(_136_),
    .B1(_142_),
    .B2(_143_),
    .ZN(_097_));
 OR2_X1 _546_ (.A1(_130_),
    .A2(net35),
    .ZN(_144_));
 NAND2_X1 _547_ (.A1(\gpio_in_sync2[11] ),
    .A2(net99),
    .ZN(_145_));
 AOI21_X1 _548_ (.A(_145_),
    .B1(\gpio_in_prev[11] ),
    .B2(net131),
    .ZN(_146_));
 OR2_X1 _549_ (.A1(\gpio_in_sync2[11] ),
    .A2(net99),
    .ZN(_147_));
 INV_X1 _550_ (.A(\gpio_in_prev[11] ),
    .ZN(_148_));
 AOI21_X1 _551_ (.A(_147_),
    .B1(_148_),
    .B2(net131),
    .ZN(_149_));
 OAI21_X1 _552_ (.A(net67),
    .B1(_146_),
    .B2(_149_),
    .ZN(_150_));
 INV_X1 _553_ (.A(net196),
    .ZN(_151_));
 AOI21_X1 _554_ (.A(_144_),
    .B1(_150_),
    .B2(_151_),
    .ZN(_098_));
 OR2_X1 _555_ (.A1(_130_),
    .A2(net36),
    .ZN(_152_));
 NAND2_X1 _556_ (.A1(\gpio_in_sync2[12] ),
    .A2(net100),
    .ZN(_153_));
 AOI21_X1 _557_ (.A(_153_),
    .B1(\gpio_in_prev[12] ),
    .B2(net132),
    .ZN(_154_));
 OR2_X1 _558_ (.A1(\gpio_in_sync2[12] ),
    .A2(net100),
    .ZN(_155_));
 INV_X1 _559_ (.A(\gpio_in_prev[12] ),
    .ZN(_156_));
 AOI21_X1 _560_ (.A(_155_),
    .B1(_156_),
    .B2(net132),
    .ZN(_157_));
 OAI21_X1 _561_ (.A(net68),
    .B1(_154_),
    .B2(_157_),
    .ZN(_158_));
 INV_X1 _562_ (.A(net197),
    .ZN(_159_));
 AOI21_X1 _563_ (.A(_152_),
    .B1(_158_),
    .B2(_159_),
    .ZN(_099_));
 OR2_X1 _564_ (.A1(_130_),
    .A2(net37),
    .ZN(_160_));
 NAND2_X1 _565_ (.A1(\gpio_in_sync2[13] ),
    .A2(net101),
    .ZN(_161_));
 AOI21_X1 _566_ (.A(_161_),
    .B1(\gpio_in_prev[13] ),
    .B2(net133),
    .ZN(_162_));
 OR2_X1 _567_ (.A1(\gpio_in_sync2[13] ),
    .A2(net101),
    .ZN(_163_));
 INV_X1 _568_ (.A(\gpio_in_prev[13] ),
    .ZN(_164_));
 AOI21_X1 _569_ (.A(_163_),
    .B1(_164_),
    .B2(net133),
    .ZN(_165_));
 OAI21_X1 _570_ (.A(net69),
    .B1(_162_),
    .B2(_165_),
    .ZN(_166_));
 INV_X1 _571_ (.A(net198),
    .ZN(_167_));
 AOI21_X1 _572_ (.A(_160_),
    .B1(_166_),
    .B2(_167_),
    .ZN(_100_));
 OR2_X1 _573_ (.A1(_130_),
    .A2(net38),
    .ZN(_168_));
 NAND2_X1 _574_ (.A1(\gpio_in_sync2[14] ),
    .A2(net102),
    .ZN(_169_));
 AOI21_X1 _575_ (.A(_169_),
    .B1(\gpio_in_prev[14] ),
    .B2(net134),
    .ZN(_170_));
 OR2_X1 _576_ (.A1(\gpio_in_sync2[14] ),
    .A2(net102),
    .ZN(_171_));
 INV_X1 _577_ (.A(\gpio_in_prev[14] ),
    .ZN(_172_));
 AOI21_X1 _578_ (.A(_171_),
    .B1(_172_),
    .B2(net134),
    .ZN(_173_));
 OAI21_X1 _579_ (.A(net70),
    .B1(_170_),
    .B2(_173_),
    .ZN(_174_));
 INV_X1 _580_ (.A(net199),
    .ZN(_175_));
 AOI21_X1 _581_ (.A(_168_),
    .B1(_174_),
    .B2(_175_),
    .ZN(_101_));
 OR2_X1 _582_ (.A1(_130_),
    .A2(net39),
    .ZN(_176_));
 NAND2_X1 _583_ (.A1(\gpio_in_sync2[15] ),
    .A2(net103),
    .ZN(_177_));
 AOI21_X1 _584_ (.A(_177_),
    .B1(\gpio_in_prev[15] ),
    .B2(net135),
    .ZN(_178_));
 OR2_X1 _585_ (.A1(\gpio_in_sync2[15] ),
    .A2(net103),
    .ZN(_179_));
 INV_X1 _586_ (.A(\gpio_in_prev[15] ),
    .ZN(_180_));
 AOI21_X1 _587_ (.A(_179_),
    .B1(_180_),
    .B2(net135),
    .ZN(_181_));
 OAI21_X1 _588_ (.A(net71),
    .B1(_178_),
    .B2(_181_),
    .ZN(_182_));
 INV_X1 _589_ (.A(net200),
    .ZN(_183_));
 AOI21_X1 _590_ (.A(_176_),
    .B1(_182_),
    .B2(_183_),
    .ZN(_102_));
 OR2_X1 _591_ (.A1(_130_),
    .A2(net40),
    .ZN(_184_));
 NAND2_X1 _592_ (.A1(\gpio_in_sync2[16] ),
    .A2(net104),
    .ZN(_185_));
 AOI21_X1 _593_ (.A(_185_),
    .B1(\gpio_in_prev[16] ),
    .B2(net136),
    .ZN(_186_));
 OR2_X1 _594_ (.A1(\gpio_in_sync2[16] ),
    .A2(net104),
    .ZN(_187_));
 INV_X1 _595_ (.A(\gpio_in_prev[16] ),
    .ZN(_188_));
 AOI21_X1 _596_ (.A(_187_),
    .B1(_188_),
    .B2(net136),
    .ZN(_189_));
 OAI21_X1 _597_ (.A(net72),
    .B1(_186_),
    .B2(_189_),
    .ZN(_190_));
 INV_X1 _598_ (.A(net201),
    .ZN(_191_));
 AOI21_X1 _599_ (.A(_184_),
    .B1(_190_),
    .B2(_191_),
    .ZN(_103_));
 BUF_X2 _600_ (.A(_129_),
    .Z(_192_));
 OR2_X1 _601_ (.A1(_192_),
    .A2(net41),
    .ZN(_193_));
 NAND2_X1 _602_ (.A1(\gpio_in_sync2[17] ),
    .A2(net105),
    .ZN(_194_));
 AOI21_X1 _603_ (.A(_194_),
    .B1(\gpio_in_prev[17] ),
    .B2(net137),
    .ZN(_195_));
 OR2_X1 _604_ (.A1(\gpio_in_sync2[17] ),
    .A2(net105),
    .ZN(_196_));
 INV_X1 _605_ (.A(\gpio_in_prev[17] ),
    .ZN(_197_));
 AOI21_X1 _606_ (.A(_196_),
    .B1(_197_),
    .B2(net137),
    .ZN(_198_));
 OAI21_X1 _607_ (.A(net73),
    .B1(_195_),
    .B2(_198_),
    .ZN(_199_));
 INV_X1 _608_ (.A(net202),
    .ZN(_200_));
 AOI21_X1 _609_ (.A(_193_),
    .B1(_199_),
    .B2(_200_),
    .ZN(_104_));
 OR2_X1 _610_ (.A1(_192_),
    .A2(net42),
    .ZN(_201_));
 NAND2_X1 _611_ (.A1(\gpio_in_sync2[18] ),
    .A2(net106),
    .ZN(_202_));
 AOI21_X1 _612_ (.A(_202_),
    .B1(\gpio_in_prev[18] ),
    .B2(net138),
    .ZN(_203_));
 OR2_X1 _613_ (.A1(\gpio_in_sync2[18] ),
    .A2(net106),
    .ZN(_204_));
 INV_X1 _614_ (.A(\gpio_in_prev[18] ),
    .ZN(_205_));
 AOI21_X1 _615_ (.A(_204_),
    .B1(_205_),
    .B2(net138),
    .ZN(_206_));
 OAI21_X1 _616_ (.A(net74),
    .B1(_203_),
    .B2(_206_),
    .ZN(_207_));
 INV_X1 _617_ (.A(net203),
    .ZN(_208_));
 AOI21_X1 _618_ (.A(_201_),
    .B1(_207_),
    .B2(_208_),
    .ZN(_105_));
 OR2_X1 _619_ (.A1(_192_),
    .A2(net43),
    .ZN(_209_));
 NAND2_X1 _620_ (.A1(\gpio_in_sync2[19] ),
    .A2(net107),
    .ZN(_210_));
 AOI21_X1 _621_ (.A(_210_),
    .B1(\gpio_in_prev[19] ),
    .B2(net139),
    .ZN(_211_));
 OR2_X1 _622_ (.A1(\gpio_in_sync2[19] ),
    .A2(net107),
    .ZN(_212_));
 INV_X1 _623_ (.A(\gpio_in_prev[19] ),
    .ZN(_213_));
 AOI21_X1 _624_ (.A(_212_),
    .B1(_213_),
    .B2(net139),
    .ZN(_214_));
 OAI21_X1 _625_ (.A(net75),
    .B1(_211_),
    .B2(_214_),
    .ZN(_215_));
 INV_X1 _626_ (.A(net204),
    .ZN(_216_));
 AOI21_X1 _627_ (.A(_209_),
    .B1(_215_),
    .B2(_216_),
    .ZN(_106_));
 XNOR2_X1 _628_ (.A(\gpio_in_sync2[1] ),
    .B(\gpio_in_prev[1] ),
    .ZN(_217_));
 NAND2_X1 _629_ (.A1(net140),
    .A2(_217_),
    .ZN(_218_));
 XNOR2_X1 _630_ (.A(\gpio_in_sync2[1] ),
    .B(net108),
    .ZN(_219_));
 AND2_X1 _631_ (.A1(net76),
    .A2(_219_),
    .ZN(_220_));
 AOI21_X1 _632_ (.A(net205),
    .B1(_218_),
    .B2(_220_),
    .ZN(_221_));
 NOR3_X1 _633_ (.A1(_130_),
    .A2(net44),
    .A3(_221_),
    .ZN(_107_));
 OR2_X1 _634_ (.A1(_192_),
    .A2(net45),
    .ZN(_222_));
 NAND2_X1 _635_ (.A1(\gpio_in_sync2[20] ),
    .A2(net109),
    .ZN(_223_));
 AOI21_X1 _636_ (.A(_223_),
    .B1(\gpio_in_prev[20] ),
    .B2(net141),
    .ZN(_224_));
 OR2_X1 _637_ (.A1(\gpio_in_sync2[20] ),
    .A2(net109),
    .ZN(_225_));
 INV_X1 _638_ (.A(\gpio_in_prev[20] ),
    .ZN(_226_));
 AOI21_X1 _639_ (.A(_225_),
    .B1(_226_),
    .B2(net141),
    .ZN(_227_));
 OAI21_X1 _640_ (.A(net77),
    .B1(_224_),
    .B2(_227_),
    .ZN(_228_));
 INV_X1 _641_ (.A(net206),
    .ZN(_229_));
 AOI21_X1 _642_ (.A(_222_),
    .B1(_228_),
    .B2(_229_),
    .ZN(_108_));
 OR2_X1 _643_ (.A1(_192_),
    .A2(net46),
    .ZN(_230_));
 NAND2_X1 _644_ (.A1(\gpio_in_sync2[21] ),
    .A2(net110),
    .ZN(_231_));
 AOI21_X1 _645_ (.A(_231_),
    .B1(\gpio_in_prev[21] ),
    .B2(net142),
    .ZN(_232_));
 OR2_X1 _646_ (.A1(\gpio_in_sync2[21] ),
    .A2(net110),
    .ZN(_233_));
 INV_X1 _647_ (.A(\gpio_in_prev[21] ),
    .ZN(_234_));
 AOI21_X1 _648_ (.A(_233_),
    .B1(_234_),
    .B2(net142),
    .ZN(_235_));
 OAI21_X1 _649_ (.A(net78),
    .B1(_232_),
    .B2(_235_),
    .ZN(_236_));
 INV_X1 _650_ (.A(net207),
    .ZN(_237_));
 AOI21_X1 _651_ (.A(_230_),
    .B1(_236_),
    .B2(_237_),
    .ZN(_109_));
 OR2_X1 _652_ (.A1(_192_),
    .A2(net47),
    .ZN(_238_));
 NAND2_X1 _653_ (.A1(\gpio_in_sync2[22] ),
    .A2(net111),
    .ZN(_239_));
 AOI21_X1 _654_ (.A(_239_),
    .B1(\gpio_in_prev[22] ),
    .B2(net143),
    .ZN(_240_));
 OR2_X1 _655_ (.A1(\gpio_in_sync2[22] ),
    .A2(net111),
    .ZN(_241_));
 INV_X1 _656_ (.A(\gpio_in_prev[22] ),
    .ZN(_242_));
 AOI21_X1 _657_ (.A(_241_),
    .B1(_242_),
    .B2(net143),
    .ZN(_243_));
 OAI21_X1 _658_ (.A(net79),
    .B1(_240_),
    .B2(_243_),
    .ZN(_244_));
 INV_X1 _659_ (.A(net208),
    .ZN(_245_));
 AOI21_X1 _660_ (.A(_238_),
    .B1(_244_),
    .B2(_245_),
    .ZN(_110_));
 OR2_X1 _661_ (.A1(_192_),
    .A2(net48),
    .ZN(_246_));
 NAND2_X1 _662_ (.A1(\gpio_in_sync2[23] ),
    .A2(net112),
    .ZN(_247_));
 AOI21_X1 _663_ (.A(_247_),
    .B1(\gpio_in_prev[23] ),
    .B2(net144),
    .ZN(_248_));
 OR2_X1 _664_ (.A1(\gpio_in_sync2[23] ),
    .A2(net112),
    .ZN(_249_));
 INV_X1 _665_ (.A(\gpio_in_prev[23] ),
    .ZN(_250_));
 AOI21_X1 _666_ (.A(_249_),
    .B1(_250_),
    .B2(net144),
    .ZN(_251_));
 OAI21_X1 _667_ (.A(net80),
    .B1(_248_),
    .B2(_251_),
    .ZN(_252_));
 INV_X1 _668_ (.A(net209),
    .ZN(_253_));
 AOI21_X1 _669_ (.A(_246_),
    .B1(_252_),
    .B2(_253_),
    .ZN(_111_));
 OR2_X1 _670_ (.A1(_192_),
    .A2(net49),
    .ZN(_254_));
 NAND2_X1 _671_ (.A1(\gpio_in_sync2[24] ),
    .A2(net113),
    .ZN(_255_));
 AOI21_X1 _672_ (.A(_255_),
    .B1(\gpio_in_prev[24] ),
    .B2(net145),
    .ZN(_256_));
 OR2_X1 _673_ (.A1(\gpio_in_sync2[24] ),
    .A2(net113),
    .ZN(_257_));
 INV_X1 _674_ (.A(\gpio_in_prev[24] ),
    .ZN(_258_));
 AOI21_X1 _675_ (.A(_257_),
    .B1(_258_),
    .B2(net145),
    .ZN(_259_));
 OAI21_X1 _676_ (.A(net81),
    .B1(_256_),
    .B2(_259_),
    .ZN(_260_));
 INV_X1 _677_ (.A(net210),
    .ZN(_261_));
 AOI21_X1 _678_ (.A(_254_),
    .B1(_260_),
    .B2(_261_),
    .ZN(_112_));
 OR2_X1 _679_ (.A1(_192_),
    .A2(net50),
    .ZN(_262_));
 NAND2_X1 _680_ (.A1(\gpio_in_sync2[25] ),
    .A2(net114),
    .ZN(_263_));
 AOI21_X1 _681_ (.A(_263_),
    .B1(\gpio_in_prev[25] ),
    .B2(net146),
    .ZN(_264_));
 OR2_X1 _682_ (.A1(\gpio_in_sync2[25] ),
    .A2(net114),
    .ZN(_265_));
 INV_X1 _683_ (.A(\gpio_in_prev[25] ),
    .ZN(_266_));
 AOI21_X1 _684_ (.A(_265_),
    .B1(_266_),
    .B2(net146),
    .ZN(_267_));
 OAI21_X1 _685_ (.A(net82),
    .B1(_264_),
    .B2(_267_),
    .ZN(_268_));
 INV_X1 _686_ (.A(net211),
    .ZN(_269_));
 AOI21_X1 _687_ (.A(_262_),
    .B1(_268_),
    .B2(_269_),
    .ZN(_113_));
 OR2_X1 _688_ (.A1(_192_),
    .A2(net51),
    .ZN(_270_));
 NAND2_X1 _689_ (.A1(\gpio_in_sync2[26] ),
    .A2(net115),
    .ZN(_271_));
 AOI21_X1 _690_ (.A(_271_),
    .B1(\gpio_in_prev[26] ),
    .B2(net147),
    .ZN(_272_));
 OR2_X1 _691_ (.A1(\gpio_in_sync2[26] ),
    .A2(net115),
    .ZN(_273_));
 INV_X1 _692_ (.A(\gpio_in_prev[26] ),
    .ZN(_274_));
 AOI21_X1 _693_ (.A(_273_),
    .B1(_274_),
    .B2(net147),
    .ZN(_275_));
 OAI21_X1 _694_ (.A(net83),
    .B1(_272_),
    .B2(_275_),
    .ZN(_276_));
 INV_X1 _695_ (.A(net212),
    .ZN(_277_));
 AOI21_X1 _696_ (.A(_270_),
    .B1(_276_),
    .B2(_277_),
    .ZN(_114_));
 BUF_X2 _697_ (.A(_129_),
    .Z(_278_));
 OR2_X1 _698_ (.A1(_278_),
    .A2(net52),
    .ZN(_279_));
 NAND2_X1 _699_ (.A1(\gpio_in_sync2[27] ),
    .A2(net116),
    .ZN(_280_));
 AOI21_X1 _700_ (.A(_280_),
    .B1(\gpio_in_prev[27] ),
    .B2(net148),
    .ZN(_281_));
 OR2_X1 _701_ (.A1(\gpio_in_sync2[27] ),
    .A2(net116),
    .ZN(_282_));
 INV_X1 _702_ (.A(\gpio_in_prev[27] ),
    .ZN(_283_));
 AOI21_X1 _703_ (.A(_282_),
    .B1(_283_),
    .B2(net148),
    .ZN(_284_));
 OAI21_X1 _704_ (.A(net84),
    .B1(_281_),
    .B2(_284_),
    .ZN(_285_));
 INV_X1 _705_ (.A(net213),
    .ZN(_286_));
 AOI21_X1 _706_ (.A(_279_),
    .B1(_285_),
    .B2(_286_),
    .ZN(_115_));
 OR2_X1 _707_ (.A1(_278_),
    .A2(net53),
    .ZN(_287_));
 NAND2_X1 _708_ (.A1(\gpio_in_sync2[28] ),
    .A2(net117),
    .ZN(_288_));
 AOI21_X1 _709_ (.A(_288_),
    .B1(\gpio_in_prev[28] ),
    .B2(net149),
    .ZN(_289_));
 OR2_X1 _710_ (.A1(\gpio_in_sync2[28] ),
    .A2(net117),
    .ZN(_290_));
 INV_X1 _711_ (.A(\gpio_in_prev[28] ),
    .ZN(_291_));
 AOI21_X1 _712_ (.A(_290_),
    .B1(_291_),
    .B2(net149),
    .ZN(_292_));
 OAI21_X1 _713_ (.A(net85),
    .B1(_289_),
    .B2(_292_),
    .ZN(_293_));
 INV_X1 _714_ (.A(net214),
    .ZN(_294_));
 AOI21_X1 _715_ (.A(_287_),
    .B1(_293_),
    .B2(_294_),
    .ZN(_116_));
 OR2_X1 _716_ (.A1(_278_),
    .A2(net54),
    .ZN(_295_));
 NAND2_X1 _717_ (.A1(\gpio_in_sync2[29] ),
    .A2(net118),
    .ZN(_296_));
 AOI21_X1 _718_ (.A(_296_),
    .B1(\gpio_in_prev[29] ),
    .B2(net150),
    .ZN(_297_));
 OR2_X1 _719_ (.A1(\gpio_in_sync2[29] ),
    .A2(net118),
    .ZN(_298_));
 INV_X1 _720_ (.A(\gpio_in_prev[29] ),
    .ZN(_299_));
 AOI21_X1 _721_ (.A(_298_),
    .B1(_299_),
    .B2(net150),
    .ZN(_300_));
 OAI21_X1 _722_ (.A(net86),
    .B1(_297_),
    .B2(_300_),
    .ZN(_301_));
 INV_X1 _723_ (.A(net215),
    .ZN(_302_));
 AOI21_X1 _724_ (.A(_295_),
    .B1(_301_),
    .B2(_302_),
    .ZN(_117_));
 XNOR2_X1 _725_ (.A(\gpio_in_sync2[2] ),
    .B(\gpio_in_prev[2] ),
    .ZN(_303_));
 NAND2_X1 _726_ (.A1(net151),
    .A2(_303_),
    .ZN(_304_));
 XNOR2_X1 _727_ (.A(\gpio_in_sync2[2] ),
    .B(net119),
    .ZN(_305_));
 AND2_X1 _728_ (.A1(net87),
    .A2(_305_),
    .ZN(_306_));
 AOI21_X1 _729_ (.A(net216),
    .B1(_304_),
    .B2(_306_),
    .ZN(_307_));
 NOR3_X1 _730_ (.A1(_130_),
    .A2(net55),
    .A3(_307_),
    .ZN(_118_));
 OR2_X1 _731_ (.A1(_278_),
    .A2(net56),
    .ZN(_308_));
 NAND2_X1 _732_ (.A1(\gpio_in_sync2[30] ),
    .A2(net120),
    .ZN(_309_));
 AOI21_X1 _733_ (.A(_309_),
    .B1(\gpio_in_prev[30] ),
    .B2(net152),
    .ZN(_310_));
 OR2_X1 _734_ (.A1(\gpio_in_sync2[30] ),
    .A2(net120),
    .ZN(_311_));
 INV_X1 _735_ (.A(\gpio_in_prev[30] ),
    .ZN(_312_));
 AOI21_X1 _736_ (.A(_311_),
    .B1(_312_),
    .B2(net152),
    .ZN(_313_));
 OAI21_X1 _737_ (.A(net88),
    .B1(_310_),
    .B2(_313_),
    .ZN(_314_));
 INV_X1 _738_ (.A(net217),
    .ZN(_315_));
 AOI21_X1 _739_ (.A(_308_),
    .B1(_314_),
    .B2(_315_),
    .ZN(_119_));
 OR2_X1 _740_ (.A1(_278_),
    .A2(net57),
    .ZN(_316_));
 NAND2_X1 _741_ (.A1(\gpio_in_sync2[31] ),
    .A2(net121),
    .ZN(_317_));
 AOI21_X1 _742_ (.A(_317_),
    .B1(\gpio_in_prev[31] ),
    .B2(net153),
    .ZN(_318_));
 OR2_X1 _743_ (.A1(\gpio_in_sync2[31] ),
    .A2(net121),
    .ZN(_319_));
 INV_X1 _744_ (.A(\gpio_in_prev[31] ),
    .ZN(_320_));
 AOI21_X1 _745_ (.A(_319_),
    .B1(_320_),
    .B2(net153),
    .ZN(_321_));
 OAI21_X1 _746_ (.A(net89),
    .B1(_318_),
    .B2(_321_),
    .ZN(_322_));
 INV_X1 _747_ (.A(net218),
    .ZN(_323_));
 AOI21_X1 _748_ (.A(_316_),
    .B1(_322_),
    .B2(_323_),
    .ZN(_120_));
 OR2_X1 _749_ (.A1(_278_),
    .A2(net58),
    .ZN(_324_));
 NAND2_X1 _750_ (.A1(\gpio_in_sync2[3] ),
    .A2(net122),
    .ZN(_325_));
 AOI21_X1 _751_ (.A(_325_),
    .B1(net154),
    .B2(\gpio_in_prev[3] ),
    .ZN(_326_));
 OR2_X1 _752_ (.A1(\gpio_in_sync2[3] ),
    .A2(net122),
    .ZN(_327_));
 INV_X1 _753_ (.A(\gpio_in_prev[3] ),
    .ZN(_328_));
 AOI21_X1 _754_ (.A(_327_),
    .B1(net154),
    .B2(_328_),
    .ZN(_329_));
 OAI21_X1 _755_ (.A(net90),
    .B1(_326_),
    .B2(_329_),
    .ZN(_330_));
 INV_X1 _756_ (.A(net219),
    .ZN(_331_));
 AOI21_X1 _757_ (.A(_324_),
    .B1(_330_),
    .B2(_331_),
    .ZN(_121_));
 OR2_X1 _758_ (.A1(_278_),
    .A2(net59),
    .ZN(_332_));
 NAND2_X1 _759_ (.A1(\gpio_in_sync2[4] ),
    .A2(net123),
    .ZN(_333_));
 AOI21_X1 _760_ (.A(_333_),
    .B1(net155),
    .B2(\gpio_in_prev[4] ),
    .ZN(_334_));
 OR2_X1 _761_ (.A1(\gpio_in_sync2[4] ),
    .A2(net123),
    .ZN(_335_));
 INV_X1 _762_ (.A(\gpio_in_prev[4] ),
    .ZN(_336_));
 AOI21_X1 _763_ (.A(_335_),
    .B1(net155),
    .B2(_336_),
    .ZN(_337_));
 OAI21_X1 _764_ (.A(net91),
    .B1(_334_),
    .B2(_337_),
    .ZN(_338_));
 INV_X1 _765_ (.A(net220),
    .ZN(_339_));
 AOI21_X1 _766_ (.A(_332_),
    .B1(_338_),
    .B2(_339_),
    .ZN(_122_));
 OR2_X1 _767_ (.A1(_278_),
    .A2(net60),
    .ZN(_340_));
 NAND2_X1 _768_ (.A1(\gpio_in_sync2[5] ),
    .A2(net124),
    .ZN(_341_));
 AOI21_X1 _769_ (.A(_341_),
    .B1(net156),
    .B2(\gpio_in_prev[5] ),
    .ZN(_342_));
 OR2_X1 _770_ (.A1(\gpio_in_sync2[5] ),
    .A2(net124),
    .ZN(_343_));
 INV_X1 _771_ (.A(\gpio_in_prev[5] ),
    .ZN(_344_));
 AOI21_X1 _772_ (.A(_343_),
    .B1(net156),
    .B2(_344_),
    .ZN(_345_));
 OAI21_X1 _773_ (.A(net92),
    .B1(_342_),
    .B2(_345_),
    .ZN(_346_));
 INV_X1 _774_ (.A(net221),
    .ZN(_347_));
 AOI21_X1 _775_ (.A(_340_),
    .B1(_346_),
    .B2(_347_),
    .ZN(_123_));
 OR2_X1 _776_ (.A1(_278_),
    .A2(net61),
    .ZN(_348_));
 NAND2_X1 _777_ (.A1(\gpio_in_sync2[6] ),
    .A2(net125),
    .ZN(_349_));
 AOI21_X1 _778_ (.A(_349_),
    .B1(net157),
    .B2(\gpio_in_prev[6] ),
    .ZN(_350_));
 OR2_X1 _779_ (.A1(\gpio_in_sync2[6] ),
    .A2(net125),
    .ZN(_351_));
 INV_X1 _780_ (.A(\gpio_in_prev[6] ),
    .ZN(_352_));
 AOI21_X1 _781_ (.A(_351_),
    .B1(net157),
    .B2(_352_),
    .ZN(_353_));
 OAI21_X1 _782_ (.A(net93),
    .B1(_350_),
    .B2(_353_),
    .ZN(_354_));
 INV_X1 _783_ (.A(net222),
    .ZN(_355_));
 AOI21_X1 _784_ (.A(_348_),
    .B1(_354_),
    .B2(_355_),
    .ZN(_124_));
 OR2_X1 _785_ (.A1(_278_),
    .A2(net62),
    .ZN(_356_));
 NAND2_X1 _786_ (.A1(\gpio_in_sync2[7] ),
    .A2(net126),
    .ZN(_357_));
 AOI21_X1 _787_ (.A(_357_),
    .B1(net158),
    .B2(\gpio_in_prev[7] ),
    .ZN(_358_));
 OR2_X1 _788_ (.A1(\gpio_in_sync2[7] ),
    .A2(net126),
    .ZN(_359_));
 INV_X1 _789_ (.A(\gpio_in_prev[7] ),
    .ZN(_360_));
 AOI21_X1 _790_ (.A(_359_),
    .B1(net158),
    .B2(_360_),
    .ZN(_361_));
 OAI21_X1 _791_ (.A(net94),
    .B1(_358_),
    .B2(_361_),
    .ZN(_362_));
 INV_X1 _792_ (.A(net223),
    .ZN(_363_));
 AOI21_X1 _793_ (.A(_356_),
    .B1(_362_),
    .B2(_363_),
    .ZN(_125_));
 OR2_X1 _794_ (.A1(_129_),
    .A2(net63),
    .ZN(_364_));
 NAND2_X1 _795_ (.A1(\gpio_in_sync2[8] ),
    .A2(net127),
    .ZN(_365_));
 AOI21_X1 _796_ (.A(_365_),
    .B1(net159),
    .B2(\gpio_in_prev[8] ),
    .ZN(_366_));
 OR2_X1 _797_ (.A1(\gpio_in_sync2[8] ),
    .A2(net127),
    .ZN(_367_));
 INV_X1 _798_ (.A(\gpio_in_prev[8] ),
    .ZN(_368_));
 AOI21_X1 _799_ (.A(_367_),
    .B1(net159),
    .B2(_368_),
    .ZN(_369_));
 OAI21_X1 _800_ (.A(net95),
    .B1(_366_),
    .B2(_369_),
    .ZN(_370_));
 INV_X1 _801_ (.A(net224),
    .ZN(_371_));
 AOI21_X1 _802_ (.A(_364_),
    .B1(_370_),
    .B2(_371_),
    .ZN(_126_));
 OR2_X1 _803_ (.A1(_129_),
    .A2(net64),
    .ZN(_372_));
 NAND2_X1 _804_ (.A1(\gpio_in_sync2[9] ),
    .A2(net128),
    .ZN(_373_));
 AOI21_X1 _805_ (.A(_373_),
    .B1(\gpio_in_prev[9] ),
    .B2(net160),
    .ZN(_374_));
 OR2_X1 _806_ (.A1(\gpio_in_sync2[9] ),
    .A2(net128),
    .ZN(_375_));
 INV_X1 _807_ (.A(\gpio_in_prev[9] ),
    .ZN(_376_));
 AOI21_X1 _808_ (.A(_375_),
    .B1(_376_),
    .B2(net160),
    .ZN(_377_));
 OAI21_X1 _809_ (.A(net96),
    .B1(_374_),
    .B2(_377_),
    .ZN(_378_));
 INV_X1 _810_ (.A(net225),
    .ZN(_379_));
 AOI21_X1 _811_ (.A(_372_),
    .B1(_378_),
    .B2(_379_),
    .ZN(_127_));
 BUF_X2 _812_ (.A(_128_),
    .Z(_380_));
 BUF_X2 _813_ (.A(_380_),
    .Z(_381_));
 AND2_X1 _814_ (.A1(_381_),
    .A2(\gpio_in_sync2[0] ),
    .ZN(_000_));
 AND2_X1 _815_ (.A1(_381_),
    .A2(\gpio_in_sync2[10] ),
    .ZN(_001_));
 AND2_X1 _816_ (.A1(_381_),
    .A2(\gpio_in_sync2[11] ),
    .ZN(_002_));
 AND2_X1 _817_ (.A1(_381_),
    .A2(\gpio_in_sync2[12] ),
    .ZN(_003_));
 AND2_X1 _818_ (.A1(_381_),
    .A2(\gpio_in_sync2[13] ),
    .ZN(_004_));
 AND2_X1 _819_ (.A1(_381_),
    .A2(\gpio_in_sync2[14] ),
    .ZN(_005_));
 AND2_X1 _820_ (.A1(_381_),
    .A2(\gpio_in_sync2[15] ),
    .ZN(_006_));
 AND2_X1 _821_ (.A1(_381_),
    .A2(\gpio_in_sync2[16] ),
    .ZN(_007_));
 AND2_X1 _822_ (.A1(_381_),
    .A2(\gpio_in_sync2[17] ),
    .ZN(_008_));
 AND2_X1 _823_ (.A1(_381_),
    .A2(\gpio_in_sync2[18] ),
    .ZN(_009_));
 BUF_X2 _824_ (.A(_380_),
    .Z(_382_));
 AND2_X1 _825_ (.A1(_382_),
    .A2(\gpio_in_sync2[19] ),
    .ZN(_010_));
 AND2_X1 _826_ (.A1(_382_),
    .A2(\gpio_in_sync2[1] ),
    .ZN(_011_));
 AND2_X1 _827_ (.A1(_382_),
    .A2(\gpio_in_sync2[20] ),
    .ZN(_012_));
 AND2_X1 _828_ (.A1(_382_),
    .A2(\gpio_in_sync2[21] ),
    .ZN(_013_));
 AND2_X1 _829_ (.A1(_382_),
    .A2(\gpio_in_sync2[22] ),
    .ZN(_014_));
 AND2_X1 _830_ (.A1(_382_),
    .A2(\gpio_in_sync2[23] ),
    .ZN(_015_));
 AND2_X1 _831_ (.A1(_382_),
    .A2(\gpio_in_sync2[24] ),
    .ZN(_016_));
 AND2_X1 _832_ (.A1(_382_),
    .A2(\gpio_in_sync2[25] ),
    .ZN(_017_));
 AND2_X1 _833_ (.A1(_382_),
    .A2(\gpio_in_sync2[26] ),
    .ZN(_018_));
 AND2_X1 _834_ (.A1(_382_),
    .A2(\gpio_in_sync2[27] ),
    .ZN(_019_));
 BUF_X2 _835_ (.A(_380_),
    .Z(_383_));
 AND2_X1 _836_ (.A1(_383_),
    .A2(\gpio_in_sync2[28] ),
    .ZN(_020_));
 AND2_X1 _837_ (.A1(_383_),
    .A2(\gpio_in_sync2[29] ),
    .ZN(_021_));
 AND2_X1 _838_ (.A1(_383_),
    .A2(\gpio_in_sync2[2] ),
    .ZN(_022_));
 AND2_X1 _839_ (.A1(_383_),
    .A2(\gpio_in_sync2[30] ),
    .ZN(_023_));
 AND2_X1 _840_ (.A1(_383_),
    .A2(\gpio_in_sync2[31] ),
    .ZN(_024_));
 AND2_X1 _841_ (.A1(\gpio_in_sync2[3] ),
    .A2(_380_),
    .ZN(_025_));
 AND2_X1 _842_ (.A1(_383_),
    .A2(\gpio_in_sync2[4] ),
    .ZN(_026_));
 AND2_X1 _843_ (.A1(_383_),
    .A2(\gpio_in_sync2[5] ),
    .ZN(_027_));
 AND2_X1 _844_ (.A1(_383_),
    .A2(\gpio_in_sync2[6] ),
    .ZN(_028_));
 AND2_X1 _845_ (.A1(_383_),
    .A2(\gpio_in_sync2[7] ),
    .ZN(_029_));
 AND2_X1 _846_ (.A1(_383_),
    .A2(\gpio_in_sync2[8] ),
    .ZN(_030_));
 BUF_X2 _847_ (.A(_380_),
    .Z(_384_));
 AND2_X1 _848_ (.A1(_384_),
    .A2(\gpio_in_sync2[9] ),
    .ZN(_031_));
 AND2_X1 _849_ (.A1(_384_),
    .A2(net1),
    .ZN(_032_));
 AND2_X1 _850_ (.A1(_384_),
    .A2(net2),
    .ZN(_033_));
 AND2_X1 _851_ (.A1(_384_),
    .A2(net3),
    .ZN(_034_));
 AND2_X1 _852_ (.A1(_384_),
    .A2(net4),
    .ZN(_035_));
 AND2_X1 _853_ (.A1(_384_),
    .A2(net5),
    .ZN(_036_));
 AND2_X1 _854_ (.A1(_384_),
    .A2(net6),
    .ZN(_037_));
 AND2_X1 _855_ (.A1(_384_),
    .A2(net7),
    .ZN(_038_));
 AND2_X1 _856_ (.A1(_384_),
    .A2(net8),
    .ZN(_039_));
 AND2_X1 _857_ (.A1(_384_),
    .A2(net9),
    .ZN(_040_));
 BUF_X2 _858_ (.A(_128_),
    .Z(_385_));
 AND2_X1 _859_ (.A1(_385_),
    .A2(net10),
    .ZN(_041_));
 AND2_X1 _860_ (.A1(_385_),
    .A2(net11),
    .ZN(_042_));
 AND2_X1 _861_ (.A1(_385_),
    .A2(net12),
    .ZN(_043_));
 AND2_X1 _862_ (.A1(_385_),
    .A2(net13),
    .ZN(_044_));
 AND2_X1 _863_ (.A1(_385_),
    .A2(net14),
    .ZN(_045_));
 AND2_X1 _864_ (.A1(_385_),
    .A2(net15),
    .ZN(_046_));
 AND2_X1 _865_ (.A1(_385_),
    .A2(net16),
    .ZN(_047_));
 AND2_X1 _866_ (.A1(_385_),
    .A2(net17),
    .ZN(_048_));
 AND2_X1 _867_ (.A1(_385_),
    .A2(net18),
    .ZN(_049_));
 AND2_X1 _868_ (.A1(_385_),
    .A2(net19),
    .ZN(_050_));
 BUF_X2 _869_ (.A(_128_),
    .Z(_386_));
 AND2_X1 _870_ (.A1(_386_),
    .A2(net20),
    .ZN(_051_));
 AND2_X1 _871_ (.A1(_386_),
    .A2(net21),
    .ZN(_052_));
 AND2_X1 _872_ (.A1(_386_),
    .A2(net22),
    .ZN(_053_));
 AND2_X1 _873_ (.A1(_386_),
    .A2(net23),
    .ZN(_054_));
 AND2_X1 _874_ (.A1(_386_),
    .A2(net24),
    .ZN(_055_));
 AND2_X1 _875_ (.A1(_386_),
    .A2(net25),
    .ZN(_056_));
 AND2_X1 _876_ (.A1(_386_),
    .A2(net26),
    .ZN(_057_));
 AND2_X1 _877_ (.A1(_386_),
    .A2(net27),
    .ZN(_058_));
 AND2_X1 _878_ (.A1(_386_),
    .A2(net28),
    .ZN(_059_));
 AND2_X1 _879_ (.A1(_386_),
    .A2(net29),
    .ZN(_060_));
 BUF_X2 _880_ (.A(_128_),
    .Z(_387_));
 AND2_X1 _881_ (.A1(_387_),
    .A2(net30),
    .ZN(_061_));
 AND2_X1 _882_ (.A1(_387_),
    .A2(net31),
    .ZN(_062_));
 AND2_X1 _883_ (.A1(_387_),
    .A2(net32),
    .ZN(_063_));
 AND2_X1 _884_ (.A1(_387_),
    .A2(\gpio_in_sync1[0] ),
    .ZN(_064_));
 AND2_X1 _885_ (.A1(_387_),
    .A2(\gpio_in_sync1[10] ),
    .ZN(_065_));
 AND2_X1 _886_ (.A1(_387_),
    .A2(\gpio_in_sync1[11] ),
    .ZN(_066_));
 AND2_X1 _887_ (.A1(_387_),
    .A2(\gpio_in_sync1[12] ),
    .ZN(_067_));
 AND2_X1 _888_ (.A1(_387_),
    .A2(\gpio_in_sync1[13] ),
    .ZN(_068_));
 AND2_X1 _889_ (.A1(_387_),
    .A2(\gpio_in_sync1[14] ),
    .ZN(_069_));
 AND2_X1 _890_ (.A1(_387_),
    .A2(\gpio_in_sync1[15] ),
    .ZN(_070_));
 BUF_X2 _891_ (.A(_128_),
    .Z(_388_));
 AND2_X1 _892_ (.A1(_388_),
    .A2(\gpio_in_sync1[16] ),
    .ZN(_071_));
 AND2_X1 _893_ (.A1(_388_),
    .A2(\gpio_in_sync1[17] ),
    .ZN(_072_));
 AND2_X1 _894_ (.A1(_388_),
    .A2(\gpio_in_sync1[18] ),
    .ZN(_073_));
 AND2_X1 _895_ (.A1(_388_),
    .A2(\gpio_in_sync1[19] ),
    .ZN(_074_));
 AND2_X1 _896_ (.A1(_388_),
    .A2(\gpio_in_sync1[1] ),
    .ZN(_075_));
 AND2_X1 _897_ (.A1(_388_),
    .A2(\gpio_in_sync1[20] ),
    .ZN(_076_));
 AND2_X1 _898_ (.A1(_388_),
    .A2(\gpio_in_sync1[21] ),
    .ZN(_077_));
 AND2_X1 _899_ (.A1(_388_),
    .A2(\gpio_in_sync1[22] ),
    .ZN(_078_));
 AND2_X1 _900_ (.A1(_388_),
    .A2(\gpio_in_sync1[23] ),
    .ZN(_079_));
 AND2_X1 _901_ (.A1(_388_),
    .A2(\gpio_in_sync1[24] ),
    .ZN(_080_));
 BUF_X2 _902_ (.A(_128_),
    .Z(_389_));
 AND2_X1 _903_ (.A1(_389_),
    .A2(\gpio_in_sync1[25] ),
    .ZN(_081_));
 AND2_X1 _904_ (.A1(_389_),
    .A2(\gpio_in_sync1[26] ),
    .ZN(_082_));
 AND2_X1 _905_ (.A1(_389_),
    .A2(\gpio_in_sync1[27] ),
    .ZN(_083_));
 AND2_X1 _906_ (.A1(_389_),
    .A2(\gpio_in_sync1[28] ),
    .ZN(_084_));
 AND2_X1 _907_ (.A1(_389_),
    .A2(\gpio_in_sync1[29] ),
    .ZN(_085_));
 AND2_X1 _908_ (.A1(_389_),
    .A2(\gpio_in_sync1[2] ),
    .ZN(_086_));
 AND2_X1 _909_ (.A1(_389_),
    .A2(\gpio_in_sync1[30] ),
    .ZN(_087_));
 AND2_X1 _910_ (.A1(_389_),
    .A2(\gpio_in_sync1[31] ),
    .ZN(_088_));
 AND2_X1 _911_ (.A1(_389_),
    .A2(\gpio_in_sync1[3] ),
    .ZN(_089_));
 AND2_X1 _912_ (.A1(_389_),
    .A2(\gpio_in_sync1[4] ),
    .ZN(_090_));
 AND2_X1 _913_ (.A1(_380_),
    .A2(\gpio_in_sync1[5] ),
    .ZN(_091_));
 AND2_X1 _914_ (.A1(_380_),
    .A2(\gpio_in_sync1[6] ),
    .ZN(_092_));
 AND2_X1 _915_ (.A1(_380_),
    .A2(\gpio_in_sync1[7] ),
    .ZN(_093_));
 AND2_X1 _916_ (.A1(_380_),
    .A2(\gpio_in_sync1[8] ),
    .ZN(_094_));
 AND2_X1 _917_ (.A1(_380_),
    .A2(\gpio_in_sync1[9] ),
    .ZN(_095_));
 NOR4_X1 _918_ (.A1(net202),
    .A2(net206),
    .A3(net209),
    .A4(net208),
    .ZN(_390_));
 NOR4_X2 _919_ (.A1(net201),
    .A2(net204),
    .A3(net203),
    .A4(net207),
    .ZN(_391_));
 NOR4_X1 _920_ (.A1(net211),
    .A2(net214),
    .A3(net218),
    .A4(net217),
    .ZN(_392_));
 NOR4_X1 _921_ (.A1(net210),
    .A2(net213),
    .A3(net212),
    .A4(net215),
    .ZN(_393_));
 NAND4_X1 _922_ (.A1(_390_),
    .A2(_391_),
    .A3(_392_),
    .A4(_393_),
    .ZN(_394_));
 NOR4_X1 _923_ (.A1(net221),
    .A2(net220),
    .A3(net223),
    .A4(net199),
    .ZN(_395_));
 NOR4_X2 _924_ (.A1(net205),
    .A2(net194),
    .A3(net219),
    .A4(net216),
    .ZN(_396_));
 NOR4_X1 _925_ (.A1(net222),
    .A2(net198),
    .A3(net197),
    .A4(net200),
    .ZN(_397_));
 NOR4_X1 _926_ (.A1(net225),
    .A2(net224),
    .A3(net196),
    .A4(net195),
    .ZN(_398_));
 NAND4_X1 _927_ (.A1(_395_),
    .A2(_396_),
    .A3(_397_),
    .A4(_398_),
    .ZN(_399_));
 OR2_X1 _928_ (.A1(_394_),
    .A2(_399_),
    .ZN(net193));
 BUF_X1 _929_ (.A(net1),
    .Z(net161));
 BUF_X1 _930_ (.A(net12),
    .Z(net172));
 BUF_X1 _931_ (.A(net23),
    .Z(net183));
 BUF_X1 _932_ (.A(net26),
    .Z(net186));
 BUF_X1 _933_ (.A(net27),
    .Z(net187));
 BUF_X1 _934_ (.A(net28),
    .Z(net188));
 BUF_X1 _935_ (.A(net29),
    .Z(net189));
 BUF_X1 _936_ (.A(net30),
    .Z(net190));
 BUF_X1 _937_ (.A(net31),
    .Z(net191));
 BUF_X1 _938_ (.A(net32),
    .Z(net192));
 BUF_X1 _939_ (.A(net2),
    .Z(net162));
 BUF_X1 _940_ (.A(net3),
    .Z(net163));
 BUF_X1 _941_ (.A(net4),
    .Z(net164));
 BUF_X1 _942_ (.A(net5),
    .Z(net165));
 BUF_X1 _943_ (.A(net6),
    .Z(net166));
 BUF_X1 _944_ (.A(net7),
    .Z(net167));
 BUF_X1 _945_ (.A(net8),
    .Z(net168));
 BUF_X1 _946_ (.A(net9),
    .Z(net169));
 BUF_X1 _947_ (.A(net10),
    .Z(net170));
 BUF_X1 _948_ (.A(net11),
    .Z(net171));
 BUF_X1 _949_ (.A(net13),
    .Z(net173));
 BUF_X1 _950_ (.A(net14),
    .Z(net174));
 BUF_X1 _951_ (.A(net15),
    .Z(net175));
 BUF_X1 _952_ (.A(net16),
    .Z(net176));
 BUF_X1 _953_ (.A(net17),
    .Z(net177));
 BUF_X1 _954_ (.A(net18),
    .Z(net178));
 BUF_X1 _955_ (.A(net19),
    .Z(net179));
 BUF_X1 _956_ (.A(net20),
    .Z(net180));
 BUF_X1 _957_ (.A(net21),
    .Z(net181));
 BUF_X1 _958_ (.A(net22),
    .Z(net182));
 BUF_X1 _959_ (.A(net24),
    .Z(net184));
 BUF_X1 _960_ (.A(net25),
    .Z(net185));
 BUF_X1 _961_ (.A(net1),
    .Z(gpio_pins[0]));
 BUF_X1 _962_ (.A(net12),
    .Z(gpio_pins[1]));
 BUF_X1 _963_ (.A(net23),
    .Z(gpio_pins[2]));
 BUF_X1 _964_ (.A(net26),
    .Z(gpio_pins[3]));
 BUF_X1 _965_ (.A(net27),
    .Z(gpio_pins[4]));
 BUF_X1 _966_ (.A(net28),
    .Z(gpio_pins[5]));
 BUF_X1 _967_ (.A(net29),
    .Z(gpio_pins[6]));
 BUF_X1 _968_ (.A(net30),
    .Z(gpio_pins[7]));
 BUF_X1 _969_ (.A(net31),
    .Z(gpio_pins[8]));
 BUF_X1 _970_ (.A(net32),
    .Z(gpio_pins[9]));
 BUF_X1 _971_ (.A(net2),
    .Z(gpio_pins[10]));
 BUF_X1 _972_ (.A(net3),
    .Z(gpio_pins[11]));
 BUF_X1 _973_ (.A(net4),
    .Z(gpio_pins[12]));
 BUF_X1 _974_ (.A(net5),
    .Z(gpio_pins[13]));
 BUF_X1 _975_ (.A(net6),
    .Z(gpio_pins[14]));
 BUF_X1 _976_ (.A(net7),
    .Z(gpio_pins[15]));
 BUF_X1 _977_ (.A(net8),
    .Z(gpio_pins[16]));
 BUF_X1 _978_ (.A(net9),
    .Z(gpio_pins[17]));
 BUF_X1 _979_ (.A(net10),
    .Z(gpio_pins[18]));
 BUF_X1 _980_ (.A(net11),
    .Z(gpio_pins[19]));
 BUF_X1 _981_ (.A(net13),
    .Z(gpio_pins[20]));
 BUF_X1 _982_ (.A(net14),
    .Z(gpio_pins[21]));
 BUF_X1 _983_ (.A(net15),
    .Z(gpio_pins[22]));
 BUF_X1 _984_ (.A(net16),
    .Z(gpio_pins[23]));
 BUF_X1 _985_ (.A(net17),
    .Z(gpio_pins[24]));
 BUF_X1 _986_ (.A(net18),
    .Z(gpio_pins[25]));
 BUF_X1 _987_ (.A(net19),
    .Z(gpio_pins[26]));
 BUF_X1 _988_ (.A(net20),
    .Z(gpio_pins[27]));
 BUF_X1 _989_ (.A(net21),
    .Z(gpio_pins[28]));
 BUF_X1 _990_ (.A(net22),
    .Z(gpio_pins[29]));
 BUF_X1 _991_ (.A(net24),
    .Z(gpio_pins[30]));
 BUF_X1 _992_ (.A(net25),
    .Z(gpio_pins[31]));
 DFF_X1 \gpio_in_prev[0]$_SDFF_PN0_  (.D(_000_),
    .CK(clknet_4_14_0_clk),
    .Q(\gpio_in_prev[0] ),
    .QN(_527_));
 DFF_X1 \gpio_in_prev[10]$_SDFF_PN0_  (.D(_001_),
    .CK(clknet_4_10_0_clk),
    .Q(\gpio_in_prev[10] ),
    .QN(_526_));
 DFF_X1 \gpio_in_prev[11]$_SDFF_PN0_  (.D(_002_),
    .CK(clknet_4_10_0_clk),
    .Q(\gpio_in_prev[11] ),
    .QN(_525_));
 DFF_X1 \gpio_in_prev[12]$_SDFF_PN0_  (.D(_003_),
    .CK(clknet_4_11_0_clk),
    .Q(\gpio_in_prev[12] ),
    .QN(_524_));
 DFF_X1 \gpio_in_prev[13]$_SDFF_PN0_  (.D(_004_),
    .CK(clknet_4_14_0_clk),
    .Q(\gpio_in_prev[13] ),
    .QN(_523_));
 DFF_X1 \gpio_in_prev[14]$_SDFF_PN0_  (.D(_005_),
    .CK(clknet_4_15_0_clk),
    .Q(\gpio_in_prev[14] ),
    .QN(_522_));
 DFF_X1 \gpio_in_prev[15]$_SDFF_PN0_  (.D(_006_),
    .CK(clknet_4_10_0_clk),
    .Q(\gpio_in_prev[15] ),
    .QN(_521_));
 DFF_X1 \gpio_in_prev[16]$_SDFF_PN0_  (.D(_007_),
    .CK(clknet_4_8_0_clk),
    .Q(\gpio_in_prev[16] ),
    .QN(_520_));
 DFF_X1 \gpio_in_prev[17]$_SDFF_PN0_  (.D(_008_),
    .CK(clknet_4_9_0_clk),
    .Q(\gpio_in_prev[17] ),
    .QN(_519_));
 DFF_X1 \gpio_in_prev[18]$_SDFF_PN0_  (.D(_009_),
    .CK(clknet_4_8_0_clk),
    .Q(\gpio_in_prev[18] ),
    .QN(_518_));
 DFF_X1 \gpio_in_prev[19]$_SDFF_PN0_  (.D(_010_),
    .CK(clknet_4_2_0_clk),
    .Q(\gpio_in_prev[19] ),
    .QN(_517_));
 DFF_X1 \gpio_in_prev[1]$_SDFF_PN0_  (.D(_011_),
    .CK(clknet_4_6_0_clk),
    .Q(\gpio_in_prev[1] ),
    .QN(_516_));
 DFF_X1 \gpio_in_prev[20]$_SDFF_PN0_  (.D(_012_),
    .CK(clknet_4_1_0_clk),
    .Q(\gpio_in_prev[20] ),
    .QN(_515_));
 DFF_X1 \gpio_in_prev[21]$_SDFF_PN0_  (.D(_013_),
    .CK(clknet_4_3_0_clk),
    .Q(\gpio_in_prev[21] ),
    .QN(_514_));
 DFF_X1 \gpio_in_prev[22]$_SDFF_PN0_  (.D(_014_),
    .CK(clknet_4_0_0_clk),
    .Q(\gpio_in_prev[22] ),
    .QN(_513_));
 DFF_X1 \gpio_in_prev[23]$_SDFF_PN0_  (.D(_015_),
    .CK(clknet_4_0_0_clk),
    .Q(\gpio_in_prev[23] ),
    .QN(_512_));
 DFF_X1 \gpio_in_prev[24]$_SDFF_PN0_  (.D(_016_),
    .CK(clknet_4_1_0_clk),
    .Q(\gpio_in_prev[24] ),
    .QN(_511_));
 DFF_X1 \gpio_in_prev[25]$_SDFF_PN0_  (.D(_017_),
    .CK(clknet_4_6_0_clk),
    .Q(\gpio_in_prev[25] ),
    .QN(_510_));
 DFF_X1 \gpio_in_prev[26]$_SDFF_PN0_  (.D(_018_),
    .CK(clknet_4_4_0_clk),
    .Q(\gpio_in_prev[26] ),
    .QN(_509_));
 DFF_X1 \gpio_in_prev[27]$_SDFF_PN0_  (.D(_019_),
    .CK(clknet_4_5_0_clk),
    .Q(\gpio_in_prev[27] ),
    .QN(_508_));
 DFF_X1 \gpio_in_prev[28]$_SDFF_PN0_  (.D(_020_),
    .CK(clknet_4_5_0_clk),
    .Q(\gpio_in_prev[28] ),
    .QN(_507_));
 DFF_X1 \gpio_in_prev[29]$_SDFF_PN0_  (.D(_021_),
    .CK(clknet_4_7_0_clk),
    .Q(\gpio_in_prev[29] ),
    .QN(_506_));
 DFF_X1 \gpio_in_prev[2]$_SDFF_PN0_  (.D(_022_),
    .CK(clknet_4_13_0_clk),
    .Q(\gpio_in_prev[2] ),
    .QN(_505_));
 DFF_X1 \gpio_in_prev[30]$_SDFF_PN0_  (.D(_023_),
    .CK(clknet_4_7_0_clk),
    .Q(\gpio_in_prev[30] ),
    .QN(_504_));
 DFF_X1 \gpio_in_prev[31]$_SDFF_PN0_  (.D(_024_),
    .CK(clknet_4_5_0_clk),
    .Q(\gpio_in_prev[31] ),
    .QN(_503_));
 DFF_X1 \gpio_in_prev[3]$_SDFF_PN0_  (.D(_025_),
    .CK(clknet_4_7_0_clk),
    .Q(\gpio_in_prev[3] ),
    .QN(_502_));
 DFF_X1 \gpio_in_prev[4]$_SDFF_PN0_  (.D(_026_),
    .CK(clknet_4_7_0_clk),
    .Q(\gpio_in_prev[4] ),
    .QN(_501_));
 DFF_X1 \gpio_in_prev[5]$_SDFF_PN0_  (.D(_027_),
    .CK(clknet_4_13_0_clk),
    .Q(\gpio_in_prev[5] ),
    .QN(_500_));
 DFF_X1 \gpio_in_prev[6]$_SDFF_PN0_  (.D(_028_),
    .CK(clknet_4_15_0_clk),
    .Q(\gpio_in_prev[6] ),
    .QN(_499_));
 DFF_X1 \gpio_in_prev[7]$_SDFF_PN0_  (.D(_029_),
    .CK(clknet_4_15_0_clk),
    .Q(\gpio_in_prev[7] ),
    .QN(_498_));
 DFF_X1 \gpio_in_prev[8]$_SDFF_PN0_  (.D(_030_),
    .CK(clknet_4_15_0_clk),
    .Q(\gpio_in_prev[8] ),
    .QN(_497_));
 DFF_X1 \gpio_in_prev[9]$_SDFF_PN0_  (.D(_031_),
    .CK(clknet_4_11_0_clk),
    .Q(\gpio_in_prev[9] ),
    .QN(_496_));
 DFF_X1 \gpio_in_sync1[0]$_SDFF_PN0_  (.D(_032_),
    .CK(clknet_4_9_0_clk),
    .Q(\gpio_in_sync1[0] ),
    .QN(_495_));
 DFF_X1 \gpio_in_sync1[10]$_SDFF_PN0_  (.D(_033_),
    .CK(clknet_4_10_0_clk),
    .Q(\gpio_in_sync1[10] ),
    .QN(_494_));
 DFF_X1 \gpio_in_sync1[11]$_SDFF_PN0_  (.D(_034_),
    .CK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync1[11] ),
    .QN(_493_));
 DFF_X1 \gpio_in_sync1[12]$_SDFF_PN0_  (.D(_035_),
    .CK(clknet_4_10_0_clk),
    .Q(\gpio_in_sync1[12] ),
    .QN(_492_));
 DFF_X1 \gpio_in_sync1[13]$_SDFF_PN0_  (.D(_036_),
    .CK(clknet_4_11_0_clk),
    .Q(\gpio_in_sync1[13] ),
    .QN(_491_));
 DFF_X1 \gpio_in_sync1[14]$_SDFF_PN0_  (.D(_037_),
    .CK(clknet_4_14_0_clk),
    .Q(\gpio_in_sync1[14] ),
    .QN(_490_));
 DFF_X1 \gpio_in_sync1[15]$_SDFF_PN0_  (.D(_038_),
    .CK(clknet_4_10_0_clk),
    .Q(\gpio_in_sync1[15] ),
    .QN(_489_));
 DFF_X1 \gpio_in_sync1[16]$_SDFF_PN0_  (.D(_039_),
    .CK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync1[16] ),
    .QN(_488_));
 DFF_X1 \gpio_in_sync1[17]$_SDFF_PN0_  (.D(_040_),
    .CK(clknet_4_9_0_clk),
    .Q(\gpio_in_sync1[17] ),
    .QN(_487_));
 DFF_X1 \gpio_in_sync1[18]$_SDFF_PN0_  (.D(_041_),
    .CK(clknet_4_2_0_clk),
    .Q(\gpio_in_sync1[18] ),
    .QN(_486_));
 DFF_X1 \gpio_in_sync1[19]$_SDFF_PN0_  (.D(_042_),
    .CK(clknet_4_3_0_clk),
    .Q(\gpio_in_sync1[19] ),
    .QN(_485_));
 DFF_X1 \gpio_in_sync1[1]$_SDFF_PN0_  (.D(_043_),
    .CK(clknet_4_3_0_clk),
    .Q(\gpio_in_sync1[1] ),
    .QN(_484_));
 DFF_X1 \gpio_in_sync1[20]$_SDFF_PN0_  (.D(_044_),
    .CK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync1[20] ),
    .QN(_483_));
 DFF_X1 \gpio_in_sync1[21]$_SDFF_PN0_  (.D(_045_),
    .CK(clknet_4_3_0_clk),
    .Q(\gpio_in_sync1[21] ),
    .QN(_482_));
 DFF_X1 \gpio_in_sync1[22]$_SDFF_PN0_  (.D(_046_),
    .CK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync1[22] ),
    .QN(_481_));
 DFF_X1 \gpio_in_sync1[23]$_SDFF_PN0_  (.D(_047_),
    .CK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync1[23] ),
    .QN(_480_));
 DFF_X1 \gpio_in_sync1[24]$_SDFF_PN0_  (.D(_048_),
    .CK(clknet_4_1_0_clk),
    .Q(\gpio_in_sync1[24] ),
    .QN(_479_));
 DFF_X1 \gpio_in_sync1[25]$_SDFF_PN0_  (.D(_049_),
    .CK(clknet_4_1_0_clk),
    .Q(\gpio_in_sync1[25] ),
    .QN(_478_));
 DFF_X1 \gpio_in_sync1[26]$_SDFF_PN0_  (.D(_050_),
    .CK(clknet_4_1_0_clk),
    .Q(\gpio_in_sync1[26] ),
    .QN(_477_));
 DFF_X1 \gpio_in_sync1[27]$_SDFF_PN0_  (.D(_051_),
    .CK(clknet_4_4_0_clk),
    .Q(\gpio_in_sync1[27] ),
    .QN(_476_));
 DFF_X1 \gpio_in_sync1[28]$_SDFF_PN0_  (.D(_052_),
    .CK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync1[28] ),
    .QN(_475_));
 DFF_X1 \gpio_in_sync1[29]$_SDFF_PN0_  (.D(_053_),
    .CK(clknet_4_4_0_clk),
    .Q(\gpio_in_sync1[29] ),
    .QN(_474_));
 DFF_X1 \gpio_in_sync1[2]$_SDFF_PN0_  (.D(_054_),
    .CK(clknet_4_6_0_clk),
    .Q(\gpio_in_sync1[2] ),
    .QN(_473_));
 DFF_X1 \gpio_in_sync1[30]$_SDFF_PN0_  (.D(_055_),
    .CK(clknet_4_7_0_clk),
    .Q(\gpio_in_sync1[30] ),
    .QN(_472_));
 DFF_X1 \gpio_in_sync1[31]$_SDFF_PN0_  (.D(_056_),
    .CK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync1[31] ),
    .QN(_471_));
 DFF_X1 \gpio_in_sync1[3]$_SDFF_PN0_  (.D(_057_),
    .CK(clknet_4_6_0_clk),
    .Q(\gpio_in_sync1[3] ),
    .QN(_470_));
 DFF_X1 \gpio_in_sync1[4]$_SDFF_PN0_  (.D(_058_),
    .CK(clknet_4_7_0_clk),
    .Q(\gpio_in_sync1[4] ),
    .QN(_469_));
 DFF_X1 \gpio_in_sync1[5]$_SDFF_PN0_  (.D(_059_),
    .CK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync1[5] ),
    .QN(_468_));
 DFF_X1 \gpio_in_sync1[6]$_SDFF_PN0_  (.D(_060_),
    .CK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync1[6] ),
    .QN(_467_));
 DFF_X1 \gpio_in_sync1[7]$_SDFF_PN0_  (.D(_061_),
    .CK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync1[7] ),
    .QN(_466_));
 DFF_X1 \gpio_in_sync1[8]$_SDFF_PN0_  (.D(_062_),
    .CK(clknet_4_14_0_clk),
    .Q(\gpio_in_sync1[8] ),
    .QN(_465_));
 DFF_X1 \gpio_in_sync1[9]$_SDFF_PN0_  (.D(_063_),
    .CK(clknet_4_9_0_clk),
    .Q(\gpio_in_sync1[9] ),
    .QN(_464_));
 DFF_X1 \gpio_in_sync2[0]$_SDFF_PN0_  (.D(_064_),
    .CK(clknet_4_9_0_clk),
    .Q(\gpio_in_sync2[0] ),
    .QN(_463_));
 DFF_X1 \gpio_in_sync2[10]$_SDFF_PN0_  (.D(_065_),
    .CK(clknet_4_10_0_clk),
    .Q(\gpio_in_sync2[10] ),
    .QN(_462_));
 DFF_X1 \gpio_in_sync2[11]$_SDFF_PN0_  (.D(_066_),
    .CK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync2[11] ),
    .QN(_461_));
 DFF_X1 \gpio_in_sync2[12]$_SDFF_PN0_  (.D(_067_),
    .CK(clknet_4_10_0_clk),
    .Q(\gpio_in_sync2[12] ),
    .QN(_460_));
 DFF_X1 \gpio_in_sync2[13]$_SDFF_PN0_  (.D(_068_),
    .CK(clknet_4_14_0_clk),
    .Q(\gpio_in_sync2[13] ),
    .QN(_459_));
 DFF_X1 \gpio_in_sync2[14]$_SDFF_PN0_  (.D(_069_),
    .CK(clknet_4_14_0_clk),
    .Q(\gpio_in_sync2[14] ),
    .QN(_458_));
 DFF_X1 \gpio_in_sync2[15]$_SDFF_PN0_  (.D(_070_),
    .CK(clknet_4_10_0_clk),
    .Q(\gpio_in_sync2[15] ),
    .QN(_457_));
 DFF_X1 \gpio_in_sync2[16]$_SDFF_PN0_  (.D(_071_),
    .CK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync2[16] ),
    .QN(_456_));
 DFF_X1 \gpio_in_sync2[17]$_SDFF_PN0_  (.D(_072_),
    .CK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync2[17] ),
    .QN(_455_));
 DFF_X1 \gpio_in_sync2[18]$_SDFF_PN0_  (.D(_073_),
    .CK(clknet_4_3_0_clk),
    .Q(\gpio_in_sync2[18] ),
    .QN(_454_));
 DFF_X1 \gpio_in_sync2[19]$_SDFF_PN0_  (.D(_074_),
    .CK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync2[19] ),
    .QN(_453_));
 DFF_X1 \gpio_in_sync2[1]$_SDFF_PN0_  (.D(_075_),
    .CK(clknet_4_2_0_clk),
    .Q(\gpio_in_sync2[1] ),
    .QN(_452_));
 DFF_X1 \gpio_in_sync2[20]$_SDFF_PN0_  (.D(_076_),
    .CK(clknet_4_1_0_clk),
    .Q(\gpio_in_sync2[20] ),
    .QN(_451_));
 DFF_X1 \gpio_in_sync2[21]$_SDFF_PN0_  (.D(_077_),
    .CK(clknet_4_3_0_clk),
    .Q(\gpio_in_sync2[21] ),
    .QN(_450_));
 DFF_X1 \gpio_in_sync2[22]$_SDFF_PN0_  (.D(_078_),
    .CK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync2[22] ),
    .QN(_449_));
 DFF_X1 \gpio_in_sync2[23]$_SDFF_PN0_  (.D(_079_),
    .CK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync2[23] ),
    .QN(_448_));
 DFF_X1 \gpio_in_sync2[24]$_SDFF_PN0_  (.D(_080_),
    .CK(clknet_4_1_0_clk),
    .Q(\gpio_in_sync2[24] ),
    .QN(_447_));
 DFF_X1 \gpio_in_sync2[25]$_SDFF_PN0_  (.D(_081_),
    .CK(clknet_4_4_0_clk),
    .Q(\gpio_in_sync2[25] ),
    .QN(_446_));
 DFF_X1 \gpio_in_sync2[26]$_SDFF_PN0_  (.D(_082_),
    .CK(clknet_4_4_0_clk),
    .Q(\gpio_in_sync2[26] ),
    .QN(_445_));
 DFF_X1 \gpio_in_sync2[27]$_SDFF_PN0_  (.D(_083_),
    .CK(clknet_4_4_0_clk),
    .Q(\gpio_in_sync2[27] ),
    .QN(_444_));
 DFF_X1 \gpio_in_sync2[28]$_SDFF_PN0_  (.D(_084_),
    .CK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync2[28] ),
    .QN(_443_));
 DFF_X1 \gpio_in_sync2[29]$_SDFF_PN0_  (.D(_085_),
    .CK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync2[29] ),
    .QN(_442_));
 DFF_X1 \gpio_in_sync2[2]$_SDFF_PN0_  (.D(_086_),
    .CK(clknet_4_13_0_clk),
    .Q(\gpio_in_sync2[2] ),
    .QN(_441_));
 DFF_X1 \gpio_in_sync2[30]$_SDFF_PN0_  (.D(_087_),
    .CK(clknet_4_7_0_clk),
    .Q(\gpio_in_sync2[30] ),
    .QN(_440_));
 DFF_X1 \gpio_in_sync2[31]$_SDFF_PN0_  (.D(_088_),
    .CK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync2[31] ),
    .QN(_439_));
 DFF_X1 \gpio_in_sync2[3]$_SDFF_PN0_  (.D(_089_),
    .CK(clknet_4_6_0_clk),
    .Q(\gpio_in_sync2[3] ),
    .QN(_438_));
 DFF_X1 \gpio_in_sync2[4]$_SDFF_PN0_  (.D(_090_),
    .CK(clknet_4_7_0_clk),
    .Q(\gpio_in_sync2[4] ),
    .QN(_437_));
 DFF_X1 \gpio_in_sync2[5]$_SDFF_PN0_  (.D(_091_),
    .CK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync2[5] ),
    .QN(_436_));
 DFF_X1 \gpio_in_sync2[6]$_SDFF_PN0_  (.D(_092_),
    .CK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync2[6] ),
    .QN(_435_));
 DFF_X1 \gpio_in_sync2[7]$_SDFF_PN0_  (.D(_093_),
    .CK(clknet_4_15_0_clk),
    .Q(\gpio_in_sync2[7] ),
    .QN(_434_));
 DFF_X1 \gpio_in_sync2[8]$_SDFF_PN0_  (.D(_094_),
    .CK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync2[8] ),
    .QN(_433_));
 DFF_X1 \gpio_in_sync2[9]$_SDFF_PN0_  (.D(_095_),
    .CK(clknet_4_11_0_clk),
    .Q(\gpio_in_sync2[9] ),
    .QN(_432_));
 DFF_X1 \int_status_reg[0]$_SDFFE_PP0P_  (.D(_096_),
    .CK(clknet_4_15_0_clk),
    .Q(net194),
    .QN(_431_));
 DFF_X1 \int_status_reg[10]$_SDFFE_PP0P_  (.D(_097_),
    .CK(clknet_4_11_0_clk),
    .Q(net195),
    .QN(_430_));
 DFF_X1 \int_status_reg[11]$_SDFFE_PP0P_  (.D(_098_),
    .CK(clknet_4_10_0_clk),
    .Q(net196),
    .QN(_429_));
 DFF_X1 \int_status_reg[12]$_SDFFE_PP0P_  (.D(_099_),
    .CK(clknet_4_11_0_clk),
    .Q(net197),
    .QN(_428_));
 DFF_X1 \int_status_reg[13]$_SDFFE_PP0P_  (.D(_100_),
    .CK(clknet_4_11_0_clk),
    .Q(net198),
    .QN(_427_));
 DFF_X1 \int_status_reg[14]$_SDFFE_PP0P_  (.D(_101_),
    .CK(clknet_4_15_0_clk),
    .Q(net199),
    .QN(_426_));
 DFF_X1 \int_status_reg[15]$_SDFFE_PP0P_  (.D(_102_),
    .CK(clknet_4_11_0_clk),
    .Q(net200),
    .QN(_425_));
 DFF_X1 \int_status_reg[16]$_SDFFE_PP0P_  (.D(_103_),
    .CK(clknet_4_8_0_clk),
    .Q(net201),
    .QN(_424_));
 DFF_X1 \int_status_reg[17]$_SDFFE_PP0P_  (.D(_104_),
    .CK(clknet_4_3_0_clk),
    .Q(net202),
    .QN(_423_));
 DFF_X1 \int_status_reg[18]$_SDFFE_PP0P_  (.D(_105_),
    .CK(clknet_4_2_0_clk),
    .Q(net203),
    .QN(_422_));
 DFF_X1 \int_status_reg[19]$_SDFFE_PP0P_  (.D(_106_),
    .CK(clknet_4_2_0_clk),
    .Q(net204),
    .QN(_421_));
 DFF_X1 \int_status_reg[1]$_SDFFE_PP0P_  (.D(_107_),
    .CK(clknet_4_13_0_clk),
    .Q(net205),
    .QN(_420_));
 DFF_X1 \int_status_reg[20]$_SDFFE_PP0P_  (.D(_108_),
    .CK(clknet_4_0_0_clk),
    .Q(net206),
    .QN(_419_));
 DFF_X1 \int_status_reg[21]$_SDFFE_PP0P_  (.D(_109_),
    .CK(clknet_4_2_0_clk),
    .Q(net207),
    .QN(_418_));
 DFF_X1 \int_status_reg[22]$_SDFFE_PP0P_  (.D(_110_),
    .CK(clknet_4_0_0_clk),
    .Q(net208),
    .QN(_417_));
 DFF_X1 \int_status_reg[23]$_SDFFE_PP0P_  (.D(_111_),
    .CK(clknet_4_0_0_clk),
    .Q(net209),
    .QN(_416_));
 DFF_X1 \int_status_reg[24]$_SDFFE_PP0P_  (.D(_112_),
    .CK(clknet_4_1_0_clk),
    .Q(net210),
    .QN(_415_));
 DFF_X1 \int_status_reg[25]$_SDFFE_PP0P_  (.D(_113_),
    .CK(clknet_4_6_0_clk),
    .Q(net211),
    .QN(_414_));
 DFF_X1 \int_status_reg[26]$_SDFFE_PP0P_  (.D(_114_),
    .CK(clknet_4_4_0_clk),
    .Q(net212),
    .QN(_413_));
 DFF_X1 \int_status_reg[27]$_SDFFE_PP0P_  (.D(_115_),
    .CK(clknet_4_4_0_clk),
    .Q(net213),
    .QN(_412_));
 DFF_X1 \int_status_reg[28]$_SDFFE_PP0P_  (.D(_116_),
    .CK(clknet_4_5_0_clk),
    .Q(net214),
    .QN(_411_));
 DFF_X1 \int_status_reg[29]$_SDFFE_PP0P_  (.D(_117_),
    .CK(clknet_4_6_0_clk),
    .Q(net215),
    .QN(_410_));
 DFF_X1 \int_status_reg[2]$_SDFFE_PP0P_  (.D(_118_),
    .CK(clknet_4_13_0_clk),
    .Q(net216),
    .QN(_409_));
 DFF_X1 \int_status_reg[30]$_SDFFE_PP0P_  (.D(_119_),
    .CK(clknet_4_7_0_clk),
    .Q(net217),
    .QN(_408_));
 DFF_X1 \int_status_reg[31]$_SDFFE_PP0P_  (.D(_120_),
    .CK(clknet_4_5_0_clk),
    .Q(net218),
    .QN(_407_));
 DFF_X1 \int_status_reg[3]$_SDFFE_PP0P_  (.D(_121_),
    .CK(clknet_4_13_0_clk),
    .Q(net219),
    .QN(_406_));
 DFF_X1 \int_status_reg[4]$_SDFFE_PP0P_  (.D(_122_),
    .CK(clknet_4_13_0_clk),
    .Q(net220),
    .QN(_405_));
 DFF_X1 \int_status_reg[5]$_SDFFE_PP0P_  (.D(_123_),
    .CK(clknet_4_15_0_clk),
    .Q(net221),
    .QN(_404_));
 DFF_X1 \int_status_reg[6]$_SDFFE_PP0P_  (.D(_124_),
    .CK(clknet_4_15_0_clk),
    .Q(net222),
    .QN(_403_));
 DFF_X1 \int_status_reg[7]$_SDFFE_PP0P_  (.D(_125_),
    .CK(clknet_4_15_0_clk),
    .Q(net223),
    .QN(_402_));
 DFF_X1 \int_status_reg[8]$_SDFFE_PP0P_  (.D(_126_),
    .CK(clknet_4_14_0_clk),
    .Q(net224),
    .QN(_401_));
 DFF_X1 \int_status_reg[9]$_SDFFE_PP0P_  (.D(_127_),
    .CK(clknet_4_14_0_clk),
    .Q(net225),
    .QN(_400_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_63 ();
 BUF_X1 input1 (.A(gpio_out[0]),
    .Z(net1));
 BUF_X1 input2 (.A(gpio_out[10]),
    .Z(net2));
 BUF_X1 input3 (.A(gpio_out[11]),
    .Z(net3));
 BUF_X1 input4 (.A(gpio_out[12]),
    .Z(net4));
 BUF_X1 input5 (.A(gpio_out[13]),
    .Z(net5));
 BUF_X1 input6 (.A(gpio_out[14]),
    .Z(net6));
 BUF_X1 input7 (.A(gpio_out[15]),
    .Z(net7));
 BUF_X1 input8 (.A(gpio_out[16]),
    .Z(net8));
 BUF_X1 input9 (.A(gpio_out[17]),
    .Z(net9));
 BUF_X1 input10 (.A(gpio_out[18]),
    .Z(net10));
 BUF_X1 input11 (.A(gpio_out[19]),
    .Z(net11));
 BUF_X1 input12 (.A(gpio_out[1]),
    .Z(net12));
 BUF_X1 input13 (.A(gpio_out[20]),
    .Z(net13));
 BUF_X1 input14 (.A(gpio_out[21]),
    .Z(net14));
 BUF_X1 input15 (.A(gpio_out[22]),
    .Z(net15));
 BUF_X1 input16 (.A(gpio_out[23]),
    .Z(net16));
 BUF_X1 input17 (.A(gpio_out[24]),
    .Z(net17));
 BUF_X1 input18 (.A(gpio_out[25]),
    .Z(net18));
 BUF_X1 input19 (.A(gpio_out[26]),
    .Z(net19));
 BUF_X1 input20 (.A(gpio_out[27]),
    .Z(net20));
 BUF_X1 input21 (.A(gpio_out[28]),
    .Z(net21));
 BUF_X1 input22 (.A(gpio_out[29]),
    .Z(net22));
 BUF_X1 input23 (.A(gpio_out[2]),
    .Z(net23));
 BUF_X1 input24 (.A(gpio_out[30]),
    .Z(net24));
 BUF_X1 input25 (.A(gpio_out[31]),
    .Z(net25));
 BUF_X1 input26 (.A(gpio_out[3]),
    .Z(net26));
 BUF_X1 input27 (.A(gpio_out[4]),
    .Z(net27));
 BUF_X1 input28 (.A(gpio_out[5]),
    .Z(net28));
 BUF_X1 input29 (.A(gpio_out[6]),
    .Z(net29));
 BUF_X1 input30 (.A(gpio_out[7]),
    .Z(net30));
 BUF_X1 input31 (.A(gpio_out[8]),
    .Z(net31));
 BUF_X1 input32 (.A(gpio_out[9]),
    .Z(net32));
 BUF_X1 input33 (.A(int_clear[0]),
    .Z(net33));
 BUF_X1 input34 (.A(int_clear[10]),
    .Z(net34));
 BUF_X1 input35 (.A(int_clear[11]),
    .Z(net35));
 BUF_X1 input36 (.A(int_clear[12]),
    .Z(net36));
 BUF_X1 input37 (.A(int_clear[13]),
    .Z(net37));
 BUF_X1 input38 (.A(int_clear[14]),
    .Z(net38));
 BUF_X1 input39 (.A(int_clear[15]),
    .Z(net39));
 BUF_X1 input40 (.A(int_clear[16]),
    .Z(net40));
 BUF_X1 input41 (.A(int_clear[17]),
    .Z(net41));
 BUF_X1 input42 (.A(int_clear[18]),
    .Z(net42));
 BUF_X1 input43 (.A(int_clear[19]),
    .Z(net43));
 BUF_X1 input44 (.A(int_clear[1]),
    .Z(net44));
 BUF_X1 input45 (.A(int_clear[20]),
    .Z(net45));
 BUF_X1 input46 (.A(int_clear[21]),
    .Z(net46));
 BUF_X1 input47 (.A(int_clear[22]),
    .Z(net47));
 BUF_X1 input48 (.A(int_clear[23]),
    .Z(net48));
 BUF_X1 input49 (.A(int_clear[24]),
    .Z(net49));
 BUF_X1 input50 (.A(int_clear[25]),
    .Z(net50));
 BUF_X1 input51 (.A(int_clear[26]),
    .Z(net51));
 BUF_X1 input52 (.A(int_clear[27]),
    .Z(net52));
 BUF_X1 input53 (.A(int_clear[28]),
    .Z(net53));
 BUF_X1 input54 (.A(int_clear[29]),
    .Z(net54));
 BUF_X1 input55 (.A(int_clear[2]),
    .Z(net55));
 BUF_X1 input56 (.A(int_clear[30]),
    .Z(net56));
 BUF_X1 input57 (.A(int_clear[31]),
    .Z(net57));
 BUF_X1 input58 (.A(int_clear[3]),
    .Z(net58));
 BUF_X1 input59 (.A(int_clear[4]),
    .Z(net59));
 BUF_X1 input60 (.A(int_clear[5]),
    .Z(net60));
 BUF_X1 input61 (.A(int_clear[6]),
    .Z(net61));
 BUF_X1 input62 (.A(int_clear[7]),
    .Z(net62));
 BUF_X1 input63 (.A(int_clear[8]),
    .Z(net63));
 BUF_X1 input64 (.A(int_clear[9]),
    .Z(net64));
 BUF_X1 input65 (.A(int_enable[0]),
    .Z(net65));
 BUF_X1 input66 (.A(int_enable[10]),
    .Z(net66));
 BUF_X1 input67 (.A(int_enable[11]),
    .Z(net67));
 BUF_X1 input68 (.A(int_enable[12]),
    .Z(net68));
 BUF_X1 input69 (.A(int_enable[13]),
    .Z(net69));
 BUF_X1 input70 (.A(int_enable[14]),
    .Z(net70));
 BUF_X1 input71 (.A(int_enable[15]),
    .Z(net71));
 BUF_X1 input72 (.A(int_enable[16]),
    .Z(net72));
 BUF_X1 input73 (.A(int_enable[17]),
    .Z(net73));
 BUF_X1 input74 (.A(int_enable[18]),
    .Z(net74));
 BUF_X1 input75 (.A(int_enable[19]),
    .Z(net75));
 BUF_X1 input76 (.A(int_enable[1]),
    .Z(net76));
 BUF_X1 input77 (.A(int_enable[20]),
    .Z(net77));
 BUF_X1 input78 (.A(int_enable[21]),
    .Z(net78));
 BUF_X1 input79 (.A(int_enable[22]),
    .Z(net79));
 BUF_X1 input80 (.A(int_enable[23]),
    .Z(net80));
 BUF_X1 input81 (.A(int_enable[24]),
    .Z(net81));
 BUF_X1 input82 (.A(int_enable[25]),
    .Z(net82));
 BUF_X1 input83 (.A(int_enable[26]),
    .Z(net83));
 BUF_X1 input84 (.A(int_enable[27]),
    .Z(net84));
 BUF_X1 input85 (.A(int_enable[28]),
    .Z(net85));
 BUF_X1 input86 (.A(int_enable[29]),
    .Z(net86));
 BUF_X1 input87 (.A(int_enable[2]),
    .Z(net87));
 BUF_X1 input88 (.A(int_enable[30]),
    .Z(net88));
 BUF_X1 input89 (.A(int_enable[31]),
    .Z(net89));
 BUF_X1 input90 (.A(int_enable[3]),
    .Z(net90));
 BUF_X1 input91 (.A(int_enable[4]),
    .Z(net91));
 BUF_X1 input92 (.A(int_enable[5]),
    .Z(net92));
 BUF_X1 input93 (.A(int_enable[6]),
    .Z(net93));
 BUF_X1 input94 (.A(int_enable[7]),
    .Z(net94));
 BUF_X1 input95 (.A(int_enable[8]),
    .Z(net95));
 BUF_X1 input96 (.A(int_enable[9]),
    .Z(net96));
 BUF_X1 input97 (.A(int_polarity[0]),
    .Z(net97));
 BUF_X1 input98 (.A(int_polarity[10]),
    .Z(net98));
 BUF_X1 input99 (.A(int_polarity[11]),
    .Z(net99));
 BUF_X1 input100 (.A(int_polarity[12]),
    .Z(net100));
 BUF_X1 input101 (.A(int_polarity[13]),
    .Z(net101));
 BUF_X1 input102 (.A(int_polarity[14]),
    .Z(net102));
 BUF_X1 input103 (.A(int_polarity[15]),
    .Z(net103));
 BUF_X1 input104 (.A(int_polarity[16]),
    .Z(net104));
 BUF_X1 input105 (.A(int_polarity[17]),
    .Z(net105));
 BUF_X1 input106 (.A(int_polarity[18]),
    .Z(net106));
 BUF_X1 input107 (.A(int_polarity[19]),
    .Z(net107));
 BUF_X1 input108 (.A(int_polarity[1]),
    .Z(net108));
 BUF_X1 input109 (.A(int_polarity[20]),
    .Z(net109));
 BUF_X1 input110 (.A(int_polarity[21]),
    .Z(net110));
 BUF_X1 input111 (.A(int_polarity[22]),
    .Z(net111));
 BUF_X1 input112 (.A(int_polarity[23]),
    .Z(net112));
 BUF_X1 input113 (.A(int_polarity[24]),
    .Z(net113));
 BUF_X1 input114 (.A(int_polarity[25]),
    .Z(net114));
 BUF_X1 input115 (.A(int_polarity[26]),
    .Z(net115));
 BUF_X1 input116 (.A(int_polarity[27]),
    .Z(net116));
 BUF_X1 input117 (.A(int_polarity[28]),
    .Z(net117));
 BUF_X1 input118 (.A(int_polarity[29]),
    .Z(net118));
 BUF_X1 input119 (.A(int_polarity[2]),
    .Z(net119));
 BUF_X1 input120 (.A(int_polarity[30]),
    .Z(net120));
 BUF_X1 input121 (.A(int_polarity[31]),
    .Z(net121));
 BUF_X1 input122 (.A(int_polarity[3]),
    .Z(net122));
 BUF_X1 input123 (.A(int_polarity[4]),
    .Z(net123));
 BUF_X1 input124 (.A(int_polarity[5]),
    .Z(net124));
 BUF_X1 input125 (.A(int_polarity[6]),
    .Z(net125));
 BUF_X1 input126 (.A(int_polarity[7]),
    .Z(net126));
 BUF_X1 input127 (.A(int_polarity[8]),
    .Z(net127));
 BUF_X1 input128 (.A(int_polarity[9]),
    .Z(net128));
 BUF_X1 input129 (.A(int_type[0]),
    .Z(net129));
 BUF_X1 input130 (.A(int_type[10]),
    .Z(net130));
 BUF_X1 input131 (.A(int_type[11]),
    .Z(net131));
 BUF_X1 input132 (.A(int_type[12]),
    .Z(net132));
 BUF_X1 input133 (.A(int_type[13]),
    .Z(net133));
 BUF_X1 input134 (.A(int_type[14]),
    .Z(net134));
 BUF_X1 input135 (.A(int_type[15]),
    .Z(net135));
 BUF_X1 input136 (.A(int_type[16]),
    .Z(net136));
 BUF_X1 input137 (.A(int_type[17]),
    .Z(net137));
 BUF_X1 input138 (.A(int_type[18]),
    .Z(net138));
 BUF_X1 input139 (.A(int_type[19]),
    .Z(net139));
 BUF_X1 input140 (.A(int_type[1]),
    .Z(net140));
 BUF_X1 input141 (.A(int_type[20]),
    .Z(net141));
 BUF_X1 input142 (.A(int_type[21]),
    .Z(net142));
 BUF_X1 input143 (.A(int_type[22]),
    .Z(net143));
 BUF_X1 input144 (.A(int_type[23]),
    .Z(net144));
 BUF_X1 input145 (.A(int_type[24]),
    .Z(net145));
 BUF_X1 input146 (.A(int_type[25]),
    .Z(net146));
 BUF_X1 input147 (.A(int_type[26]),
    .Z(net147));
 BUF_X1 input148 (.A(int_type[27]),
    .Z(net148));
 BUF_X1 input149 (.A(int_type[28]),
    .Z(net149));
 BUF_X1 input150 (.A(int_type[29]),
    .Z(net150));
 BUF_X1 input151 (.A(int_type[2]),
    .Z(net151));
 BUF_X1 input152 (.A(int_type[30]),
    .Z(net152));
 BUF_X1 input153 (.A(int_type[31]),
    .Z(net153));
 BUF_X1 input154 (.A(int_type[3]),
    .Z(net154));
 BUF_X1 input155 (.A(int_type[4]),
    .Z(net155));
 BUF_X1 input156 (.A(int_type[5]),
    .Z(net156));
 BUF_X1 input157 (.A(int_type[6]),
    .Z(net157));
 BUF_X1 input158 (.A(int_type[7]),
    .Z(net158));
 BUF_X1 input159 (.A(int_type[8]),
    .Z(net159));
 BUF_X1 input160 (.A(int_type[9]),
    .Z(net160));
 BUF_X1 output161 (.A(net161),
    .Z(gpio_in[0]));
 BUF_X1 output162 (.A(net162),
    .Z(gpio_in[10]));
 BUF_X1 output163 (.A(net163),
    .Z(gpio_in[11]));
 BUF_X1 output164 (.A(net164),
    .Z(gpio_in[12]));
 BUF_X1 output165 (.A(net165),
    .Z(gpio_in[13]));
 BUF_X1 output166 (.A(net166),
    .Z(gpio_in[14]));
 BUF_X1 output167 (.A(net167),
    .Z(gpio_in[15]));
 BUF_X1 output168 (.A(net168),
    .Z(gpio_in[16]));
 BUF_X1 output169 (.A(net169),
    .Z(gpio_in[17]));
 BUF_X1 output170 (.A(net170),
    .Z(gpio_in[18]));
 BUF_X1 output171 (.A(net171),
    .Z(gpio_in[19]));
 BUF_X1 output172 (.A(net172),
    .Z(gpio_in[1]));
 BUF_X1 output173 (.A(net173),
    .Z(gpio_in[20]));
 BUF_X1 output174 (.A(net174),
    .Z(gpio_in[21]));
 BUF_X1 output175 (.A(net175),
    .Z(gpio_in[22]));
 BUF_X1 output176 (.A(net176),
    .Z(gpio_in[23]));
 BUF_X1 output177 (.A(net177),
    .Z(gpio_in[24]));
 BUF_X1 output178 (.A(net178),
    .Z(gpio_in[25]));
 BUF_X1 output179 (.A(net179),
    .Z(gpio_in[26]));
 BUF_X1 output180 (.A(net180),
    .Z(gpio_in[27]));
 BUF_X1 output181 (.A(net181),
    .Z(gpio_in[28]));
 BUF_X1 output182 (.A(net182),
    .Z(gpio_in[29]));
 BUF_X1 output183 (.A(net183),
    .Z(gpio_in[2]));
 BUF_X1 output184 (.A(net184),
    .Z(gpio_in[30]));
 BUF_X1 output185 (.A(net185),
    .Z(gpio_in[31]));
 BUF_X1 output186 (.A(net186),
    .Z(gpio_in[3]));
 BUF_X1 output187 (.A(net187),
    .Z(gpio_in[4]));
 BUF_X1 output188 (.A(net188),
    .Z(gpio_in[5]));
 BUF_X1 output189 (.A(net189),
    .Z(gpio_in[6]));
 BUF_X1 output190 (.A(net190),
    .Z(gpio_in[7]));
 BUF_X1 output191 (.A(net191),
    .Z(gpio_in[8]));
 BUF_X1 output192 (.A(net192),
    .Z(gpio_in[9]));
 BUF_X1 output193 (.A(net193),
    .Z(int_out));
 BUF_X1 output194 (.A(net194),
    .Z(int_status[0]));
 BUF_X1 output195 (.A(net195),
    .Z(int_status[10]));
 BUF_X1 output196 (.A(net196),
    .Z(int_status[11]));
 BUF_X1 output197 (.A(net197),
    .Z(int_status[12]));
 BUF_X1 output198 (.A(net198),
    .Z(int_status[13]));
 BUF_X1 output199 (.A(net199),
    .Z(int_status[14]));
 BUF_X1 output200 (.A(net200),
    .Z(int_status[15]));
 BUF_X1 output201 (.A(net201),
    .Z(int_status[16]));
 BUF_X1 output202 (.A(net202),
    .Z(int_status[17]));
 BUF_X1 output203 (.A(net203),
    .Z(int_status[18]));
 BUF_X1 output204 (.A(net204),
    .Z(int_status[19]));
 BUF_X1 output205 (.A(net205),
    .Z(int_status[1]));
 BUF_X1 output206 (.A(net206),
    .Z(int_status[20]));
 BUF_X1 output207 (.A(net207),
    .Z(int_status[21]));
 BUF_X1 output208 (.A(net208),
    .Z(int_status[22]));
 BUF_X1 output209 (.A(net209),
    .Z(int_status[23]));
 BUF_X1 output210 (.A(net210),
    .Z(int_status[24]));
 BUF_X1 output211 (.A(net211),
    .Z(int_status[25]));
 BUF_X1 output212 (.A(net212),
    .Z(int_status[26]));
 BUF_X1 output213 (.A(net213),
    .Z(int_status[27]));
 BUF_X1 output214 (.A(net214),
    .Z(int_status[28]));
 BUF_X1 output215 (.A(net215),
    .Z(int_status[29]));
 BUF_X1 output216 (.A(net216),
    .Z(int_status[2]));
 BUF_X1 output217 (.A(net217),
    .Z(int_status[30]));
 BUF_X1 output218 (.A(net218),
    .Z(int_status[31]));
 BUF_X1 output219 (.A(net219),
    .Z(int_status[3]));
 BUF_X1 output220 (.A(net220),
    .Z(int_status[4]));
 BUF_X1 output221 (.A(net221),
    .Z(int_status[5]));
 BUF_X1 output222 (.A(net222),
    .Z(int_status[6]));
 BUF_X1 output223 (.A(net223),
    .Z(int_status[7]));
 BUF_X1 output224 (.A(net224),
    .Z(int_status[8]));
 BUF_X1 output225 (.A(net225),
    .Z(int_status[9]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X2 clkload0 (.A(clknet_4_1_0_clk));
 INV_X2 clkload1 (.A(clknet_4_2_0_clk));
 INV_X2 clkload2 (.A(clknet_4_3_0_clk));
 INV_X2 clkload3 (.A(clknet_4_4_0_clk));
 CLKBUF_X1 clkload4 (.A(clknet_4_5_0_clk));
 INV_X2 clkload5 (.A(clknet_4_6_0_clk));
 INV_X1 clkload6 (.A(clknet_4_7_0_clk));
 INV_X2 clkload7 (.A(clknet_4_8_0_clk));
 INV_X4 clkload8 (.A(clknet_4_9_0_clk));
 CLKBUF_X1 clkload9 (.A(clknet_4_10_0_clk));
 INV_X2 clkload10 (.A(clknet_4_11_0_clk));
 INV_X2 clkload11 (.A(clknet_4_12_0_clk));
 INV_X2 clkload12 (.A(clknet_4_13_0_clk));
 INV_X2 clkload13 (.A(clknet_4_14_0_clk));
 CLKBUF_X1 clkload14 (.A(clknet_4_15_0_clk));
 FILLCELL_X2 FILLER_0_7 ();
 FILLCELL_X8 FILLER_0_15 ();
 FILLCELL_X4 FILLER_0_23 ();
 FILLCELL_X2 FILLER_0_27 ();
 FILLCELL_X1 FILLER_0_29 ();
 FILLCELL_X2 FILLER_0_107 ();
 FILLCELL_X2 FILLER_0_133 ();
 FILLCELL_X16 FILLER_0_200 ();
 FILLCELL_X4 FILLER_0_216 ();
 FILLCELL_X1 FILLER_0_220 ();
 FILLCELL_X1 FILLER_0_226 ();
 FILLCELL_X1 FILLER_0_231 ();
 FILLCELL_X8 FILLER_1_17 ();
 FILLCELL_X2 FILLER_1_29 ();
 FILLCELL_X1 FILLER_1_51 ();
 FILLCELL_X1 FILLER_1_60 ();
 FILLCELL_X2 FILLER_1_90 ();
 FILLCELL_X1 FILLER_1_98 ();
 FILLCELL_X4 FILLER_1_102 ();
 FILLCELL_X2 FILLER_1_106 ();
 FILLCELL_X1 FILLER_1_108 ();
 FILLCELL_X2 FILLER_1_117 ();
 FILLCELL_X2 FILLER_1_122 ();
 FILLCELL_X2 FILLER_1_129 ();
 FILLCELL_X1 FILLER_1_148 ();
 FILLCELL_X2 FILLER_1_153 ();
 FILLCELL_X1 FILLER_1_172 ();
 FILLCELL_X2 FILLER_1_183 ();
 FILLCELL_X4 FILLER_1_208 ();
 FILLCELL_X2 FILLER_1_212 ();
 FILLCELL_X1 FILLER_1_214 ();
 FILLCELL_X1 FILLER_2_1 ();
 FILLCELL_X1 FILLER_2_51 ();
 FILLCELL_X8 FILLER_2_58 ();
 FILLCELL_X4 FILLER_2_66 ();
 FILLCELL_X2 FILLER_2_70 ();
 FILLCELL_X1 FILLER_2_72 ();
 FILLCELL_X1 FILLER_2_76 ();
 FILLCELL_X2 FILLER_2_99 ();
 FILLCELL_X1 FILLER_2_101 ();
 FILLCELL_X1 FILLER_2_106 ();
 FILLCELL_X8 FILLER_2_128 ();
 FILLCELL_X2 FILLER_2_136 ();
 FILLCELL_X1 FILLER_2_138 ();
 FILLCELL_X1 FILLER_2_232 ();
 FILLCELL_X1 FILLER_2_237 ();
 FILLCELL_X1 FILLER_3_4 ();
 FILLCELL_X2 FILLER_3_8 ();
 FILLCELL_X1 FILLER_3_10 ();
 FILLCELL_X8 FILLER_3_15 ();
 FILLCELL_X4 FILLER_3_23 ();
 FILLCELL_X2 FILLER_3_27 ();
 FILLCELL_X2 FILLER_3_32 ();
 FILLCELL_X1 FILLER_3_34 ();
 FILLCELL_X2 FILLER_3_38 ();
 FILLCELL_X4 FILLER_3_63 ();
 FILLCELL_X1 FILLER_3_67 ();
 FILLCELL_X4 FILLER_3_73 ();
 FILLCELL_X2 FILLER_3_94 ();
 FILLCELL_X4 FILLER_3_120 ();
 FILLCELL_X8 FILLER_3_128 ();
 FILLCELL_X4 FILLER_3_136 ();
 FILLCELL_X1 FILLER_3_140 ();
 FILLCELL_X4 FILLER_3_145 ();
 FILLCELL_X2 FILLER_3_149 ();
 FILLCELL_X1 FILLER_3_151 ();
 FILLCELL_X2 FILLER_3_156 ();
 FILLCELL_X1 FILLER_3_158 ();
 FILLCELL_X2 FILLER_3_165 ();
 FILLCELL_X1 FILLER_3_167 ();
 FILLCELL_X16 FILLER_3_172 ();
 FILLCELL_X2 FILLER_3_188 ();
 FILLCELL_X1 FILLER_3_190 ();
 FILLCELL_X8 FILLER_3_202 ();
 FILLCELL_X2 FILLER_3_210 ();
 FILLCELL_X4 FILLER_4_4 ();
 FILLCELL_X4 FILLER_4_32 ();
 FILLCELL_X1 FILLER_4_36 ();
 FILLCELL_X8 FILLER_4_40 ();
 FILLCELL_X2 FILLER_4_48 ();
 FILLCELL_X4 FILLER_4_67 ();
 FILLCELL_X1 FILLER_4_71 ();
 FILLCELL_X16 FILLER_4_76 ();
 FILLCELL_X4 FILLER_4_92 ();
 FILLCELL_X1 FILLER_4_96 ();
 FILLCELL_X4 FILLER_4_101 ();
 FILLCELL_X2 FILLER_4_105 ();
 FILLCELL_X1 FILLER_4_107 ();
 FILLCELL_X2 FILLER_4_114 ();
 FILLCELL_X1 FILLER_4_116 ();
 FILLCELL_X1 FILLER_4_132 ();
 FILLCELL_X16 FILLER_4_137 ();
 FILLCELL_X2 FILLER_4_153 ();
 FILLCELL_X1 FILLER_4_155 ();
 FILLCELL_X2 FILLER_4_160 ();
 FILLCELL_X8 FILLER_4_181 ();
 FILLCELL_X2 FILLER_4_189 ();
 FILLCELL_X4 FILLER_4_212 ();
 FILLCELL_X1 FILLER_4_216 ();
 FILLCELL_X1 FILLER_5_1 ();
 FILLCELL_X1 FILLER_5_23 ();
 FILLCELL_X8 FILLER_5_45 ();
 FILLCELL_X2 FILLER_5_53 ();
 FILLCELL_X8 FILLER_5_59 ();
 FILLCELL_X32 FILLER_5_84 ();
 FILLCELL_X4 FILLER_5_116 ();
 FILLCELL_X2 FILLER_5_120 ();
 FILLCELL_X2 FILLER_5_126 ();
 FILLCELL_X4 FILLER_5_138 ();
 FILLCELL_X8 FILLER_5_144 ();
 FILLCELL_X1 FILLER_5_152 ();
 FILLCELL_X8 FILLER_5_170 ();
 FILLCELL_X2 FILLER_5_178 ();
 FILLCELL_X8 FILLER_5_184 ();
 FILLCELL_X4 FILLER_5_192 ();
 FILLCELL_X2 FILLER_5_196 ();
 FILLCELL_X1 FILLER_5_198 ();
 FILLCELL_X4 FILLER_5_202 ();
 FILLCELL_X1 FILLER_5_206 ();
 FILLCELL_X1 FILLER_5_234 ();
 FILLCELL_X8 FILLER_6_23 ();
 FILLCELL_X4 FILLER_6_31 ();
 FILLCELL_X2 FILLER_6_52 ();
 FILLCELL_X16 FILLER_6_75 ();
 FILLCELL_X4 FILLER_6_91 ();
 FILLCELL_X2 FILLER_6_95 ();
 FILLCELL_X4 FILLER_6_114 ();
 FILLCELL_X8 FILLER_6_152 ();
 FILLCELL_X8 FILLER_6_165 ();
 FILLCELL_X2 FILLER_6_173 ();
 FILLCELL_X4 FILLER_6_201 ();
 FILLCELL_X1 FILLER_6_205 ();
 FILLCELL_X1 FILLER_6_219 ();
 FILLCELL_X1 FILLER_6_224 ();
 FILLCELL_X1 FILLER_6_234 ();
 FILLCELL_X1 FILLER_7_16 ();
 FILLCELL_X4 FILLER_7_24 ();
 FILLCELL_X2 FILLER_7_28 ();
 FILLCELL_X1 FILLER_7_30 ();
 FILLCELL_X8 FILLER_7_48 ();
 FILLCELL_X4 FILLER_7_56 ();
 FILLCELL_X4 FILLER_7_65 ();
 FILLCELL_X2 FILLER_7_69 ();
 FILLCELL_X2 FILLER_7_110 ();
 FILLCELL_X4 FILLER_7_129 ();
 FILLCELL_X1 FILLER_7_133 ();
 FILLCELL_X4 FILLER_7_139 ();
 FILLCELL_X1 FILLER_7_143 ();
 FILLCELL_X2 FILLER_7_156 ();
 FILLCELL_X2 FILLER_7_179 ();
 FILLCELL_X1 FILLER_7_190 ();
 FILLCELL_X8 FILLER_7_195 ();
 FILLCELL_X1 FILLER_7_234 ();
 FILLCELL_X4 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_9 ();
 FILLCELL_X1 FILLER_8_14 ();
 FILLCELL_X4 FILLER_8_36 ();
 FILLCELL_X1 FILLER_8_40 ();
 FILLCELL_X1 FILLER_8_45 ();
 FILLCELL_X16 FILLER_8_69 ();
 FILLCELL_X2 FILLER_8_85 ();
 FILLCELL_X4 FILLER_8_91 ();
 FILLCELL_X2 FILLER_8_95 ();
 FILLCELL_X4 FILLER_8_104 ();
 FILLCELL_X32 FILLER_8_112 ();
 FILLCELL_X16 FILLER_8_144 ();
 FILLCELL_X1 FILLER_8_160 ();
 FILLCELL_X1 FILLER_8_180 ();
 FILLCELL_X8 FILLER_8_201 ();
 FILLCELL_X4 FILLER_8_209 ();
 FILLCELL_X2 FILLER_8_213 ();
 FILLCELL_X1 FILLER_8_215 ();
 FILLCELL_X1 FILLER_8_219 ();
 FILLCELL_X2 FILLER_8_224 ();
 FILLCELL_X1 FILLER_8_231 ();
 FILLCELL_X1 FILLER_9_11 ();
 FILLCELL_X2 FILLER_9_35 ();
 FILLCELL_X1 FILLER_9_37 ();
 FILLCELL_X32 FILLER_9_59 ();
 FILLCELL_X8 FILLER_9_91 ();
 FILLCELL_X4 FILLER_9_99 ();
 FILLCELL_X2 FILLER_9_120 ();
 FILLCELL_X1 FILLER_9_143 ();
 FILLCELL_X4 FILLER_9_148 ();
 FILLCELL_X1 FILLER_9_152 ();
 FILLCELL_X2 FILLER_9_160 ();
 FILLCELL_X8 FILLER_9_170 ();
 FILLCELL_X4 FILLER_9_178 ();
 FILLCELL_X1 FILLER_9_182 ();
 FILLCELL_X16 FILLER_9_187 ();
 FILLCELL_X4 FILLER_9_203 ();
 FILLCELL_X2 FILLER_9_210 ();
 FILLCELL_X1 FILLER_9_212 ();
 FILLCELL_X1 FILLER_9_237 ();
 FILLCELL_X1 FILLER_10_20 ();
 FILLCELL_X16 FILLER_10_28 ();
 FILLCELL_X4 FILLER_10_44 ();
 FILLCELL_X32 FILLER_10_56 ();
 FILLCELL_X32 FILLER_10_88 ();
 FILLCELL_X8 FILLER_10_120 ();
 FILLCELL_X4 FILLER_10_128 ();
 FILLCELL_X2 FILLER_10_132 ();
 FILLCELL_X1 FILLER_10_134 ();
 FILLCELL_X2 FILLER_10_139 ();
 FILLCELL_X1 FILLER_10_141 ();
 FILLCELL_X8 FILLER_10_169 ();
 FILLCELL_X2 FILLER_10_177 ();
 FILLCELL_X8 FILLER_10_200 ();
 FILLCELL_X1 FILLER_10_208 ();
 FILLCELL_X4 FILLER_10_213 ();
 FILLCELL_X2 FILLER_11_7 ();
 FILLCELL_X4 FILLER_11_23 ();
 FILLCELL_X32 FILLER_11_64 ();
 FILLCELL_X32 FILLER_11_96 ();
 FILLCELL_X4 FILLER_11_128 ();
 FILLCELL_X2 FILLER_11_132 ();
 FILLCELL_X1 FILLER_11_134 ();
 FILLCELL_X2 FILLER_11_152 ();
 FILLCELL_X16 FILLER_11_162 ();
 FILLCELL_X4 FILLER_11_178 ();
 FILLCELL_X2 FILLER_11_182 ();
 FILLCELL_X1 FILLER_11_184 ();
 FILLCELL_X1 FILLER_12_10 ();
 FILLCELL_X2 FILLER_12_41 ();
 FILLCELL_X1 FILLER_12_43 ();
 FILLCELL_X32 FILLER_12_57 ();
 FILLCELL_X32 FILLER_12_89 ();
 FILLCELL_X16 FILLER_12_121 ();
 FILLCELL_X8 FILLER_12_137 ();
 FILLCELL_X4 FILLER_12_145 ();
 FILLCELL_X2 FILLER_12_149 ();
 FILLCELL_X1 FILLER_12_151 ();
 FILLCELL_X4 FILLER_12_156 ();
 FILLCELL_X1 FILLER_12_181 ();
 FILLCELL_X32 FILLER_12_186 ();
 FILLCELL_X2 FILLER_12_227 ();
 FILLCELL_X1 FILLER_12_231 ();
 FILLCELL_X2 FILLER_13_4 ();
 FILLCELL_X1 FILLER_13_6 ();
 FILLCELL_X8 FILLER_13_22 ();
 FILLCELL_X2 FILLER_13_30 ();
 FILLCELL_X1 FILLER_13_32 ();
 FILLCELL_X4 FILLER_13_67 ();
 FILLCELL_X32 FILLER_13_75 ();
 FILLCELL_X32 FILLER_13_107 ();
 FILLCELL_X8 FILLER_13_139 ();
 FILLCELL_X4 FILLER_13_147 ();
 FILLCELL_X2 FILLER_13_151 ();
 FILLCELL_X1 FILLER_13_153 ();
 FILLCELL_X2 FILLER_13_171 ();
 FILLCELL_X1 FILLER_13_173 ();
 FILLCELL_X8 FILLER_13_199 ();
 FILLCELL_X4 FILLER_13_211 ();
 FILLCELL_X2 FILLER_13_215 ();
 FILLCELL_X1 FILLER_13_217 ();
 FILLCELL_X1 FILLER_13_227 ();
 FILLCELL_X1 FILLER_13_234 ();
 FILLCELL_X2 FILLER_14_15 ();
 FILLCELL_X8 FILLER_14_34 ();
 FILLCELL_X1 FILLER_14_42 ();
 FILLCELL_X16 FILLER_14_47 ();
 FILLCELL_X8 FILLER_14_63 ();
 FILLCELL_X4 FILLER_14_88 ();
 FILLCELL_X2 FILLER_14_92 ();
 FILLCELL_X1 FILLER_14_94 ();
 FILLCELL_X16 FILLER_14_99 ();
 FILLCELL_X4 FILLER_14_115 ();
 FILLCELL_X2 FILLER_14_119 ();
 FILLCELL_X8 FILLER_14_125 ();
 FILLCELL_X1 FILLER_14_137 ();
 FILLCELL_X4 FILLER_14_142 ();
 FILLCELL_X2 FILLER_14_146 ();
 FILLCELL_X16 FILLER_14_152 ();
 FILLCELL_X8 FILLER_14_168 ();
 FILLCELL_X8 FILLER_14_180 ();
 FILLCELL_X2 FILLER_14_188 ();
 FILLCELL_X1 FILLER_14_190 ();
 FILLCELL_X1 FILLER_14_225 ();
 FILLCELL_X2 FILLER_14_236 ();
 FILLCELL_X1 FILLER_15_7 ();
 FILLCELL_X1 FILLER_15_11 ();
 FILLCELL_X2 FILLER_15_40 ();
 FILLCELL_X32 FILLER_15_59 ();
 FILLCELL_X32 FILLER_15_91 ();
 FILLCELL_X8 FILLER_15_123 ();
 FILLCELL_X4 FILLER_15_131 ();
 FILLCELL_X1 FILLER_15_135 ();
 FILLCELL_X8 FILLER_15_159 ();
 FILLCELL_X4 FILLER_15_167 ();
 FILLCELL_X2 FILLER_15_171 ();
 FILLCELL_X1 FILLER_15_173 ();
 FILLCELL_X16 FILLER_15_195 ();
 FILLCELL_X1 FILLER_15_237 ();
 FILLCELL_X2 FILLER_16_4 ();
 FILLCELL_X2 FILLER_16_23 ();
 FILLCELL_X1 FILLER_16_29 ();
 FILLCELL_X16 FILLER_16_47 ();
 FILLCELL_X4 FILLER_16_63 ();
 FILLCELL_X2 FILLER_16_67 ();
 FILLCELL_X2 FILLER_16_76 ();
 FILLCELL_X32 FILLER_16_84 ();
 FILLCELL_X4 FILLER_16_116 ();
 FILLCELL_X2 FILLER_16_120 ();
 FILLCELL_X1 FILLER_16_122 ();
 FILLCELL_X4 FILLER_16_128 ();
 FILLCELL_X1 FILLER_16_132 ();
 FILLCELL_X4 FILLER_16_137 ();
 FILLCELL_X1 FILLER_16_141 ();
 FILLCELL_X16 FILLER_16_145 ();
 FILLCELL_X8 FILLER_16_161 ();
 FILLCELL_X2 FILLER_16_169 ();
 FILLCELL_X16 FILLER_16_195 ();
 FILLCELL_X8 FILLER_16_211 ();
 FILLCELL_X1 FILLER_16_234 ();
 FILLCELL_X32 FILLER_17_29 ();
 FILLCELL_X32 FILLER_17_61 ();
 FILLCELL_X16 FILLER_17_93 ();
 FILLCELL_X8 FILLER_17_109 ();
 FILLCELL_X4 FILLER_17_117 ();
 FILLCELL_X2 FILLER_17_121 ();
 FILLCELL_X16 FILLER_17_127 ();
 FILLCELL_X8 FILLER_17_143 ();
 FILLCELL_X1 FILLER_17_151 ();
 FILLCELL_X16 FILLER_17_156 ();
 FILLCELL_X8 FILLER_17_172 ();
 FILLCELL_X4 FILLER_17_180 ();
 FILLCELL_X2 FILLER_17_184 ();
 FILLCELL_X1 FILLER_17_203 ();
 FILLCELL_X4 FILLER_17_213 ();
 FILLCELL_X1 FILLER_17_217 ();
 FILLCELL_X2 FILLER_17_231 ();
 FILLCELL_X2 FILLER_17_236 ();
 FILLCELL_X1 FILLER_18_12 ();
 FILLCELL_X16 FILLER_18_30 ();
 FILLCELL_X4 FILLER_18_46 ();
 FILLCELL_X2 FILLER_18_50 ();
 FILLCELL_X1 FILLER_18_52 ();
 FILLCELL_X8 FILLER_18_67 ();
 FILLCELL_X4 FILLER_18_75 ();
 FILLCELL_X1 FILLER_18_79 ();
 FILLCELL_X32 FILLER_18_88 ();
 FILLCELL_X32 FILLER_18_120 ();
 FILLCELL_X32 FILLER_18_152 ();
 FILLCELL_X16 FILLER_18_184 ();
 FILLCELL_X8 FILLER_18_200 ();
 FILLCELL_X1 FILLER_18_237 ();
 FILLCELL_X2 FILLER_19_10 ();
 FILLCELL_X2 FILLER_19_19 ();
 FILLCELL_X4 FILLER_19_25 ();
 FILLCELL_X2 FILLER_19_29 ();
 FILLCELL_X1 FILLER_19_31 ();
 FILLCELL_X1 FILLER_19_53 ();
 FILLCELL_X1 FILLER_19_57 ();
 FILLCELL_X32 FILLER_19_79 ();
 FILLCELL_X16 FILLER_19_111 ();
 FILLCELL_X8 FILLER_19_127 ();
 FILLCELL_X4 FILLER_19_135 ();
 FILLCELL_X8 FILLER_19_143 ();
 FILLCELL_X4 FILLER_19_151 ();
 FILLCELL_X1 FILLER_19_155 ();
 FILLCELL_X2 FILLER_19_180 ();
 FILLCELL_X1 FILLER_19_182 ();
 FILLCELL_X4 FILLER_19_187 ();
 FILLCELL_X1 FILLER_19_191 ();
 FILLCELL_X4 FILLER_19_200 ();
 FILLCELL_X2 FILLER_19_204 ();
 FILLCELL_X1 FILLER_19_237 ();
 FILLCELL_X2 FILLER_20_36 ();
 FILLCELL_X32 FILLER_20_59 ();
 FILLCELL_X32 FILLER_20_91 ();
 FILLCELL_X4 FILLER_20_123 ();
 FILLCELL_X8 FILLER_20_131 ();
 FILLCELL_X4 FILLER_20_139 ();
 FILLCELL_X2 FILLER_20_143 ();
 FILLCELL_X1 FILLER_20_145 ();
 FILLCELL_X2 FILLER_20_167 ();
 FILLCELL_X4 FILLER_20_173 ();
 FILLCELL_X4 FILLER_20_181 ();
 FILLCELL_X2 FILLER_20_185 ();
 FILLCELL_X1 FILLER_20_187 ();
 FILLCELL_X4 FILLER_20_217 ();
 FILLCELL_X1 FILLER_21_10 ();
 FILLCELL_X1 FILLER_21_18 ();
 FILLCELL_X8 FILLER_21_22 ();
 FILLCELL_X1 FILLER_21_34 ();
 FILLCELL_X1 FILLER_21_38 ();
 FILLCELL_X16 FILLER_21_59 ();
 FILLCELL_X4 FILLER_21_75 ();
 FILLCELL_X2 FILLER_21_79 ();
 FILLCELL_X2 FILLER_21_95 ();
 FILLCELL_X1 FILLER_21_97 ();
 FILLCELL_X4 FILLER_21_115 ();
 FILLCELL_X16 FILLER_21_123 ();
 FILLCELL_X8 FILLER_21_139 ();
 FILLCELL_X4 FILLER_21_147 ();
 FILLCELL_X2 FILLER_21_151 ();
 FILLCELL_X1 FILLER_21_153 ();
 FILLCELL_X4 FILLER_21_217 ();
 FILLCELL_X1 FILLER_21_221 ();
 FILLCELL_X4 FILLER_21_224 ();
 FILLCELL_X1 FILLER_21_228 ();
 FILLCELL_X8 FILLER_22_10 ();
 FILLCELL_X1 FILLER_22_18 ();
 FILLCELL_X8 FILLER_22_22 ();
 FILLCELL_X2 FILLER_22_30 ();
 FILLCELL_X8 FILLER_22_36 ();
 FILLCELL_X4 FILLER_22_44 ();
 FILLCELL_X2 FILLER_22_53 ();
 FILLCELL_X1 FILLER_22_55 ();
 FILLCELL_X4 FILLER_22_60 ();
 FILLCELL_X2 FILLER_22_64 ();
 FILLCELL_X1 FILLER_22_66 ();
 FILLCELL_X4 FILLER_22_105 ();
 FILLCELL_X2 FILLER_22_109 ();
 FILLCELL_X4 FILLER_22_115 ();
 FILLCELL_X4 FILLER_22_142 ();
 FILLCELL_X2 FILLER_22_146 ();
 FILLCELL_X1 FILLER_22_148 ();
 FILLCELL_X16 FILLER_22_153 ();
 FILLCELL_X8 FILLER_22_169 ();
 FILLCELL_X2 FILLER_22_177 ();
 FILLCELL_X4 FILLER_22_183 ();
 FILLCELL_X1 FILLER_22_187 ();
 FILLCELL_X1 FILLER_22_210 ();
 FILLCELL_X2 FILLER_22_214 ();
 FILLCELL_X1 FILLER_22_219 ();
 FILLCELL_X1 FILLER_22_224 ();
 FILLCELL_X2 FILLER_23_7 ();
 FILLCELL_X8 FILLER_23_51 ();
 FILLCELL_X4 FILLER_23_59 ();
 FILLCELL_X2 FILLER_23_63 ();
 FILLCELL_X8 FILLER_23_69 ();
 FILLCELL_X4 FILLER_23_77 ();
 FILLCELL_X2 FILLER_23_81 ();
 FILLCELL_X1 FILLER_23_83 ();
 FILLCELL_X8 FILLER_23_88 ();
 FILLCELL_X4 FILLER_23_96 ();
 FILLCELL_X16 FILLER_23_117 ();
 FILLCELL_X8 FILLER_23_167 ();
 FILLCELL_X2 FILLER_23_175 ();
 FILLCELL_X4 FILLER_23_194 ();
 FILLCELL_X2 FILLER_23_198 ();
 FILLCELL_X2 FILLER_23_207 ();
 FILLCELL_X1 FILLER_23_209 ();
 FILLCELL_X1 FILLER_23_215 ();
 FILLCELL_X1 FILLER_24_10 ();
 FILLCELL_X8 FILLER_24_32 ();
 FILLCELL_X4 FILLER_24_40 ();
 FILLCELL_X8 FILLER_24_82 ();
 FILLCELL_X4 FILLER_24_90 ();
 FILLCELL_X2 FILLER_24_94 ();
 FILLCELL_X8 FILLER_24_134 ();
 FILLCELL_X4 FILLER_24_142 ();
 FILLCELL_X2 FILLER_24_146 ();
 FILLCELL_X4 FILLER_24_152 ();
 FILLCELL_X1 FILLER_24_156 ();
 FILLCELL_X4 FILLER_24_178 ();
 FILLCELL_X4 FILLER_24_187 ();
 FILLCELL_X2 FILLER_24_191 ();
 FILLCELL_X8 FILLER_24_203 ();
 FILLCELL_X2 FILLER_24_211 ();
 FILLCELL_X1 FILLER_25_21 ();
 FILLCELL_X4 FILLER_25_25 ();
 FILLCELL_X2 FILLER_25_29 ();
 FILLCELL_X1 FILLER_25_31 ();
 FILLCELL_X2 FILLER_25_49 ();
 FILLCELL_X1 FILLER_25_51 ();
 FILLCELL_X4 FILLER_25_56 ();
 FILLCELL_X4 FILLER_25_68 ();
 FILLCELL_X2 FILLER_25_72 ();
 FILLCELL_X4 FILLER_25_91 ();
 FILLCELL_X2 FILLER_25_95 ();
 FILLCELL_X16 FILLER_25_105 ();
 FILLCELL_X1 FILLER_25_138 ();
 FILLCELL_X2 FILLER_25_143 ();
 FILLCELL_X1 FILLER_25_157 ();
 FILLCELL_X4 FILLER_25_162 ();
 FILLCELL_X2 FILLER_25_166 ();
 FILLCELL_X1 FILLER_25_168 ();
 FILLCELL_X4 FILLER_25_173 ();
 FILLCELL_X2 FILLER_25_194 ();
 FILLCELL_X8 FILLER_25_204 ();
 FILLCELL_X4 FILLER_25_212 ();
 FILLCELL_X1 FILLER_25_216 ();
 FILLCELL_X2 FILLER_25_228 ();
 FILLCELL_X1 FILLER_25_230 ();
 FILLCELL_X1 FILLER_25_234 ();
 FILLCELL_X1 FILLER_26_4 ();
 FILLCELL_X1 FILLER_26_8 ();
 FILLCELL_X1 FILLER_26_12 ();
 FILLCELL_X8 FILLER_26_38 ();
 FILLCELL_X4 FILLER_26_46 ();
 FILLCELL_X2 FILLER_26_50 ();
 FILLCELL_X1 FILLER_26_52 ();
 FILLCELL_X8 FILLER_26_70 ();
 FILLCELL_X4 FILLER_26_91 ();
 FILLCELL_X2 FILLER_26_95 ();
 FILLCELL_X1 FILLER_26_97 ();
 FILLCELL_X2 FILLER_26_102 ();
 FILLCELL_X1 FILLER_26_104 ();
 FILLCELL_X8 FILLER_26_109 ();
 FILLCELL_X2 FILLER_26_117 ();
 FILLCELL_X1 FILLER_26_119 ();
 FILLCELL_X4 FILLER_26_124 ();
 FILLCELL_X2 FILLER_26_128 ();
 FILLCELL_X1 FILLER_26_147 ();
 FILLCELL_X8 FILLER_26_185 ();
 FILLCELL_X4 FILLER_26_193 ();
 FILLCELL_X1 FILLER_26_216 ();
 FILLCELL_X2 FILLER_27_10 ();
 FILLCELL_X2 FILLER_27_29 ();
 FILLCELL_X1 FILLER_27_31 ();
 FILLCELL_X2 FILLER_27_36 ();
 FILLCELL_X1 FILLER_27_38 ();
 FILLCELL_X32 FILLER_27_43 ();
 FILLCELL_X8 FILLER_27_75 ();
 FILLCELL_X2 FILLER_27_83 ();
 FILLCELL_X8 FILLER_27_93 ();
 FILLCELL_X2 FILLER_27_101 ();
 FILLCELL_X16 FILLER_27_120 ();
 FILLCELL_X4 FILLER_27_136 ();
 FILLCELL_X16 FILLER_27_145 ();
 FILLCELL_X4 FILLER_27_161 ();
 FILLCELL_X16 FILLER_27_169 ();
 FILLCELL_X4 FILLER_27_185 ();
 FILLCELL_X2 FILLER_27_189 ();
 FILLCELL_X4 FILLER_27_201 ();
 FILLCELL_X1 FILLER_27_205 ();
 FILLCELL_X2 FILLER_27_209 ();
 FILLCELL_X4 FILLER_28_17 ();
 FILLCELL_X1 FILLER_28_21 ();
 FILLCELL_X1 FILLER_28_60 ();
 FILLCELL_X1 FILLER_28_64 ();
 FILLCELL_X16 FILLER_28_67 ();
 FILLCELL_X2 FILLER_28_83 ();
 FILLCELL_X1 FILLER_28_85 ();
 FILLCELL_X16 FILLER_28_90 ();
 FILLCELL_X2 FILLER_28_106 ();
 FILLCELL_X1 FILLER_28_108 ();
 FILLCELL_X1 FILLER_28_116 ();
 FILLCELL_X16 FILLER_28_123 ();
 FILLCELL_X4 FILLER_28_139 ();
 FILLCELL_X8 FILLER_28_150 ();
 FILLCELL_X4 FILLER_28_158 ();
 FILLCELL_X1 FILLER_28_162 ();
 FILLCELL_X8 FILLER_28_180 ();
 FILLCELL_X2 FILLER_28_188 ();
 FILLCELL_X1 FILLER_28_190 ();
 FILLCELL_X8 FILLER_28_208 ();
 FILLCELL_X1 FILLER_28_216 ();
 FILLCELL_X4 FILLER_28_234 ();
 FILLCELL_X2 FILLER_29_10 ();
 FILLCELL_X16 FILLER_29_15 ();
 FILLCELL_X1 FILLER_29_35 ();
 FILLCELL_X2 FILLER_29_45 ();
 FILLCELL_X1 FILLER_29_54 ();
 FILLCELL_X2 FILLER_29_84 ();
 FILLCELL_X1 FILLER_29_86 ();
 FILLCELL_X2 FILLER_29_108 ();
 FILLCELL_X1 FILLER_29_110 ();
 FILLCELL_X2 FILLER_29_150 ();
 FILLCELL_X2 FILLER_29_161 ();
 FILLCELL_X4 FILLER_29_187 ();
 FILLCELL_X2 FILLER_29_191 ();
 FILLCELL_X4 FILLER_29_199 ();
 FILLCELL_X2 FILLER_29_206 ();
 FILLCELL_X2 FILLER_29_233 ();
 FILLCELL_X16 FILLER_30_1 ();
 FILLCELL_X4 FILLER_30_17 ();
 FILLCELL_X1 FILLER_30_21 ();
 FILLCELL_X2 FILLER_30_42 ();
 FILLCELL_X2 FILLER_30_54 ();
 FILLCELL_X1 FILLER_30_100 ();
 FILLCELL_X1 FILLER_30_128 ();
 FILLCELL_X1 FILLER_30_138 ();
 FILLCELL_X2 FILLER_30_209 ();
 FILLCELL_X4 FILLER_30_232 ();
 FILLCELL_X2 FILLER_30_236 ();
 FILLCELL_X16 FILLER_31_1 ();
 FILLCELL_X8 FILLER_31_17 ();
 FILLCELL_X1 FILLER_31_130 ();
 FILLCELL_X1 FILLER_31_210 ();
 FILLCELL_X16 FILLER_31_218 ();
 FILLCELL_X4 FILLER_31_234 ();
endmodule
