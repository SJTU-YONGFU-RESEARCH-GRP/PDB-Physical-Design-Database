module loadable_updown_counter (clk,
    enable,
    load_en,
    overflow,
    rst_n,
    underflow,
    up_down,
    count,
    load_val);
 input clk;
 input enable;
 input load_en;
 output overflow;
 input rst_n;
 output underflow;
 input up_down;
 output [7:0] count;
 input [7:0] load_val;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net23;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _091_ (.I(net13),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _092_ (.I(net14),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _093_ (.I(net12),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _094_ (.I0(_074_),
    .I1(net4),
    .S(net3),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _095_ (.I(net2),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _096_ (.I0(net13),
    .I1(_030_),
    .S(_031_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _097_ (.I(_077_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _098_ (.I(net3),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _099_ (.I0(net5),
    .I1(_032_),
    .S(_033_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _100_ (.I0(net14),
    .I1(_034_),
    .S(_031_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _101_ (.A1(_082_),
    .A2(_076_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _102_ (.I0(net6),
    .I1(_035_),
    .S(_033_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _103_ (.I0(net15),
    .I1(_036_),
    .S(_031_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _104_ (.I(_031_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _105_ (.I(net7),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _106_ (.A1(net13),
    .A2(_082_),
    .A3(_080_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _107_ (.A1(_082_),
    .A2(_079_),
    .B(_081_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _108_ (.A1(_039_),
    .A2(_040_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _109_ (.A1(_086_),
    .A2(_041_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _110_ (.I0(_038_),
    .I1(_042_),
    .S(_033_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _111_ (.A1(_037_),
    .A2(net16),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _112_ (.A1(_037_),
    .A2(_043_),
    .B(_044_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _113_ (.I(_082_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _114_ (.I(_081_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _115_ (.A1(_045_),
    .A2(_076_),
    .B(_046_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _116_ (.A1(_086_),
    .A2(_047_),
    .B(_085_),
    .C(_084_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _117_ (.I(_085_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _118_ (.A1(_045_),
    .A2(_076_),
    .B(_046_),
    .C(_049_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _119_ (.A1(_086_),
    .A2(_085_),
    .B(_084_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _120_ (.I(_051_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _121_ (.A1(_050_),
    .A2(_052_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _122_ (.A1(net3),
    .A2(net8),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _123_ (.A1(net3),
    .A2(_048_),
    .A3(_053_),
    .B(_054_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _124_ (.I0(net17),
    .I1(_055_),
    .S(_031_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _125_ (.A1(_086_),
    .A2(_084_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _126_ (.A1(_084_),
    .A2(_085_),
    .B(_083_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _127_ (.A1(_041_),
    .A2(_056_),
    .B(_057_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _128_ (.A1(_088_),
    .A2(_058_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _129_ (.A1(_033_),
    .A2(_031_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _130_ (.A1(net3),
    .A2(_031_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _131_ (.A1(_037_),
    .A2(net18),
    .B1(net9),
    .B2(_061_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _132_ (.A1(_059_),
    .A2(_060_),
    .B(_062_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _133_ (.I(_076_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _134_ (.A1(_082_),
    .A2(_063_),
    .B(_081_),
    .C(_085_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _135_ (.I(_083_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _136_ (.A1(_064_),
    .A2(_051_),
    .B(_065_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _137_ (.A1(_088_),
    .A2(_066_),
    .B(_087_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _138_ (.A1(_090_),
    .A2(_060_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _139_ (.I(_088_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _140_ (.A1(_050_),
    .A2(_052_),
    .B(_083_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _141_ (.A1(_033_),
    .A2(_031_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _142_ (.A1(_090_),
    .A2(_071_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _143_ (.I(_087_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _144_ (.A1(_069_),
    .A2(_070_),
    .B(_072_),
    .C(_073_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _145_ (.A1(_037_),
    .A2(net19),
    .B1(net10),
    .B2(_061_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _146_ (.A1(_067_),
    .A2(_068_),
    .B(_008_),
    .C(_009_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _147_ (.A1(_088_),
    .A2(_090_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _148_ (.A1(_039_),
    .A2(_040_),
    .B(_056_),
    .C(_010_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _149_ (.A1(_090_),
    .A2(_087_),
    .B(_089_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _150_ (.A1(_057_),
    .A2(_010_),
    .B(_012_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _151_ (.A1(_033_),
    .A2(_031_),
    .A3(net20),
    .A4(net12),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _152_ (.A1(_011_),
    .A2(_013_),
    .B(_014_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _153_ (.A1(net2),
    .A2(net20),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _154_ (.A1(_033_),
    .A2(_078_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _155_ (.A1(_011_),
    .A2(_013_),
    .A3(_016_),
    .A4(_017_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _156_ (.A1(net3),
    .A2(net20),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _157_ (.A1(_011_),
    .A2(_013_),
    .B(_019_),
    .C(_078_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _158_ (.A1(net3),
    .A2(net20),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _159_ (.A1(_078_),
    .A2(_011_),
    .A3(_013_),
    .A4(_021_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _160_ (.A1(_015_),
    .A2(_018_),
    .A3(_020_),
    .A4(_022_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _161_ (.A1(_033_),
    .A2(_037_),
    .A3(net11),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _162_ (.A1(_031_),
    .A2(net20),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _163_ (.A1(_023_),
    .A2(_024_),
    .A3(_025_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _164_ (.A1(net18),
    .A2(net17),
    .A3(net19),
    .A4(net20),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _165_ (.A1(net14),
    .A2(net12),
    .A3(_071_),
    .A4(_026_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _166_ (.A1(net13),
    .A2(net16),
    .A3(net15),
    .A4(_027_),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _167_ (.A1(net18),
    .A2(net17),
    .A3(net19),
    .A4(net20),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _168_ (.A1(net14),
    .A2(net12),
    .A3(_060_),
    .A4(_028_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _169_ (.A1(net13),
    .A2(net16),
    .A3(net15),
    .A4(_029_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _170_ (.A(_074_),
    .B(_075_),
    .CI(net12),
    .CO(_076_),
    .S(_077_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _171_ (.A(net14),
    .B(_078_),
    .CO(_079_),
    .S(_080_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _172_ (.A(net15),
    .B(_078_),
    .CO(_081_),
    .S(_082_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _173_ (.A(net17),
    .B(_078_),
    .CO(_083_),
    .S(_084_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _174_ (.A(net16),
    .B(_078_),
    .CO(_085_),
    .S(_086_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _175_ (.A(net18),
    .B(_078_),
    .CO(_087_),
    .S(_088_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _176_ (.A(net19),
    .B(_078_),
    .CO(_089_),
    .S(_090_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[1]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[2]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[3]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[4]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[5]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[6]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[7]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 hold1 (.I(net23),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_78 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_79 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_80 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_81 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_82 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_83 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_84 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_85 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_86 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_87 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_88 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_89 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_90 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_91 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_92 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_93 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_94 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_95 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_96 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_97 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_98 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_99 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_118 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input2 (.I(load_en),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(load_val[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(load_val[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(load_val[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(load_val[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(load_val[4]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(load_val[5]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(load_val[6]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(load_val[7]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input11 (.I(up_down),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(count[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(count[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(count[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(overflow));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(underflow));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_358 ();
endmodule
