module universal_shift_register (clk,
    enable,
    load,
    rst_n,
    serial_in_left,
    serial_in_right,
    direction,
    parallel_in,
    parallel_out);
 input clk;
 input enable;
 input load;
 input rst_n;
 input serial_in_left;
 input serial_in_right;
 input [1:0] direction;
 input [7:0] parallel_in;
 output [7:0] parallel_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire \shift_right_count[0] ;
 wire \shift_right_count[1] ;
 wire \shift_right_count[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X2 _126_ (.A(net11),
    .ZN(_066_));
 BUF_X2 _127_ (.A(enable),
    .Z(_067_));
 INV_X2 _128_ (.A(_067_),
    .ZN(_068_));
 AND2_X1 _129_ (.A1(_067_),
    .A2(_113_),
    .ZN(_069_));
 INV_X2 _130_ (.A(_114_),
    .ZN(_070_));
 NAND2_X2 _131_ (.A1(_110_),
    .A2(_070_),
    .ZN(_071_));
 MUX2_X1 _132_ (.A(_069_),
    .B(\shift_right_count[1] ),
    .S(_071_),
    .Z(_072_));
 BUF_X2 _133_ (.A(load),
    .Z(_073_));
 INV_X1 _134_ (.A(_073_),
    .ZN(_074_));
 BUF_X4 _135_ (.A(_074_),
    .Z(_075_));
 AOI22_X4 _136_ (.A1(_068_),
    .A2(\shift_right_count[1] ),
    .B1(_072_),
    .B2(_075_),
    .ZN(_076_));
 NOR2_X1 _137_ (.A1(_066_),
    .A2(_076_),
    .ZN(_123_));
 NOR2_X1 _138_ (.A1(_067_),
    .A2(_014_),
    .ZN(_077_));
 NOR2_X1 _139_ (.A1(_073_),
    .A2(_014_),
    .ZN(_078_));
 INV_X1 _140_ (.A(_110_),
    .ZN(_079_));
 NOR4_X2 _141_ (.A1(_079_),
    .A2(_068_),
    .A3(\shift_right_count[0] ),
    .A4(_114_),
    .ZN(_080_));
 AOI221_X2 _142_ (.A(_077_),
    .B1(_078_),
    .B2(_071_),
    .C1(_080_),
    .C2(_074_),
    .ZN(_081_));
 OR2_X1 _143_ (.A1(_066_),
    .A2(_081_),
    .ZN(_117_));
 INV_X1 _144_ (.A(_117_),
    .ZN(_120_));
 NOR2_X1 _145_ (.A1(_067_),
    .A2(_013_),
    .ZN(_082_));
 NOR2_X1 _146_ (.A1(_073_),
    .A2(_013_),
    .ZN(_083_));
 AND4_X1 _147_ (.A1(_110_),
    .A2(_067_),
    .A3(_115_),
    .A4(_070_),
    .ZN(_084_));
 AOI221_X2 _148_ (.A(_082_),
    .B1(_083_),
    .B2(_071_),
    .C1(_084_),
    .C2(_074_),
    .ZN(_085_));
 OR2_X2 _149_ (.A1(_066_),
    .A2(_085_),
    .ZN(_086_));
 MUX2_X1 _150_ (.A(_081_),
    .B(_121_),
    .S(_086_),
    .Z(_000_));
 INV_X1 _151_ (.A(_119_),
    .ZN(_087_));
 MUX2_X1 _152_ (.A(_121_),
    .B(_087_),
    .S(_086_),
    .Z(_001_));
 MUX2_X1 _153_ (.A(_087_),
    .B(_124_),
    .S(_086_),
    .Z(_002_));
 AND2_X1 _154_ (.A1(_081_),
    .A2(_085_),
    .ZN(_088_));
 AOI221_X1 _155_ (.A(_085_),
    .B1(\shift_right_count[1] ),
    .B2(_068_),
    .C1(_075_),
    .C2(_072_),
    .ZN(_029_));
 NOR3_X1 _156_ (.A1(_066_),
    .A2(_088_),
    .A3(_029_),
    .ZN(_003_));
 AOI21_X1 _157_ (.A(_066_),
    .B1(_081_),
    .B2(_085_),
    .ZN(_030_));
 OAI21_X1 _158_ (.A(_030_),
    .B1(_085_),
    .B2(_118_),
    .ZN(_004_));
 INV_X1 _159_ (.A(net1),
    .ZN(_106_));
 OR2_X1 _160_ (.A1(_066_),
    .A2(_076_),
    .ZN(_116_));
 INV_X1 _161_ (.A(net2),
    .ZN(_109_));
 INV_X1 _162_ (.A(_121_),
    .ZN(_031_));
 NAND2_X1 _163_ (.A1(_031_),
    .A2(_086_),
    .ZN(_015_));
 NAND2_X1 _164_ (.A1(_119_),
    .A2(_086_),
    .ZN(_016_));
 AOI21_X1 _165_ (.A(_066_),
    .B1(_076_),
    .B2(_085_),
    .ZN(_017_));
 BUF_X2 _166_ (.A(net11),
    .Z(_032_));
 CLKBUF_X3 _167_ (.A(_107_),
    .Z(_033_));
 MUX2_X1 _168_ (.A(_005_),
    .B(net12),
    .S(_033_),
    .Z(_034_));
 MUX2_X1 _169_ (.A(net3),
    .B(_034_),
    .S(_075_),
    .Z(_035_));
 INV_X1 _170_ (.A(_108_),
    .ZN(_036_));
 OAI21_X4 _171_ (.A(_067_),
    .B1(_036_),
    .B2(_073_),
    .ZN(_037_));
 MUX2_X1 _172_ (.A(_035_),
    .B(net13),
    .S(_037_),
    .Z(_038_));
 AND2_X1 _173_ (.A1(_032_),
    .A2(_038_),
    .ZN(_018_));
 MUX2_X1 _174_ (.A(_006_),
    .B(net13),
    .S(_033_),
    .Z(_039_));
 MUX2_X1 _175_ (.A(net4),
    .B(_039_),
    .S(_075_),
    .Z(_040_));
 MUX2_X1 _176_ (.A(_040_),
    .B(net14),
    .S(_037_),
    .Z(_041_));
 AND2_X1 _177_ (.A1(_032_),
    .A2(_041_),
    .ZN(_019_));
 MUX2_X1 _178_ (.A(_007_),
    .B(net14),
    .S(_033_),
    .Z(_042_));
 MUX2_X1 _179_ (.A(net5),
    .B(_042_),
    .S(_075_),
    .Z(_043_));
 MUX2_X1 _180_ (.A(_043_),
    .B(net15),
    .S(_037_),
    .Z(_044_));
 AND2_X1 _181_ (.A1(_032_),
    .A2(_044_),
    .ZN(_020_));
 MUX2_X1 _182_ (.A(_008_),
    .B(net15),
    .S(_033_),
    .Z(_045_));
 MUX2_X1 _183_ (.A(net6),
    .B(_045_),
    .S(_075_),
    .Z(_046_));
 MUX2_X1 _184_ (.A(_046_),
    .B(net16),
    .S(_037_),
    .Z(_047_));
 AND2_X1 _185_ (.A1(_032_),
    .A2(_047_),
    .ZN(_021_));
 MUX2_X1 _186_ (.A(_009_),
    .B(net16),
    .S(_033_),
    .Z(_048_));
 MUX2_X1 _187_ (.A(net7),
    .B(_048_),
    .S(_075_),
    .Z(_049_));
 MUX2_X1 _188_ (.A(_049_),
    .B(net17),
    .S(_037_),
    .Z(_050_));
 AND2_X1 _189_ (.A1(_032_),
    .A2(_050_),
    .ZN(_022_));
 MUX2_X1 _190_ (.A(_010_),
    .B(net17),
    .S(_033_),
    .Z(_051_));
 MUX2_X1 _191_ (.A(net8),
    .B(_051_),
    .S(_075_),
    .Z(_052_));
 MUX2_X1 _192_ (.A(_052_),
    .B(net18),
    .S(_037_),
    .Z(_053_));
 AND2_X1 _193_ (.A1(_032_),
    .A2(_053_),
    .ZN(_023_));
 MUX2_X1 _194_ (.A(_011_),
    .B(net18),
    .S(_033_),
    .Z(_054_));
 MUX2_X1 _195_ (.A(net9),
    .B(_054_),
    .S(_075_),
    .Z(_055_));
 MUX2_X1 _196_ (.A(_055_),
    .B(net19),
    .S(_037_),
    .Z(_056_));
 AND2_X1 _197_ (.A1(_032_),
    .A2(_056_),
    .ZN(_024_));
 MUX2_X1 _198_ (.A(_012_),
    .B(net19),
    .S(_033_),
    .Z(_057_));
 MUX2_X1 _199_ (.A(net10),
    .B(_057_),
    .S(_075_),
    .Z(_058_));
 MUX2_X1 _200_ (.A(_058_),
    .B(net20),
    .S(_037_),
    .Z(_059_));
 AND2_X1 _201_ (.A1(_032_),
    .A2(_059_),
    .ZN(_025_));
 NAND2_X1 _202_ (.A1(_068_),
    .A2(\shift_right_count[0] ),
    .ZN(_060_));
 AOI21_X1 _203_ (.A(_080_),
    .B1(_071_),
    .B2(\shift_right_count[0] ),
    .ZN(_061_));
 OAI21_X1 _204_ (.A(_060_),
    .B1(_061_),
    .B2(_073_),
    .ZN(_062_));
 AND2_X1 _205_ (.A1(_032_),
    .A2(_062_),
    .ZN(_026_));
 NOR2_X1 _206_ (.A1(_066_),
    .A2(_076_),
    .ZN(_027_));
 NAND2_X1 _207_ (.A1(_068_),
    .A2(\shift_right_count[2] ),
    .ZN(_063_));
 AOI21_X1 _208_ (.A(_084_),
    .B1(_071_),
    .B2(\shift_right_count[2] ),
    .ZN(_064_));
 OAI21_X1 _209_ (.A(_063_),
    .B1(_064_),
    .B2(_073_),
    .ZN(_065_));
 AND2_X1 _210_ (.A1(_032_),
    .A2(_065_),
    .ZN(_028_));
 HA_X1 _211_ (.A(_106_),
    .B(net2),
    .CO(_107_),
    .S(_108_));
 HA_X1 _212_ (.A(net1),
    .B(_109_),
    .CO(_110_),
    .S(_111_));
 HA_X1 _213_ (.A(\shift_right_count[0] ),
    .B(\shift_right_count[1] ),
    .CO(_112_),
    .S(_113_));
 HA_X1 _214_ (.A(\shift_right_count[2] ),
    .B(_112_),
    .CO(_114_),
    .S(_115_));
 HA_X1 _215_ (.A(_116_),
    .B(_117_),
    .CO(_118_),
    .S(_119_));
 HA_X1 _216_ (.A(_116_),
    .B(_120_),
    .CO(_121_),
    .S(_122_));
 HA_X1 _217_ (.A(_123_),
    .B(_117_),
    .CO(_124_),
    .S(_125_));
 DFF_X1 _218_ (.D(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(_005_),
    .QN(_102_));
 DFF_X1 _219_ (.D(_001_),
    .CK(clknet_1_0__leaf_clk),
    .Q(_006_),
    .QN(_103_));
 DFF_X1 _220_ (.D(_002_),
    .CK(clknet_1_0__leaf_clk),
    .Q(_007_),
    .QN(_104_));
 DFF_X1 _221_ (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(_008_),
    .QN(_105_));
 DFF_X1 _222_ (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(_009_),
    .QN(_101_));
 DFF_X1 _223_ (.D(_015_),
    .CK(clknet_1_0__leaf_clk),
    .Q(_010_),
    .QN(_100_));
 DFF_X1 _224_ (.D(_016_),
    .CK(clknet_1_0__leaf_clk),
    .Q(_011_),
    .QN(_099_));
 DFF_X1 _225_ (.D(_017_),
    .CK(clknet_1_1__leaf_clk),
    .Q(_012_),
    .QN(_098_));
 DFF_X1 \parallel_out[0]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net13),
    .QN(_097_));
 DFF_X1 \parallel_out[1]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net14),
    .QN(_096_));
 DFF_X1 \parallel_out[2]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net15),
    .QN(_095_));
 DFF_X1 \parallel_out[3]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net16),
    .QN(_094_));
 DFF_X1 \parallel_out[4]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net17),
    .QN(_093_));
 DFF_X1 \parallel_out[5]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net18),
    .QN(_092_));
 DFF_X1 \parallel_out[6]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net19),
    .QN(_091_));
 DFF_X1 \parallel_out[7]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net20),
    .QN(_090_));
 DFF_X2 \shift_right_count[0]$_SDFFE_PN0N_  (.D(_026_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_right_count[0] ),
    .QN(_014_));
 DFF_X2 \shift_right_count[1]$_SDFFE_PN0N_  (.D(_027_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_right_count[1] ),
    .QN(_089_));
 DFF_X1 \shift_right_count[2]$_SDFFE_PN0N_  (.D(_028_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_right_count[2] ),
    .QN(_013_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_91 ();
 BUF_X1 input1 (.A(direction[0]),
    .Z(net1));
 BUF_X1 input2 (.A(direction[1]),
    .Z(net2));
 BUF_X1 input3 (.A(parallel_in[0]),
    .Z(net3));
 BUF_X1 input4 (.A(parallel_in[1]),
    .Z(net4));
 BUF_X1 input5 (.A(parallel_in[2]),
    .Z(net5));
 BUF_X1 input6 (.A(parallel_in[3]),
    .Z(net6));
 BUF_X1 input7 (.A(parallel_in[4]),
    .Z(net7));
 BUF_X1 input8 (.A(parallel_in[5]),
    .Z(net8));
 BUF_X1 input9 (.A(parallel_in[6]),
    .Z(net9));
 BUF_X1 input10 (.A(parallel_in[7]),
    .Z(net10));
 BUF_X1 input11 (.A(rst_n),
    .Z(net11));
 BUF_X1 input12 (.A(serial_in_right),
    .Z(net12));
 BUF_X1 output13 (.A(net13),
    .Z(parallel_out[0]));
 BUF_X1 output14 (.A(net14),
    .Z(parallel_out[1]));
 BUF_X1 output15 (.A(net15),
    .Z(parallel_out[2]));
 BUF_X1 output16 (.A(net16),
    .Z(parallel_out[3]));
 BUF_X1 output17 (.A(net17),
    .Z(parallel_out[4]));
 BUF_X1 output18 (.A(net18),
    .Z(parallel_out[5]));
 BUF_X1 output19 (.A(net19),
    .Z(parallel_out[6]));
 BUF_X1 output20 (.A(net20),
    .Z(parallel_out[7]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 INV_X2 clkload0 (.A(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X16 FILLER_0_129 ();
 FILLCELL_X8 FILLER_0_145 ();
 FILLCELL_X4 FILLER_0_153 ();
 FILLCELL_X2 FILLER_0_157 ();
 FILLCELL_X1 FILLER_0_159 ();
 FILLCELL_X2 FILLER_0_163 ();
 FILLCELL_X1 FILLER_0_165 ();
 FILLCELL_X2 FILLER_0_172 ();
 FILLCELL_X8 FILLER_0_177 ();
 FILLCELL_X4 FILLER_0_185 ();
 FILLCELL_X16 FILLER_0_192 ();
 FILLCELL_X2 FILLER_0_208 ();
 FILLCELL_X32 FILLER_0_219 ();
 FILLCELL_X32 FILLER_0_251 ();
 FILLCELL_X32 FILLER_0_283 ();
 FILLCELL_X16 FILLER_0_315 ();
 FILLCELL_X8 FILLER_0_331 ();
 FILLCELL_X4 FILLER_0_339 ();
 FILLCELL_X2 FILLER_0_343 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X16 FILLER_1_321 ();
 FILLCELL_X8 FILLER_1_337 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X16 FILLER_2_321 ();
 FILLCELL_X8 FILLER_2_337 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X16 FILLER_3_321 ();
 FILLCELL_X8 FILLER_3_337 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X16 FILLER_4_321 ();
 FILLCELL_X8 FILLER_4_337 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X16 FILLER_5_321 ();
 FILLCELL_X8 FILLER_5_337 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X16 FILLER_6_321 ();
 FILLCELL_X8 FILLER_6_337 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X16 FILLER_7_321 ();
 FILLCELL_X8 FILLER_7_337 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X16 FILLER_8_321 ();
 FILLCELL_X8 FILLER_8_337 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X16 FILLER_9_321 ();
 FILLCELL_X8 FILLER_9_337 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X2 FILLER_10_161 ();
 FILLCELL_X1 FILLER_10_163 ();
 FILLCELL_X8 FILLER_10_178 ();
 FILLCELL_X4 FILLER_10_186 ();
 FILLCELL_X32 FILLER_10_207 ();
 FILLCELL_X32 FILLER_10_239 ();
 FILLCELL_X32 FILLER_10_271 ();
 FILLCELL_X32 FILLER_10_303 ();
 FILLCELL_X8 FILLER_10_335 ();
 FILLCELL_X2 FILLER_10_343 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X16 FILLER_11_129 ();
 FILLCELL_X8 FILLER_11_145 ();
 FILLCELL_X4 FILLER_11_153 ();
 FILLCELL_X2 FILLER_11_157 ();
 FILLCELL_X1 FILLER_11_159 ();
 FILLCELL_X4 FILLER_11_181 ();
 FILLCELL_X16 FILLER_11_196 ();
 FILLCELL_X32 FILLER_11_226 ();
 FILLCELL_X32 FILLER_11_258 ();
 FILLCELL_X32 FILLER_11_290 ();
 FILLCELL_X16 FILLER_11_322 ();
 FILLCELL_X4 FILLER_11_338 ();
 FILLCELL_X2 FILLER_11_342 ();
 FILLCELL_X1 FILLER_11_344 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X2 FILLER_12_161 ();
 FILLCELL_X1 FILLER_12_163 ();
 FILLCELL_X2 FILLER_12_171 ();
 FILLCELL_X1 FILLER_12_173 ();
 FILLCELL_X8 FILLER_12_188 ();
 FILLCELL_X4 FILLER_12_196 ();
 FILLCELL_X2 FILLER_12_200 ();
 FILLCELL_X1 FILLER_12_202 ();
 FILLCELL_X32 FILLER_12_224 ();
 FILLCELL_X32 FILLER_12_256 ();
 FILLCELL_X32 FILLER_12_288 ();
 FILLCELL_X16 FILLER_12_320 ();
 FILLCELL_X8 FILLER_12_336 ();
 FILLCELL_X1 FILLER_12_344 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X16 FILLER_13_321 ();
 FILLCELL_X8 FILLER_13_337 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X16 FILLER_14_161 ();
 FILLCELL_X4 FILLER_14_177 ();
 FILLCELL_X16 FILLER_14_198 ();
 FILLCELL_X1 FILLER_14_214 ();
 FILLCELL_X32 FILLER_14_229 ();
 FILLCELL_X32 FILLER_14_261 ();
 FILLCELL_X32 FILLER_14_293 ();
 FILLCELL_X16 FILLER_14_325 ();
 FILLCELL_X4 FILLER_14_341 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X1 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_179 ();
 FILLCELL_X16 FILLER_15_211 ();
 FILLCELL_X1 FILLER_15_227 ();
 FILLCELL_X32 FILLER_15_239 ();
 FILLCELL_X32 FILLER_15_271 ();
 FILLCELL_X32 FILLER_15_303 ();
 FILLCELL_X8 FILLER_15_335 ();
 FILLCELL_X2 FILLER_15_343 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X2 FILLER_16_161 ();
 FILLCELL_X16 FILLER_16_180 ();
 FILLCELL_X4 FILLER_16_196 ();
 FILLCELL_X2 FILLER_16_200 ();
 FILLCELL_X16 FILLER_16_207 ();
 FILLCELL_X8 FILLER_16_223 ();
 FILLCELL_X4 FILLER_16_231 ();
 FILLCELL_X32 FILLER_16_252 ();
 FILLCELL_X32 FILLER_16_284 ();
 FILLCELL_X16 FILLER_16_316 ();
 FILLCELL_X8 FILLER_16_332 ();
 FILLCELL_X4 FILLER_16_340 ();
 FILLCELL_X1 FILLER_16_344 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X4 FILLER_17_161 ();
 FILLCELL_X2 FILLER_17_165 ();
 FILLCELL_X2 FILLER_17_174 ();
 FILLCELL_X32 FILLER_17_181 ();
 FILLCELL_X32 FILLER_17_213 ();
 FILLCELL_X32 FILLER_17_245 ();
 FILLCELL_X16 FILLER_17_277 ();
 FILLCELL_X8 FILLER_17_293 ();
 FILLCELL_X4 FILLER_17_301 ();
 FILLCELL_X1 FILLER_17_305 ();
 FILLCELL_X32 FILLER_17_309 ();
 FILLCELL_X4 FILLER_17_341 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X4 FILLER_18_161 ();
 FILLCELL_X2 FILLER_18_165 ();
 FILLCELL_X1 FILLER_18_227 ();
 FILLCELL_X32 FILLER_18_235 ();
 FILLCELL_X32 FILLER_18_267 ();
 FILLCELL_X32 FILLER_18_299 ();
 FILLCELL_X8 FILLER_18_331 ();
 FILLCELL_X4 FILLER_18_339 ();
 FILLCELL_X2 FILLER_18_343 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X2 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_165 ();
 FILLCELL_X32 FILLER_19_179 ();
 FILLCELL_X32 FILLER_19_211 ();
 FILLCELL_X32 FILLER_19_243 ();
 FILLCELL_X32 FILLER_19_275 ();
 FILLCELL_X32 FILLER_19_307 ();
 FILLCELL_X4 FILLER_19_339 ();
 FILLCELL_X2 FILLER_19_343 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X8 FILLER_20_181 ();
 FILLCELL_X4 FILLER_20_189 ();
 FILLCELL_X2 FILLER_20_193 ();
 FILLCELL_X8 FILLER_20_219 ();
 FILLCELL_X2 FILLER_20_227 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X16 FILLER_20_289 ();
 FILLCELL_X1 FILLER_20_305 ();
 FILLCELL_X32 FILLER_20_309 ();
 FILLCELL_X4 FILLER_20_341 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X2 FILLER_21_161 ();
 FILLCELL_X2 FILLER_21_174 ();
 FILLCELL_X1 FILLER_21_176 ();
 FILLCELL_X8 FILLER_21_186 ();
 FILLCELL_X4 FILLER_21_194 ();
 FILLCELL_X2 FILLER_21_198 ();
 FILLCELL_X16 FILLER_21_205 ();
 FILLCELL_X4 FILLER_21_221 ();
 FILLCELL_X32 FILLER_21_232 ();
 FILLCELL_X32 FILLER_21_264 ();
 FILLCELL_X8 FILLER_21_296 ();
 FILLCELL_X2 FILLER_21_304 ();
 FILLCELL_X32 FILLER_21_309 ();
 FILLCELL_X4 FILLER_21_341 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X16 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_181 ();
 FILLCELL_X16 FILLER_22_213 ();
 FILLCELL_X4 FILLER_22_229 ();
 FILLCELL_X32 FILLER_22_244 ();
 FILLCELL_X32 FILLER_22_276 ();
 FILLCELL_X32 FILLER_22_308 ();
 FILLCELL_X4 FILLER_22_340 ();
 FILLCELL_X1 FILLER_22_344 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X1 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X16 FILLER_23_289 ();
 FILLCELL_X4 FILLER_23_305 ();
 FILLCELL_X8 FILLER_23_312 ();
 FILLCELL_X2 FILLER_23_320 ();
 FILLCELL_X16 FILLER_23_325 ();
 FILLCELL_X4 FILLER_23_341 ();
 FILLCELL_X16 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_17 ();
 FILLCELL_X32 FILLER_24_22 ();
 FILLCELL_X32 FILLER_24_54 ();
 FILLCELL_X32 FILLER_24_86 ();
 FILLCELL_X32 FILLER_24_118 ();
 FILLCELL_X8 FILLER_24_150 ();
 FILLCELL_X2 FILLER_24_165 ();
 FILLCELL_X1 FILLER_24_167 ();
 FILLCELL_X4 FILLER_24_171 ();
 FILLCELL_X2 FILLER_24_175 ();
 FILLCELL_X1 FILLER_24_177 ();
 FILLCELL_X4 FILLER_24_186 ();
 FILLCELL_X2 FILLER_24_190 ();
 FILLCELL_X1 FILLER_24_192 ();
 FILLCELL_X32 FILLER_24_210 ();
 FILLCELL_X32 FILLER_24_242 ();
 FILLCELL_X32 FILLER_24_274 ();
 FILLCELL_X32 FILLER_24_306 ();
 FILLCELL_X4 FILLER_24_338 ();
 FILLCELL_X2 FILLER_24_342 ();
 FILLCELL_X1 FILLER_24_344 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X16 FILLER_25_129 ();
 FILLCELL_X8 FILLER_25_145 ();
 FILLCELL_X4 FILLER_25_153 ();
 FILLCELL_X4 FILLER_25_176 ();
 FILLCELL_X32 FILLER_25_184 ();
 FILLCELL_X32 FILLER_25_216 ();
 FILLCELL_X32 FILLER_25_248 ();
 FILLCELL_X32 FILLER_25_280 ();
 FILLCELL_X32 FILLER_25_312 ();
 FILLCELL_X1 FILLER_25_344 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X1 FILLER_26_184 ();
 FILLCELL_X16 FILLER_26_210 ();
 FILLCELL_X4 FILLER_26_226 ();
 FILLCELL_X2 FILLER_26_230 ();
 FILLCELL_X32 FILLER_26_243 ();
 FILLCELL_X16 FILLER_26_275 ();
 FILLCELL_X8 FILLER_26_291 ();
 FILLCELL_X4 FILLER_26_299 ();
 FILLCELL_X2 FILLER_26_303 ();
 FILLCELL_X1 FILLER_26_305 ();
 FILLCELL_X32 FILLER_26_309 ();
 FILLCELL_X4 FILLER_26_341 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X16 FILLER_27_129 ();
 FILLCELL_X8 FILLER_27_145 ();
 FILLCELL_X1 FILLER_27_153 ();
 FILLCELL_X2 FILLER_27_173 ();
 FILLCELL_X16 FILLER_27_186 ();
 FILLCELL_X8 FILLER_27_202 ();
 FILLCELL_X4 FILLER_27_210 ();
 FILLCELL_X2 FILLER_27_214 ();
 FILLCELL_X1 FILLER_27_216 ();
 FILLCELL_X8 FILLER_27_224 ();
 FILLCELL_X32 FILLER_27_256 ();
 FILLCELL_X16 FILLER_27_288 ();
 FILLCELL_X2 FILLER_27_304 ();
 FILLCELL_X1 FILLER_27_306 ();
 FILLCELL_X32 FILLER_27_310 ();
 FILLCELL_X2 FILLER_27_342 ();
 FILLCELL_X1 FILLER_27_344 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X16 FILLER_28_129 ();
 FILLCELL_X8 FILLER_28_145 ();
 FILLCELL_X4 FILLER_28_153 ();
 FILLCELL_X2 FILLER_28_157 ();
 FILLCELL_X32 FILLER_28_190 ();
 FILLCELL_X32 FILLER_28_222 ();
 FILLCELL_X32 FILLER_28_254 ();
 FILLCELL_X32 FILLER_28_286 ();
 FILLCELL_X16 FILLER_28_318 ();
 FILLCELL_X8 FILLER_28_334 ();
 FILLCELL_X2 FILLER_28_342 ();
 FILLCELL_X1 FILLER_28_344 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X1 FILLER_29_161 ();
 FILLCELL_X1 FILLER_29_172 ();
 FILLCELL_X16 FILLER_29_193 ();
 FILLCELL_X8 FILLER_29_209 ();
 FILLCELL_X1 FILLER_29_217 ();
 FILLCELL_X1 FILLER_29_236 ();
 FILLCELL_X32 FILLER_29_254 ();
 FILLCELL_X16 FILLER_29_286 ();
 FILLCELL_X4 FILLER_29_302 ();
 FILLCELL_X32 FILLER_29_309 ();
 FILLCELL_X4 FILLER_29_341 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X16 FILLER_30_129 ();
 FILLCELL_X8 FILLER_30_145 ();
 FILLCELL_X4 FILLER_30_153 ();
 FILLCELL_X1 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_192 ();
 FILLCELL_X32 FILLER_30_224 ();
 FILLCELL_X32 FILLER_30_256 ();
 FILLCELL_X32 FILLER_30_288 ();
 FILLCELL_X16 FILLER_30_320 ();
 FILLCELL_X8 FILLER_30_336 ();
 FILLCELL_X1 FILLER_30_344 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X8 FILLER_31_129 ();
 FILLCELL_X4 FILLER_31_137 ();
 FILLCELL_X1 FILLER_31_141 ();
 FILLCELL_X4 FILLER_31_159 ();
 FILLCELL_X1 FILLER_31_166 ();
 FILLCELL_X1 FILLER_31_170 ();
 FILLCELL_X32 FILLER_31_191 ();
 FILLCELL_X32 FILLER_31_223 ();
 FILLCELL_X32 FILLER_31_255 ();
 FILLCELL_X32 FILLER_31_287 ();
 FILLCELL_X16 FILLER_31_319 ();
 FILLCELL_X8 FILLER_31_335 ();
 FILLCELL_X2 FILLER_31_343 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X16 FILLER_32_321 ();
 FILLCELL_X8 FILLER_32_337 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X16 FILLER_33_321 ();
 FILLCELL_X8 FILLER_33_337 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X4 FILLER_34_161 ();
 FILLCELL_X1 FILLER_34_165 ();
 FILLCELL_X4 FILLER_34_179 ();
 FILLCELL_X2 FILLER_34_183 ();
 FILLCELL_X1 FILLER_34_185 ();
 FILLCELL_X32 FILLER_34_191 ();
 FILLCELL_X32 FILLER_34_223 ();
 FILLCELL_X32 FILLER_34_255 ();
 FILLCELL_X32 FILLER_34_287 ();
 FILLCELL_X16 FILLER_34_319 ();
 FILLCELL_X8 FILLER_34_335 ();
 FILLCELL_X2 FILLER_34_343 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X8 FILLER_35_161 ();
 FILLCELL_X4 FILLER_35_169 ();
 FILLCELL_X1 FILLER_35_173 ();
 FILLCELL_X4 FILLER_35_176 ();
 FILLCELL_X2 FILLER_35_180 ();
 FILLCELL_X1 FILLER_35_182 ();
 FILLCELL_X32 FILLER_35_195 ();
 FILLCELL_X32 FILLER_35_227 ();
 FILLCELL_X32 FILLER_35_259 ();
 FILLCELL_X32 FILLER_35_291 ();
 FILLCELL_X16 FILLER_35_323 ();
 FILLCELL_X4 FILLER_35_339 ();
 FILLCELL_X2 FILLER_35_343 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X16 FILLER_36_161 ();
 FILLCELL_X1 FILLER_36_177 ();
 FILLCELL_X32 FILLER_36_190 ();
 FILLCELL_X32 FILLER_36_222 ();
 FILLCELL_X32 FILLER_36_254 ();
 FILLCELL_X32 FILLER_36_286 ();
 FILLCELL_X16 FILLER_36_318 ();
 FILLCELL_X8 FILLER_36_334 ();
 FILLCELL_X2 FILLER_36_342 ();
 FILLCELL_X1 FILLER_36_344 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X4 FILLER_37_161 ();
 FILLCELL_X2 FILLER_37_165 ();
 FILLCELL_X1 FILLER_37_167 ();
 FILLCELL_X32 FILLER_37_176 ();
 FILLCELL_X32 FILLER_37_208 ();
 FILLCELL_X32 FILLER_37_240 ();
 FILLCELL_X32 FILLER_37_272 ();
 FILLCELL_X32 FILLER_37_304 ();
 FILLCELL_X8 FILLER_37_336 ();
 FILLCELL_X1 FILLER_37_344 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X16 FILLER_38_321 ();
 FILLCELL_X8 FILLER_38_337 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X16 FILLER_39_321 ();
 FILLCELL_X8 FILLER_39_337 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X16 FILLER_40_321 ();
 FILLCELL_X8 FILLER_40_337 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X16 FILLER_41_321 ();
 FILLCELL_X8 FILLER_41_337 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X16 FILLER_42_321 ();
 FILLCELL_X8 FILLER_42_337 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X16 FILLER_43_321 ();
 FILLCELL_X8 FILLER_43_337 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X16 FILLER_44_321 ();
 FILLCELL_X8 FILLER_44_337 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X16 FILLER_45_161 ();
 FILLCELL_X4 FILLER_45_177 ();
 FILLCELL_X1 FILLER_45_181 ();
 FILLCELL_X1 FILLER_45_185 ();
 FILLCELL_X16 FILLER_45_189 ();
 FILLCELL_X4 FILLER_45_205 ();
 FILLCELL_X1 FILLER_45_209 ();
 FILLCELL_X32 FILLER_45_213 ();
 FILLCELL_X32 FILLER_45_245 ();
 FILLCELL_X32 FILLER_45_277 ();
 FILLCELL_X32 FILLER_45_309 ();
 FILLCELL_X4 FILLER_45_341 ();
endmodule
