module parameterized_onehot_counter (clk,
    enable,
    rst_n,
    count);
 input clk;
 input enable;
 input rst_n;
 output [7:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16_ (.I0(net4),
    .I1(net11),
    .S(net2),
    .Z(_00_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _17_ (.I(net11),
    .ZN(_08_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18_ (.A1(net4),
    .A2(_08_),
    .Z(_09_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19_ (.I0(net5),
    .I1(_09_),
    .S(net2),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20_ (.A1(_08_),
    .A2(net5),
    .Z(_10_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21_ (.I0(net6),
    .I1(_10_),
    .S(net2),
    .Z(_02_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22_ (.A1(_08_),
    .A2(net6),
    .Z(_11_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _23_ (.I0(net7),
    .I1(_11_),
    .S(net2),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24_ (.A1(_08_),
    .A2(net7),
    .Z(_12_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _25_ (.I0(net8),
    .I1(_12_),
    .S(net2),
    .Z(_04_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26_ (.A1(_08_),
    .A2(net8),
    .Z(_13_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _27_ (.I0(net9),
    .I1(_13_),
    .S(net2),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28_ (.A1(_08_),
    .A2(net9),
    .Z(_14_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _29_ (.I0(net10),
    .I1(_14_),
    .S(net2),
    .Z(_06_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30_ (.A1(_08_),
    .A2(net10),
    .Z(_15_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31_ (.I0(net11),
    .I1(_15_),
    .S(net2),
    .Z(_07_));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \counter_reg[0]$_DFFE_PN1P_  (.D(_00_),
    .SETN(net3),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[1]$_DFFE_PN0P_  (.D(_01_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[2]$_DFFE_PN0P_  (.D(_02_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[3]$_DFFE_PN0P_  (.D(_03_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[4]$_DFFE_PN0P_  (.D(_04_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net8));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[5]$_DFFE_PN0P_  (.D(_05_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net9));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[6]$_DFFE_PN0P_  (.D(_06_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net10));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[7]$_DFFE_PN0P_  (.D(_07_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 hold1 (.I(net3),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_44 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_55 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input1 (.I(enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(rst_n),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output3 (.I(net4),
    .Z(count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output4 (.I(net5),
    .Z(count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output5 (.I(net6),
    .Z(count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output6 (.I(net7),
    .Z(count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output7 (.I(net8),
    .Z(count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output8 (.I(net9),
    .Z(count[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output9 (.I(net10),
    .Z(count[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output10 (.I(net11),
    .Z(count[7]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 clkload0 (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_196 ();
endmodule
