module parameterized_crc_generator (clk,
    crc_init,
    data_valid,
    rst_n,
    crc_out,
    data_in);
 input clk;
 input crc_init;
 input data_valid;
 input rst_n;
 output [7:0] crc_out;
 input [7:0] data_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire \crc_reflected[0] ;
 wire \crc_reflected[1] ;
 wire \crc_reflected[2] ;
 wire \crc_reflected[3] ;
 wire \crc_reflected[4] ;
 wire \crc_reflected[5] ;
 wire \crc_reflected[6] ;
 wire \crc_reflected[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X4 _085_ (.A(crc_init),
    .Z(_016_));
 INV_X1 _086_ (.A(net9),
    .ZN(_017_));
 NOR2_X2 _087_ (.A1(_016_),
    .A2(_017_),
    .ZN(_018_));
 XOR2_X2 _088_ (.A(\crc_reflected[0] ),
    .B(net1),
    .Z(_019_));
 BUF_X4 _089_ (.A(\crc_reflected[6] ),
    .Z(_020_));
 XNOR2_X1 _090_ (.A(net7),
    .B(_020_),
    .ZN(_021_));
 XNOR2_X2 _091_ (.A(_019_),
    .B(_021_),
    .ZN(_022_));
 XNOR2_X2 _092_ (.A(net8),
    .B(\crc_reflected[7] ),
    .ZN(_023_));
 XNOR2_X1 _093_ (.A(_022_),
    .B(_023_),
    .ZN(_024_));
 BUF_X2 _094_ (.A(data_valid),
    .Z(_025_));
 MUX2_X1 _095_ (.A(\crc_reflected[0] ),
    .B(_024_),
    .S(_025_),
    .Z(_026_));
 AND2_X1 _096_ (.A1(_018_),
    .A2(_026_),
    .ZN(_008_));
 CLKBUF_X3 _097_ (.A(_017_),
    .Z(_027_));
 INV_X1 _098_ (.A(\crc_reflected[1] ),
    .ZN(_028_));
 NOR3_X1 _099_ (.A1(_016_),
    .A2(_027_),
    .A3(_028_),
    .ZN(_029_));
 NOR3_X1 _100_ (.A1(_016_),
    .A2(_027_),
    .A3(\crc_reflected[1] ),
    .ZN(_030_));
 INV_X1 _101_ (.A(_025_),
    .ZN(_031_));
 XNOR2_X1 _102_ (.A(net2),
    .B(_022_),
    .ZN(_032_));
 NOR2_X1 _103_ (.A1(_031_),
    .A2(_032_),
    .ZN(_033_));
 MUX2_X1 _104_ (.A(_029_),
    .B(_030_),
    .S(_033_),
    .Z(_009_));
 OR2_X1 _105_ (.A1(\crc_reflected[2] ),
    .A2(_025_),
    .ZN(_034_));
 XNOR2_X1 _106_ (.A(net3),
    .B(\crc_reflected[2] ),
    .ZN(_035_));
 XOR2_X1 _107_ (.A(\crc_reflected[1] ),
    .B(net2),
    .Z(_036_));
 XNOR2_X1 _108_ (.A(_035_),
    .B(_036_),
    .ZN(_037_));
 XNOR2_X1 _109_ (.A(_022_),
    .B(_037_),
    .ZN(_038_));
 NAND2_X1 _110_ (.A1(_025_),
    .A2(_038_),
    .ZN(_039_));
 AND3_X1 _111_ (.A1(_018_),
    .A2(_034_),
    .A3(_039_),
    .ZN(_010_));
 INV_X1 _112_ (.A(\crc_reflected[3] ),
    .ZN(_040_));
 NOR3_X1 _113_ (.A1(_016_),
    .A2(_017_),
    .A3(_040_),
    .ZN(_041_));
 NOR3_X1 _114_ (.A1(_016_),
    .A2(_027_),
    .A3(\crc_reflected[3] ),
    .ZN(_042_));
 XNOR2_X1 _115_ (.A(net4),
    .B(_023_),
    .ZN(_043_));
 XNOR2_X1 _116_ (.A(_037_),
    .B(_043_),
    .ZN(_044_));
 NOR2_X1 _117_ (.A1(_031_),
    .A2(_044_),
    .ZN(_045_));
 MUX2_X1 _118_ (.A(_041_),
    .B(_042_),
    .S(_045_),
    .Z(_011_));
 XOR2_X2 _119_ (.A(net5),
    .B(\crc_reflected[4] ),
    .Z(_046_));
 XNOR2_X1 _120_ (.A(net4),
    .B(\crc_reflected[3] ),
    .ZN(_047_));
 XNOR2_X2 _121_ (.A(_046_),
    .B(_047_),
    .ZN(_048_));
 XNOR2_X1 _122_ (.A(_035_),
    .B(_048_),
    .ZN(_049_));
 MUX2_X1 _123_ (.A(\crc_reflected[4] ),
    .B(_049_),
    .S(_025_),
    .Z(_050_));
 AND2_X1 _124_ (.A1(_018_),
    .A2(_050_),
    .ZN(_012_));
 INV_X1 _125_ (.A(\crc_reflected[5] ),
    .ZN(_051_));
 NOR3_X1 _126_ (.A1(_016_),
    .A2(_017_),
    .A3(_051_),
    .ZN(_052_));
 NOR3_X1 _127_ (.A1(_016_),
    .A2(_027_),
    .A3(\crc_reflected[5] ),
    .ZN(_053_));
 XNOR2_X1 _128_ (.A(net6),
    .B(_048_),
    .ZN(_054_));
 NOR2_X1 _129_ (.A1(_031_),
    .A2(_054_),
    .ZN(_055_));
 MUX2_X1 _130_ (.A(_052_),
    .B(_053_),
    .S(_055_),
    .Z(_013_));
 INV_X1 _131_ (.A(_020_),
    .ZN(_056_));
 NOR3_X1 _132_ (.A1(_016_),
    .A2(_017_),
    .A3(_056_),
    .ZN(_057_));
 NOR3_X1 _133_ (.A1(_016_),
    .A2(_027_),
    .A3(_020_),
    .ZN(_058_));
 XNOR2_X2 _134_ (.A(net6),
    .B(\crc_reflected[5] ),
    .ZN(_059_));
 XNOR2_X2 _135_ (.A(net7),
    .B(_059_),
    .ZN(_060_));
 XNOR2_X1 _136_ (.A(_046_),
    .B(_060_),
    .ZN(_061_));
 NOR2_X1 _137_ (.A1(_031_),
    .A2(_061_),
    .ZN(_062_));
 MUX2_X1 _138_ (.A(_057_),
    .B(_058_),
    .S(_062_),
    .Z(_014_));
 NAND2_X1 _139_ (.A1(\crc_reflected[7] ),
    .A2(_018_),
    .ZN(_063_));
 XNOR2_X1 _140_ (.A(net8),
    .B(_020_),
    .ZN(_064_));
 XNOR2_X1 _141_ (.A(_060_),
    .B(_064_),
    .ZN(_065_));
 AOI21_X1 _142_ (.A(_063_),
    .B1(_065_),
    .B2(_025_),
    .ZN(_066_));
 INV_X1 _143_ (.A(\crc_reflected[7] ),
    .ZN(_067_));
 AND4_X1 _144_ (.A1(_067_),
    .A2(_025_),
    .A3(_018_),
    .A4(_065_),
    .ZN(_068_));
 OR2_X1 _145_ (.A1(_066_),
    .A2(_068_),
    .ZN(_015_));
 AND2_X1 _146_ (.A1(net9),
    .A2(\crc_reflected[0] ),
    .ZN(_000_));
 NOR2_X1 _147_ (.A1(_027_),
    .A2(_028_),
    .ZN(_001_));
 AND2_X1 _148_ (.A1(net9),
    .A2(\crc_reflected[2] ),
    .ZN(_002_));
 NOR2_X1 _149_ (.A1(_027_),
    .A2(_040_),
    .ZN(_003_));
 AND2_X1 _150_ (.A1(net9),
    .A2(\crc_reflected[4] ),
    .ZN(_004_));
 NOR2_X1 _151_ (.A1(_027_),
    .A2(_051_),
    .ZN(_005_));
 NOR2_X1 _152_ (.A1(_027_),
    .A2(_056_),
    .ZN(_006_));
 NOR2_X1 _153_ (.A1(_027_),
    .A2(_067_),
    .ZN(_007_));
 DFF_X1 \crc_out[0]$_SDFF_PN0_  (.D(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net10),
    .QN(_084_));
 DFF_X1 \crc_out[1]$_SDFF_PN0_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net11),
    .QN(_083_));
 DFF_X1 \crc_out[2]$_SDFF_PN0_  (.D(_002_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net12),
    .QN(_082_));
 DFF_X1 \crc_out[3]$_SDFF_PN0_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net13),
    .QN(_081_));
 DFF_X1 \crc_out[4]$_SDFF_PN0_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net14),
    .QN(_080_));
 DFF_X1 \crc_out[5]$_SDFF_PN0_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net15),
    .QN(_079_));
 DFF_X1 \crc_out[6]$_SDFF_PN0_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net16),
    .QN(_078_));
 DFF_X1 \crc_out[7]$_SDFF_PN0_  (.D(_007_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net17),
    .QN(_077_));
 DFF_X1 \crc_reg[0]$_SDFFE_PP0P_  (.D(_008_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\crc_reflected[0] ),
    .QN(_076_));
 DFF_X1 \crc_reg[1]$_SDFFE_PP0P_  (.D(_009_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\crc_reflected[1] ),
    .QN(_075_));
 DFF_X1 \crc_reg[2]$_SDFFE_PP0P_  (.D(_010_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\crc_reflected[2] ),
    .QN(_074_));
 DFF_X1 \crc_reg[3]$_SDFFE_PP0P_  (.D(_011_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\crc_reflected[3] ),
    .QN(_073_));
 DFF_X1 \crc_reg[4]$_SDFFE_PP0P_  (.D(_012_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\crc_reflected[4] ),
    .QN(_072_));
 DFF_X2 \crc_reg[5]$_SDFFE_PP0P_  (.D(_013_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\crc_reflected[5] ),
    .QN(_071_));
 DFF_X1 \crc_reg[6]$_SDFFE_PP0P_  (.D(_014_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\crc_reflected[6] ),
    .QN(_070_));
 DFF_X1 \crc_reg[7]$_SDFFE_PP0P_  (.D(_015_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\crc_reflected[7] ),
    .QN(_069_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_55 ();
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[2]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[3]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[5]),
    .Z(net6));
 BUF_X1 input7 (.A(data_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[7]),
    .Z(net8));
 BUF_X1 input9 (.A(rst_n),
    .Z(net9));
 BUF_X1 output10 (.A(net10),
    .Z(crc_out[0]));
 BUF_X1 output11 (.A(net11),
    .Z(crc_out[1]));
 BUF_X1 output12 (.A(net12),
    .Z(crc_out[2]));
 BUF_X1 output13 (.A(net13),
    .Z(crc_out[3]));
 BUF_X1 output14 (.A(net14),
    .Z(crc_out[4]));
 BUF_X1 output15 (.A(net15),
    .Z(crc_out[5]));
 BUF_X1 output16 (.A(net16),
    .Z(crc_out[6]));
 BUF_X1 output17 (.A(net17),
    .Z(crc_out[7]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_73 ();
 FILLCELL_X8 FILLER_0_80 ();
 FILLCELL_X4 FILLER_0_88 ();
 FILLCELL_X16 FILLER_0_95 ();
 FILLCELL_X1 FILLER_0_111 ();
 FILLCELL_X8 FILLER_0_115 ();
 FILLCELL_X4 FILLER_0_123 ();
 FILLCELL_X8 FILLER_0_130 ();
 FILLCELL_X4 FILLER_0_138 ();
 FILLCELL_X1 FILLER_0_142 ();
 FILLCELL_X32 FILLER_0_146 ();
 FILLCELL_X32 FILLER_0_178 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X16 FILLER_1_65 ();
 FILLCELL_X1 FILLER_1_81 ();
 FILLCELL_X32 FILLER_1_85 ();
 FILLCELL_X32 FILLER_1_117 ();
 FILLCELL_X32 FILLER_1_149 ();
 FILLCELL_X16 FILLER_1_181 ();
 FILLCELL_X8 FILLER_1_197 ();
 FILLCELL_X4 FILLER_1_205 ();
 FILLCELL_X1 FILLER_1_209 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X16 FILLER_2_193 ();
 FILLCELL_X1 FILLER_2_209 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_65 ();
 FILLCELL_X4 FILLER_3_73 ();
 FILLCELL_X1 FILLER_3_77 ();
 FILLCELL_X16 FILLER_3_95 ();
 FILLCELL_X8 FILLER_3_111 ();
 FILLCELL_X4 FILLER_3_119 ();
 FILLCELL_X2 FILLER_3_123 ();
 FILLCELL_X1 FILLER_3_125 ();
 FILLCELL_X32 FILLER_3_143 ();
 FILLCELL_X32 FILLER_3_175 ();
 FILLCELL_X2 FILLER_3_207 ();
 FILLCELL_X1 FILLER_3_209 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X16 FILLER_4_97 ();
 FILLCELL_X8 FILLER_4_113 ();
 FILLCELL_X2 FILLER_4_121 ();
 FILLCELL_X32 FILLER_4_127 ();
 FILLCELL_X32 FILLER_4_159 ();
 FILLCELL_X16 FILLER_4_191 ();
 FILLCELL_X2 FILLER_4_207 ();
 FILLCELL_X1 FILLER_4_209 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X16 FILLER_5_65 ();
 FILLCELL_X16 FILLER_5_85 ();
 FILLCELL_X8 FILLER_5_101 ();
 FILLCELL_X2 FILLER_5_109 ();
 FILLCELL_X32 FILLER_5_120 ();
 FILLCELL_X32 FILLER_5_152 ();
 FILLCELL_X16 FILLER_5_184 ();
 FILLCELL_X8 FILLER_5_200 ();
 FILLCELL_X2 FILLER_5_208 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X4 FILLER_6_65 ();
 FILLCELL_X2 FILLER_6_69 ();
 FILLCELL_X1 FILLER_6_71 ();
 FILLCELL_X16 FILLER_6_85 ();
 FILLCELL_X4 FILLER_6_101 ();
 FILLCELL_X1 FILLER_6_105 ();
 FILLCELL_X32 FILLER_6_123 ();
 FILLCELL_X32 FILLER_6_155 ();
 FILLCELL_X16 FILLER_6_187 ();
 FILLCELL_X4 FILLER_6_203 ();
 FILLCELL_X2 FILLER_6_207 ();
 FILLCELL_X1 FILLER_6_209 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X4 FILLER_7_65 ();
 FILLCELL_X16 FILLER_7_86 ();
 FILLCELL_X4 FILLER_7_102 ();
 FILLCELL_X2 FILLER_7_106 ();
 FILLCELL_X1 FILLER_7_108 ();
 FILLCELL_X8 FILLER_7_134 ();
 FILLCELL_X2 FILLER_7_142 ();
 FILLCELL_X1 FILLER_7_144 ();
 FILLCELL_X8 FILLER_7_162 ();
 FILLCELL_X4 FILLER_7_170 ();
 FILLCELL_X1 FILLER_7_174 ();
 FILLCELL_X32 FILLER_7_178 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X8 FILLER_8_65 ();
 FILLCELL_X1 FILLER_8_73 ();
 FILLCELL_X16 FILLER_8_85 ();
 FILLCELL_X8 FILLER_8_101 ();
 FILLCELL_X2 FILLER_8_109 ();
 FILLCELL_X32 FILLER_8_133 ();
 FILLCELL_X32 FILLER_8_165 ();
 FILLCELL_X8 FILLER_8_197 ();
 FILLCELL_X4 FILLER_8_205 ();
 FILLCELL_X1 FILLER_8_209 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X2 FILLER_9_97 ();
 FILLCELL_X1 FILLER_9_99 ();
 FILLCELL_X16 FILLER_9_102 ();
 FILLCELL_X32 FILLER_9_124 ();
 FILLCELL_X32 FILLER_9_156 ();
 FILLCELL_X16 FILLER_9_188 ();
 FILLCELL_X4 FILLER_9_204 ();
 FILLCELL_X2 FILLER_9_208 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X8 FILLER_10_65 ();
 FILLCELL_X2 FILLER_10_73 ();
 FILLCELL_X16 FILLER_10_85 ();
 FILLCELL_X8 FILLER_10_101 ();
 FILLCELL_X4 FILLER_10_109 ();
 FILLCELL_X2 FILLER_10_113 ();
 FILLCELL_X32 FILLER_10_120 ();
 FILLCELL_X32 FILLER_10_152 ();
 FILLCELL_X16 FILLER_10_184 ();
 FILLCELL_X8 FILLER_10_200 ();
 FILLCELL_X2 FILLER_10_208 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X8 FILLER_11_65 ();
 FILLCELL_X2 FILLER_11_73 ();
 FILLCELL_X16 FILLER_11_91 ();
 FILLCELL_X4 FILLER_11_107 ();
 FILLCELL_X2 FILLER_11_111 ();
 FILLCELL_X1 FILLER_11_113 ();
 FILLCELL_X1 FILLER_11_123 ();
 FILLCELL_X32 FILLER_11_130 ();
 FILLCELL_X32 FILLER_11_162 ();
 FILLCELL_X16 FILLER_11_194 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_33 ();
 FILLCELL_X8 FILLER_12_49 ();
 FILLCELL_X4 FILLER_12_57 ();
 FILLCELL_X2 FILLER_12_61 ();
 FILLCELL_X1 FILLER_12_63 ();
 FILLCELL_X16 FILLER_12_88 ();
 FILLCELL_X8 FILLER_12_104 ();
 FILLCELL_X8 FILLER_12_114 ();
 FILLCELL_X2 FILLER_12_140 ();
 FILLCELL_X16 FILLER_12_148 ();
 FILLCELL_X4 FILLER_12_164 ();
 FILLCELL_X2 FILLER_12_168 ();
 FILLCELL_X32 FILLER_12_173 ();
 FILLCELL_X4 FILLER_12_205 ();
 FILLCELL_X1 FILLER_12_209 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_17 ();
 FILLCELL_X1 FILLER_13_19 ();
 FILLCELL_X32 FILLER_13_23 ();
 FILLCELL_X16 FILLER_13_55 ();
 FILLCELL_X4 FILLER_13_79 ();
 FILLCELL_X8 FILLER_13_93 ();
 FILLCELL_X4 FILLER_13_101 ();
 FILLCELL_X2 FILLER_13_105 ();
 FILLCELL_X1 FILLER_13_107 ();
 FILLCELL_X2 FILLER_13_123 ();
 FILLCELL_X1 FILLER_13_125 ();
 FILLCELL_X2 FILLER_13_135 ();
 FILLCELL_X16 FILLER_13_140 ();
 FILLCELL_X8 FILLER_13_156 ();
 FILLCELL_X4 FILLER_13_164 ();
 FILLCELL_X2 FILLER_13_168 ();
 FILLCELL_X1 FILLER_13_170 ();
 FILLCELL_X32 FILLER_13_174 ();
 FILLCELL_X4 FILLER_13_206 ();
 FILLCELL_X32 FILLER_14_4 ();
 FILLCELL_X32 FILLER_14_36 ();
 FILLCELL_X4 FILLER_14_90 ();
 FILLCELL_X16 FILLER_14_100 ();
 FILLCELL_X8 FILLER_14_116 ();
 FILLCELL_X4 FILLER_14_124 ();
 FILLCELL_X2 FILLER_14_135 ();
 FILLCELL_X1 FILLER_14_137 ();
 FILLCELL_X2 FILLER_14_145 ();
 FILLCELL_X32 FILLER_14_164 ();
 FILLCELL_X8 FILLER_14_196 ();
 FILLCELL_X4 FILLER_14_204 ();
 FILLCELL_X2 FILLER_14_208 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X8 FILLER_15_65 ();
 FILLCELL_X2 FILLER_15_73 ();
 FILLCELL_X1 FILLER_15_75 ();
 FILLCELL_X8 FILLER_15_79 ();
 FILLCELL_X4 FILLER_15_87 ();
 FILLCELL_X2 FILLER_15_91 ();
 FILLCELL_X1 FILLER_15_93 ();
 FILLCELL_X8 FILLER_15_107 ();
 FILLCELL_X1 FILLER_15_115 ();
 FILLCELL_X4 FILLER_15_121 ();
 FILLCELL_X2 FILLER_15_125 ();
 FILLCELL_X1 FILLER_15_127 ();
 FILLCELL_X32 FILLER_15_151 ();
 FILLCELL_X16 FILLER_15_183 ();
 FILLCELL_X8 FILLER_15_199 ();
 FILLCELL_X2 FILLER_15_207 ();
 FILLCELL_X1 FILLER_15_209 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X8 FILLER_16_17 ();
 FILLCELL_X32 FILLER_16_28 ();
 FILLCELL_X4 FILLER_16_60 ();
 FILLCELL_X1 FILLER_16_64 ();
 FILLCELL_X8 FILLER_16_82 ();
 FILLCELL_X4 FILLER_16_90 ();
 FILLCELL_X2 FILLER_16_101 ();
 FILLCELL_X8 FILLER_16_106 ();
 FILLCELL_X4 FILLER_16_114 ();
 FILLCELL_X2 FILLER_16_118 ();
 FILLCELL_X1 FILLER_16_120 ();
 FILLCELL_X1 FILLER_16_132 ();
 FILLCELL_X2 FILLER_16_137 ();
 FILLCELL_X4 FILLER_16_143 ();
 FILLCELL_X32 FILLER_16_150 ();
 FILLCELL_X16 FILLER_16_182 ();
 FILLCELL_X8 FILLER_16_198 ();
 FILLCELL_X4 FILLER_16_206 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X4 FILLER_17_65 ();
 FILLCELL_X2 FILLER_17_69 ();
 FILLCELL_X1 FILLER_17_71 ();
 FILLCELL_X16 FILLER_17_106 ();
 FILLCELL_X8 FILLER_17_122 ();
 FILLCELL_X1 FILLER_17_130 ();
 FILLCELL_X16 FILLER_17_134 ();
 FILLCELL_X1 FILLER_17_150 ();
 FILLCELL_X2 FILLER_17_168 ();
 FILLCELL_X1 FILLER_17_170 ();
 FILLCELL_X32 FILLER_17_174 ();
 FILLCELL_X4 FILLER_17_206 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X16 FILLER_18_65 ();
 FILLCELL_X4 FILLER_18_81 ();
 FILLCELL_X2 FILLER_18_85 ();
 FILLCELL_X1 FILLER_18_87 ();
 FILLCELL_X2 FILLER_18_90 ();
 FILLCELL_X1 FILLER_18_96 ();
 FILLCELL_X32 FILLER_18_114 ();
 FILLCELL_X32 FILLER_18_146 ();
 FILLCELL_X32 FILLER_18_178 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X16 FILLER_19_124 ();
 FILLCELL_X1 FILLER_19_140 ();
 FILLCELL_X32 FILLER_19_148 ();
 FILLCELL_X16 FILLER_19_180 ();
 FILLCELL_X8 FILLER_19_196 ();
 FILLCELL_X4 FILLER_19_204 ();
 FILLCELL_X2 FILLER_19_208 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X16 FILLER_20_65 ();
 FILLCELL_X4 FILLER_20_81 ();
 FILLCELL_X2 FILLER_20_85 ();
 FILLCELL_X8 FILLER_20_90 ();
 FILLCELL_X2 FILLER_20_98 ();
 FILLCELL_X32 FILLER_20_103 ();
 FILLCELL_X32 FILLER_20_135 ();
 FILLCELL_X32 FILLER_20_167 ();
 FILLCELL_X8 FILLER_20_199 ();
 FILLCELL_X2 FILLER_20_207 ();
 FILLCELL_X1 FILLER_20_209 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X16 FILLER_21_193 ();
 FILLCELL_X1 FILLER_21_209 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X16 FILLER_22_193 ();
 FILLCELL_X1 FILLER_22_209 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X16 FILLER_23_193 ();
 FILLCELL_X1 FILLER_23_209 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X2 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_148 ();
 FILLCELL_X16 FILLER_24_180 ();
 FILLCELL_X8 FILLER_24_196 ();
 FILLCELL_X4 FILLER_24_204 ();
 FILLCELL_X2 FILLER_24_208 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X16 FILLER_25_65 ();
 FILLCELL_X1 FILLER_25_81 ();
 FILLCELL_X32 FILLER_25_116 ();
 FILLCELL_X32 FILLER_25_148 ();
 FILLCELL_X16 FILLER_25_180 ();
 FILLCELL_X8 FILLER_25_196 ();
 FILLCELL_X4 FILLER_25_204 ();
 FILLCELL_X2 FILLER_25_208 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X4 FILLER_26_97 ();
 FILLCELL_X1 FILLER_26_101 ();
 FILLCELL_X32 FILLER_26_105 ();
 FILLCELL_X8 FILLER_26_137 ();
 FILLCELL_X2 FILLER_26_145 ();
 FILLCELL_X1 FILLER_26_147 ();
 FILLCELL_X32 FILLER_26_151 ();
 FILLCELL_X16 FILLER_26_183 ();
 FILLCELL_X8 FILLER_26_199 ();
 FILLCELL_X2 FILLER_26_207 ();
 FILLCELL_X1 FILLER_26_209 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X8 FILLER_27_65 ();
 FILLCELL_X4 FILLER_27_73 ();
 FILLCELL_X2 FILLER_27_77 ();
 FILLCELL_X1 FILLER_27_79 ();
 FILLCELL_X32 FILLER_27_83 ();
 FILLCELL_X32 FILLER_27_118 ();
 FILLCELL_X32 FILLER_27_150 ();
 FILLCELL_X16 FILLER_27_182 ();
 FILLCELL_X8 FILLER_27_198 ();
 FILLCELL_X4 FILLER_27_206 ();
endmodule
