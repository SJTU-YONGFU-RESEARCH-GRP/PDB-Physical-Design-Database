module bidirectional_fifo (a_almost_empty,
    a_almost_full,
    a_empty,
    a_full,
    a_rd_en,
    a_wr_en,
    b_almost_empty,
    b_almost_full,
    b_empty,
    b_full,
    b_rd_en,
    b_wr_en,
    clk,
    rst_n,
    a_rd_data,
    a_to_b_count,
    a_wr_data,
    b_rd_data,
    b_to_a_count,
    b_wr_data);
 output a_almost_empty;
 output a_almost_full;
 output a_empty;
 output a_full;
 input a_rd_en;
 input a_wr_en;
 output b_almost_empty;
 output b_almost_full;
 output b_empty;
 output b_full;
 input b_rd_en;
 input b_wr_en;
 input clk;
 input rst_n;
 output [7:0] a_rd_data;
 output [4:0] a_to_b_count;
 input [7:0] a_wr_data;
 output [7:0] b_rd_data;
 output [4:0] b_to_a_count;
 input [7:0] b_wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire \a_rd_ptr[0] ;
 wire \a_rd_ptr[1] ;
 wire \a_rd_ptr[2] ;
 wire \a_rd_ptr[3] ;
 wire \a_rd_ptr[4] ;
 wire \a_to_b_mem[0][0] ;
 wire \a_to_b_mem[0][1] ;
 wire \a_to_b_mem[0][2] ;
 wire \a_to_b_mem[0][3] ;
 wire \a_to_b_mem[0][4] ;
 wire \a_to_b_mem[0][5] ;
 wire \a_to_b_mem[0][6] ;
 wire \a_to_b_mem[0][7] ;
 wire \a_to_b_mem[10][0] ;
 wire \a_to_b_mem[10][1] ;
 wire \a_to_b_mem[10][2] ;
 wire \a_to_b_mem[10][3] ;
 wire \a_to_b_mem[10][4] ;
 wire \a_to_b_mem[10][5] ;
 wire \a_to_b_mem[10][6] ;
 wire \a_to_b_mem[10][7] ;
 wire \a_to_b_mem[11][0] ;
 wire \a_to_b_mem[11][1] ;
 wire \a_to_b_mem[11][2] ;
 wire \a_to_b_mem[11][3] ;
 wire \a_to_b_mem[11][4] ;
 wire \a_to_b_mem[11][5] ;
 wire \a_to_b_mem[11][6] ;
 wire \a_to_b_mem[11][7] ;
 wire \a_to_b_mem[12][0] ;
 wire \a_to_b_mem[12][1] ;
 wire \a_to_b_mem[12][2] ;
 wire \a_to_b_mem[12][3] ;
 wire \a_to_b_mem[12][4] ;
 wire \a_to_b_mem[12][5] ;
 wire \a_to_b_mem[12][6] ;
 wire \a_to_b_mem[12][7] ;
 wire \a_to_b_mem[13][0] ;
 wire \a_to_b_mem[13][1] ;
 wire \a_to_b_mem[13][2] ;
 wire \a_to_b_mem[13][3] ;
 wire \a_to_b_mem[13][4] ;
 wire \a_to_b_mem[13][5] ;
 wire \a_to_b_mem[13][6] ;
 wire \a_to_b_mem[13][7] ;
 wire \a_to_b_mem[14][0] ;
 wire \a_to_b_mem[14][1] ;
 wire \a_to_b_mem[14][2] ;
 wire \a_to_b_mem[14][3] ;
 wire \a_to_b_mem[14][4] ;
 wire \a_to_b_mem[14][5] ;
 wire \a_to_b_mem[14][6] ;
 wire \a_to_b_mem[14][7] ;
 wire \a_to_b_mem[15][0] ;
 wire \a_to_b_mem[15][1] ;
 wire \a_to_b_mem[15][2] ;
 wire \a_to_b_mem[15][3] ;
 wire \a_to_b_mem[15][4] ;
 wire \a_to_b_mem[15][5] ;
 wire \a_to_b_mem[15][6] ;
 wire \a_to_b_mem[15][7] ;
 wire \a_to_b_mem[1][0] ;
 wire \a_to_b_mem[1][1] ;
 wire \a_to_b_mem[1][2] ;
 wire \a_to_b_mem[1][3] ;
 wire \a_to_b_mem[1][4] ;
 wire \a_to_b_mem[1][5] ;
 wire \a_to_b_mem[1][6] ;
 wire \a_to_b_mem[1][7] ;
 wire \a_to_b_mem[2][0] ;
 wire \a_to_b_mem[2][1] ;
 wire \a_to_b_mem[2][2] ;
 wire \a_to_b_mem[2][3] ;
 wire \a_to_b_mem[2][4] ;
 wire \a_to_b_mem[2][5] ;
 wire \a_to_b_mem[2][6] ;
 wire \a_to_b_mem[2][7] ;
 wire \a_to_b_mem[3][0] ;
 wire \a_to_b_mem[3][1] ;
 wire \a_to_b_mem[3][2] ;
 wire \a_to_b_mem[3][3] ;
 wire \a_to_b_mem[3][4] ;
 wire \a_to_b_mem[3][5] ;
 wire \a_to_b_mem[3][6] ;
 wire \a_to_b_mem[3][7] ;
 wire \a_to_b_mem[4][0] ;
 wire \a_to_b_mem[4][1] ;
 wire \a_to_b_mem[4][2] ;
 wire \a_to_b_mem[4][3] ;
 wire \a_to_b_mem[4][4] ;
 wire \a_to_b_mem[4][5] ;
 wire \a_to_b_mem[4][6] ;
 wire \a_to_b_mem[4][7] ;
 wire \a_to_b_mem[5][0] ;
 wire \a_to_b_mem[5][1] ;
 wire \a_to_b_mem[5][2] ;
 wire \a_to_b_mem[5][3] ;
 wire \a_to_b_mem[5][4] ;
 wire \a_to_b_mem[5][5] ;
 wire \a_to_b_mem[5][6] ;
 wire \a_to_b_mem[5][7] ;
 wire \a_to_b_mem[6][0] ;
 wire \a_to_b_mem[6][1] ;
 wire \a_to_b_mem[6][2] ;
 wire \a_to_b_mem[6][3] ;
 wire \a_to_b_mem[6][4] ;
 wire \a_to_b_mem[6][5] ;
 wire \a_to_b_mem[6][6] ;
 wire \a_to_b_mem[6][7] ;
 wire \a_to_b_mem[7][0] ;
 wire \a_to_b_mem[7][1] ;
 wire \a_to_b_mem[7][2] ;
 wire \a_to_b_mem[7][3] ;
 wire \a_to_b_mem[7][4] ;
 wire \a_to_b_mem[7][5] ;
 wire \a_to_b_mem[7][6] ;
 wire \a_to_b_mem[7][7] ;
 wire \a_to_b_mem[8][0] ;
 wire \a_to_b_mem[8][1] ;
 wire \a_to_b_mem[8][2] ;
 wire \a_to_b_mem[8][3] ;
 wire \a_to_b_mem[8][4] ;
 wire \a_to_b_mem[8][5] ;
 wire \a_to_b_mem[8][6] ;
 wire \a_to_b_mem[8][7] ;
 wire \a_to_b_mem[9][0] ;
 wire \a_to_b_mem[9][1] ;
 wire \a_to_b_mem[9][2] ;
 wire \a_to_b_mem[9][3] ;
 wire \a_to_b_mem[9][4] ;
 wire \a_to_b_mem[9][5] ;
 wire \a_to_b_mem[9][6] ;
 wire \a_to_b_mem[9][7] ;
 wire \a_wr_ptr[0] ;
 wire \a_wr_ptr[1] ;
 wire \a_wr_ptr[2] ;
 wire \a_wr_ptr[3] ;
 wire \a_wr_ptr[4] ;
 wire \b_rd_ptr[0] ;
 wire \b_rd_ptr[1] ;
 wire \b_rd_ptr[2] ;
 wire \b_rd_ptr[3] ;
 wire \b_rd_ptr[4] ;
 wire \b_to_a_mem[0][0] ;
 wire \b_to_a_mem[0][1] ;
 wire \b_to_a_mem[0][2] ;
 wire \b_to_a_mem[0][3] ;
 wire \b_to_a_mem[0][4] ;
 wire \b_to_a_mem[0][5] ;
 wire \b_to_a_mem[0][6] ;
 wire \b_to_a_mem[0][7] ;
 wire \b_to_a_mem[10][0] ;
 wire \b_to_a_mem[10][1] ;
 wire \b_to_a_mem[10][2] ;
 wire \b_to_a_mem[10][3] ;
 wire \b_to_a_mem[10][4] ;
 wire \b_to_a_mem[10][5] ;
 wire \b_to_a_mem[10][6] ;
 wire \b_to_a_mem[10][7] ;
 wire \b_to_a_mem[11][0] ;
 wire \b_to_a_mem[11][1] ;
 wire \b_to_a_mem[11][2] ;
 wire \b_to_a_mem[11][3] ;
 wire \b_to_a_mem[11][4] ;
 wire \b_to_a_mem[11][5] ;
 wire \b_to_a_mem[11][6] ;
 wire \b_to_a_mem[11][7] ;
 wire \b_to_a_mem[12][0] ;
 wire \b_to_a_mem[12][1] ;
 wire \b_to_a_mem[12][2] ;
 wire \b_to_a_mem[12][3] ;
 wire \b_to_a_mem[12][4] ;
 wire \b_to_a_mem[12][5] ;
 wire \b_to_a_mem[12][6] ;
 wire \b_to_a_mem[12][7] ;
 wire \b_to_a_mem[13][0] ;
 wire \b_to_a_mem[13][1] ;
 wire \b_to_a_mem[13][2] ;
 wire \b_to_a_mem[13][3] ;
 wire \b_to_a_mem[13][4] ;
 wire \b_to_a_mem[13][5] ;
 wire \b_to_a_mem[13][6] ;
 wire \b_to_a_mem[13][7] ;
 wire \b_to_a_mem[14][0] ;
 wire \b_to_a_mem[14][1] ;
 wire \b_to_a_mem[14][2] ;
 wire \b_to_a_mem[14][3] ;
 wire \b_to_a_mem[14][4] ;
 wire \b_to_a_mem[14][5] ;
 wire \b_to_a_mem[14][6] ;
 wire \b_to_a_mem[14][7] ;
 wire \b_to_a_mem[15][0] ;
 wire \b_to_a_mem[15][1] ;
 wire \b_to_a_mem[15][2] ;
 wire \b_to_a_mem[15][3] ;
 wire \b_to_a_mem[15][4] ;
 wire \b_to_a_mem[15][5] ;
 wire \b_to_a_mem[15][6] ;
 wire \b_to_a_mem[15][7] ;
 wire \b_to_a_mem[1][0] ;
 wire \b_to_a_mem[1][1] ;
 wire \b_to_a_mem[1][2] ;
 wire \b_to_a_mem[1][3] ;
 wire \b_to_a_mem[1][4] ;
 wire \b_to_a_mem[1][5] ;
 wire \b_to_a_mem[1][6] ;
 wire \b_to_a_mem[1][7] ;
 wire \b_to_a_mem[2][0] ;
 wire \b_to_a_mem[2][1] ;
 wire \b_to_a_mem[2][2] ;
 wire \b_to_a_mem[2][3] ;
 wire \b_to_a_mem[2][4] ;
 wire \b_to_a_mem[2][5] ;
 wire \b_to_a_mem[2][6] ;
 wire \b_to_a_mem[2][7] ;
 wire \b_to_a_mem[3][0] ;
 wire \b_to_a_mem[3][1] ;
 wire \b_to_a_mem[3][2] ;
 wire \b_to_a_mem[3][3] ;
 wire \b_to_a_mem[3][4] ;
 wire \b_to_a_mem[3][5] ;
 wire \b_to_a_mem[3][6] ;
 wire \b_to_a_mem[3][7] ;
 wire \b_to_a_mem[4][0] ;
 wire \b_to_a_mem[4][1] ;
 wire \b_to_a_mem[4][2] ;
 wire \b_to_a_mem[4][3] ;
 wire \b_to_a_mem[4][4] ;
 wire \b_to_a_mem[4][5] ;
 wire \b_to_a_mem[4][6] ;
 wire \b_to_a_mem[4][7] ;
 wire \b_to_a_mem[5][0] ;
 wire \b_to_a_mem[5][1] ;
 wire \b_to_a_mem[5][2] ;
 wire \b_to_a_mem[5][3] ;
 wire \b_to_a_mem[5][4] ;
 wire \b_to_a_mem[5][5] ;
 wire \b_to_a_mem[5][6] ;
 wire \b_to_a_mem[5][7] ;
 wire \b_to_a_mem[6][0] ;
 wire \b_to_a_mem[6][1] ;
 wire \b_to_a_mem[6][2] ;
 wire \b_to_a_mem[6][3] ;
 wire \b_to_a_mem[6][4] ;
 wire \b_to_a_mem[6][5] ;
 wire \b_to_a_mem[6][6] ;
 wire \b_to_a_mem[6][7] ;
 wire \b_to_a_mem[7][0] ;
 wire \b_to_a_mem[7][1] ;
 wire \b_to_a_mem[7][2] ;
 wire \b_to_a_mem[7][3] ;
 wire \b_to_a_mem[7][4] ;
 wire \b_to_a_mem[7][5] ;
 wire \b_to_a_mem[7][6] ;
 wire \b_to_a_mem[7][7] ;
 wire \b_to_a_mem[8][0] ;
 wire \b_to_a_mem[8][1] ;
 wire \b_to_a_mem[8][2] ;
 wire \b_to_a_mem[8][3] ;
 wire \b_to_a_mem[8][4] ;
 wire \b_to_a_mem[8][5] ;
 wire \b_to_a_mem[8][6] ;
 wire \b_to_a_mem[8][7] ;
 wire \b_to_a_mem[9][0] ;
 wire \b_to_a_mem[9][1] ;
 wire \b_to_a_mem[9][2] ;
 wire \b_to_a_mem[9][3] ;
 wire \b_to_a_mem[9][4] ;
 wire \b_to_a_mem[9][5] ;
 wire \b_to_a_mem[9][6] ;
 wire \b_to_a_mem[9][7] ;
 wire \b_wr_ptr[0] ;
 wire \b_wr_ptr[1] ;
 wire \b_wr_ptr[2] ;
 wire \b_wr_ptr[3] ;
 wire \b_wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;

 sky130_fd_sc_hd__inv_1 _316_ (.A(_315_),
    .Y(net51));
 sky130_fd_sc_hd__xor2_2 _317_ (.A(_290_),
    .B(_274_),
    .X(net53));
 sky130_fd_sc_hd__inv_1 _318_ (.A(_280_),
    .Y(_074_));
 sky130_fd_sc_hd__nand2_1 _319_ (.A(_290_),
    .B(_282_),
    .Y(_075_));
 sky130_fd_sc_hd__a21oi_1 _320_ (.A1(_290_),
    .A2(_281_),
    .B1(_289_),
    .Y(_076_));
 sky130_fd_sc_hd__o21ai_4 _321_ (.A1(_314_),
    .A2(_075_),
    .B1(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__xnor2_1 _322_ (.A(_074_),
    .B(_077_),
    .Y(net54));
 sky130_fd_sc_hd__a21o_1 _323_ (.A1(_290_),
    .A2(_274_),
    .B1(_289_),
    .X(_078_));
 sky130_fd_sc_hd__a21oi_2 _324_ (.A1(_280_),
    .A2(_078_),
    .B1(_279_),
    .Y(_079_));
 sky130_fd_sc_hd__xnor2_2 _325_ (.A(\b_wr_ptr[4] ),
    .B(\a_rd_ptr[4] ),
    .Y(_080_));
 sky130_fd_sc_hd__xnor2_4 _326_ (.A(_079_),
    .B(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__clkbuf_4 _327_ (.A(_081_),
    .X(net55));
 sky130_fd_sc_hd__inv_1 _328_ (.A(_313_),
    .Y(net34));
 sky130_fd_sc_hd__inv_1 _329_ (.A(_285_),
    .Y(_082_));
 sky130_fd_sc_hd__nand2_1 _330_ (.A(_293_),
    .B(_287_),
    .Y(_083_));
 sky130_fd_sc_hd__a21oi_1 _331_ (.A1(_293_),
    .A2(_286_),
    .B1(_292_),
    .Y(_084_));
 sky130_fd_sc_hd__o21ai_4 _332_ (.A1(_312_),
    .A2(_083_),
    .B1(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__xnor2_1 _333_ (.A(_082_),
    .B(_085_),
    .Y(net37));
 sky130_fd_sc_hd__xor2_4 _334_ (.A(_293_),
    .B(_277_),
    .X(net36));
 sky130_fd_sc_hd__a21o_1 _335_ (.A1(_293_),
    .A2(_277_),
    .B1(_292_),
    .X(_086_));
 sky130_fd_sc_hd__a21oi_2 _336_ (.A1(_285_),
    .A2(_086_),
    .B1(_284_),
    .Y(_087_));
 sky130_fd_sc_hd__xnor2_2 _337_ (.A(\a_wr_ptr[4] ),
    .B(\b_rd_ptr[4] ),
    .Y(_088_));
 sky130_fd_sc_hd__xnor2_4 _338_ (.A(_087_),
    .B(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__buf_4 _339_ (.A(_089_),
    .X(net38));
 sky130_fd_sc_hd__nor4_2 _340_ (.A(_285_),
    .B(net34),
    .C(net35),
    .D(net36),
    .Y(_090_));
 sky130_fd_sc_hd__nor4_2 _341_ (.A(_082_),
    .B(net34),
    .C(net35),
    .D(net36),
    .Y(_091_));
 sky130_fd_sc_hd__mux2_4 _342_ (.A0(_090_),
    .A1(_091_),
    .S(_085_),
    .X(_092_));
 sky130_fd_sc_hd__and2_0 _343_ (.A(net38),
    .B(_092_),
    .X(net42));
 sky130_fd_sc_hd__nor4_1 _344_ (.A(_280_),
    .B(net51),
    .C(net52),
    .D(net53),
    .Y(_093_));
 sky130_fd_sc_hd__nor4_1 _345_ (.A(_074_),
    .B(net51),
    .C(net52),
    .D(net53),
    .Y(_094_));
 sky130_fd_sc_hd__mux2_2 _346_ (.A0(_093_),
    .A1(_094_),
    .S(_077_),
    .X(_095_));
 sky130_fd_sc_hd__and2_0 _347_ (.A(net55),
    .B(_095_),
    .X(net25));
 sky130_fd_sc_hd__mux2i_4 _348_ (.A0(_093_),
    .A1(_094_),
    .S(_077_),
    .Y(_096_));
 sky130_fd_sc_hd__nor2_1 _349_ (.A(net55),
    .B(_096_),
    .Y(net24));
 sky130_fd_sc_hd__mux2i_4 _350_ (.A0(_090_),
    .A1(_091_),
    .S(_085_),
    .Y(_097_));
 sky130_fd_sc_hd__nor2_1 _351_ (.A(net38),
    .B(_097_),
    .Y(net41));
 sky130_fd_sc_hd__nor2_1 _352_ (.A(\a_wr_ptr[3] ),
    .B(\a_wr_ptr[2] ),
    .Y(_098_));
 sky130_fd_sc_hd__a21boi_2 _353_ (.A1(_089_),
    .A2(_092_),
    .B1_N(net11),
    .Y(_099_));
 sky130_fd_sc_hd__and3_4 _354_ (.A(_305_),
    .B(_098_),
    .C(_099_),
    .X(_000_));
 sky130_fd_sc_hd__and3_4 _355_ (.A(_308_),
    .B(_098_),
    .C(_099_),
    .X(_007_));
 sky130_fd_sc_hd__and3_4 _356_ (.A(_306_),
    .B(_098_),
    .C(_099_),
    .X(_008_));
 sky130_fd_sc_hd__nand2_1 _357_ (.A(net11),
    .B(_310_),
    .Y(_100_));
 sky130_fd_sc_hd__a21oi_2 _358_ (.A1(_089_),
    .A2(_092_),
    .B1(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__and2_4 _359_ (.A(_098_),
    .B(_101_),
    .X(_009_));
 sky130_fd_sc_hd__buf_4 _360_ (.A(_099_),
    .X(_102_));
 sky130_fd_sc_hd__nor2b_1 _361_ (.A(\a_wr_ptr[3] ),
    .B_N(\a_wr_ptr[2] ),
    .Y(_103_));
 sky130_fd_sc_hd__and3_4 _362_ (.A(_305_),
    .B(_102_),
    .C(_103_),
    .X(_010_));
 sky130_fd_sc_hd__and3_4 _363_ (.A(_308_),
    .B(_102_),
    .C(_103_),
    .X(_011_));
 sky130_fd_sc_hd__and3_4 _364_ (.A(_306_),
    .B(_102_),
    .C(_103_),
    .X(_012_));
 sky130_fd_sc_hd__and2_4 _365_ (.A(_101_),
    .B(_103_),
    .X(_013_));
 sky130_fd_sc_hd__nor2b_1 _366_ (.A(\a_wr_ptr[2] ),
    .B_N(\a_wr_ptr[3] ),
    .Y(_104_));
 sky130_fd_sc_hd__and3_4 _367_ (.A(_305_),
    .B(_102_),
    .C(_104_),
    .X(_014_));
 sky130_fd_sc_hd__and3_4 _368_ (.A(_308_),
    .B(_102_),
    .C(_104_),
    .X(_015_));
 sky130_fd_sc_hd__and3_4 _369_ (.A(_306_),
    .B(_102_),
    .C(_104_),
    .X(_001_));
 sky130_fd_sc_hd__and2_4 _370_ (.A(_101_),
    .B(_104_),
    .X(_002_));
 sky130_fd_sc_hd__and2_0 _371_ (.A(\a_wr_ptr[3] ),
    .B(\a_wr_ptr[2] ),
    .X(_105_));
 sky130_fd_sc_hd__and3_4 _372_ (.A(_305_),
    .B(_102_),
    .C(_105_),
    .X(_003_));
 sky130_fd_sc_hd__and3_4 _373_ (.A(_308_),
    .B(_102_),
    .C(_105_),
    .X(_004_));
 sky130_fd_sc_hd__and3_4 _374_ (.A(_306_),
    .B(_102_),
    .C(_105_),
    .X(_005_));
 sky130_fd_sc_hd__nand3_1 _375_ (.A(net11),
    .B(_310_),
    .C(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__a21oi_4 _376_ (.A1(net38),
    .A2(_092_),
    .B1(_106_),
    .Y(_006_));
 sky130_fd_sc_hd__nor2_1 _377_ (.A(\b_wr_ptr[3] ),
    .B(\b_wr_ptr[2] ),
    .Y(_107_));
 sky130_fd_sc_hd__a21boi_2 _378_ (.A1(_081_),
    .A2(_095_),
    .B1_N(net21),
    .Y(_108_));
 sky130_fd_sc_hd__and3_4 _379_ (.A(_296_),
    .B(_107_),
    .C(_108_),
    .X(_016_));
 sky130_fd_sc_hd__and3_4 _380_ (.A(_299_),
    .B(_107_),
    .C(_108_),
    .X(_023_));
 sky130_fd_sc_hd__and3_4 _381_ (.A(_297_),
    .B(_107_),
    .C(_108_),
    .X(_024_));
 sky130_fd_sc_hd__nand2_1 _382_ (.A(net21),
    .B(_301_),
    .Y(_109_));
 sky130_fd_sc_hd__a21oi_2 _383_ (.A1(_081_),
    .A2(_095_),
    .B1(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__and2_4 _384_ (.A(_107_),
    .B(_110_),
    .X(_025_));
 sky130_fd_sc_hd__buf_4 _385_ (.A(_108_),
    .X(_111_));
 sky130_fd_sc_hd__nor2b_1 _386_ (.A(\b_wr_ptr[3] ),
    .B_N(\b_wr_ptr[2] ),
    .Y(_112_));
 sky130_fd_sc_hd__and3_4 _387_ (.A(_296_),
    .B(_111_),
    .C(_112_),
    .X(_026_));
 sky130_fd_sc_hd__and3_4 _388_ (.A(_299_),
    .B(_111_),
    .C(_112_),
    .X(_027_));
 sky130_fd_sc_hd__and3_4 _389_ (.A(_297_),
    .B(_111_),
    .C(_112_),
    .X(_028_));
 sky130_fd_sc_hd__and2_4 _390_ (.A(_110_),
    .B(_112_),
    .X(_029_));
 sky130_fd_sc_hd__nor2b_1 _391_ (.A(\b_wr_ptr[2] ),
    .B_N(\b_wr_ptr[3] ),
    .Y(_113_));
 sky130_fd_sc_hd__and3_4 _392_ (.A(_296_),
    .B(_111_),
    .C(_113_),
    .X(_030_));
 sky130_fd_sc_hd__and3_4 _393_ (.A(_299_),
    .B(_111_),
    .C(_113_),
    .X(_031_));
 sky130_fd_sc_hd__and3_4 _394_ (.A(_297_),
    .B(_111_),
    .C(_113_),
    .X(_017_));
 sky130_fd_sc_hd__and2_4 _395_ (.A(_110_),
    .B(_113_),
    .X(_018_));
 sky130_fd_sc_hd__and2_0 _396_ (.A(\b_wr_ptr[3] ),
    .B(\b_wr_ptr[2] ),
    .X(_114_));
 sky130_fd_sc_hd__and3_4 _397_ (.A(_296_),
    .B(_111_),
    .C(_114_),
    .X(_019_));
 sky130_fd_sc_hd__and3_4 _398_ (.A(_299_),
    .B(_111_),
    .C(_114_),
    .X(_020_));
 sky130_fd_sc_hd__and3_4 _399_ (.A(_297_),
    .B(_111_),
    .C(_114_),
    .X(_021_));
 sky130_fd_sc_hd__nand3_1 _400_ (.A(net21),
    .B(_301_),
    .C(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__a21oi_4 _401_ (.A1(net55),
    .A2(_095_),
    .B1(_115_),
    .Y(_022_));
 sky130_fd_sc_hd__clkinvlp_4 _402_ (.A(\a_rd_ptr[3] ),
    .Y(_278_));
 sky130_fd_sc_hd__buf_4 _403_ (.A(\a_rd_ptr[1] ),
    .X(_116_));
 sky130_fd_sc_hd__clkinvlp_4 _404_ (.A(_116_),
    .Y(_272_));
 sky130_fd_sc_hd__inv_1 _405_ (.A(_314_),
    .Y(_273_));
 sky130_fd_sc_hd__buf_4 _406_ (.A(\a_rd_ptr[2] ),
    .X(_117_));
 sky130_fd_sc_hd__inv_1 _407_ (.A(_117_),
    .Y(_288_));
 sky130_fd_sc_hd__inv_1 _408_ (.A(_312_),
    .Y(_276_));
 sky130_fd_sc_hd__inv_1 _409_ (.A(\b_wr_ptr[0] ),
    .Y(_035_));
 sky130_fd_sc_hd__inv_1 _410_ (.A(\a_wr_ptr[0] ),
    .Y(_032_));
 sky130_fd_sc_hd__clkinvlp_4 _411_ (.A(\b_rd_ptr[3] ),
    .Y(_283_));
 sky130_fd_sc_hd__buf_4 _412_ (.A(\b_rd_ptr[1] ),
    .X(_118_));
 sky130_fd_sc_hd__clkinvlp_4 _413_ (.A(_118_),
    .Y(_275_));
 sky130_fd_sc_hd__buf_6 _414_ (.A(\b_rd_ptr[2] ),
    .X(_119_));
 sky130_fd_sc_hd__clkinvlp_4 _415_ (.A(_119_),
    .Y(_291_));
 sky130_fd_sc_hd__inv_1 _416_ (.A(\b_wr_ptr[1] ),
    .Y(_295_));
 sky130_fd_sc_hd__inv_1 _417_ (.A(\a_wr_ptr[1] ),
    .Y(_304_));
 sky130_fd_sc_hd__clkbuf_4 _418_ (.A(\a_rd_ptr[0] ),
    .X(_120_));
 sky130_fd_sc_hd__clkbuf_4 _419_ (.A(\a_rd_ptr[2] ),
    .X(_121_));
 sky130_fd_sc_hd__mux4_1 _420_ (.A0(\b_to_a_mem[0][0] ),
    .A1(\b_to_a_mem[1][0] ),
    .A2(\b_to_a_mem[4][0] ),
    .A3(\b_to_a_mem[5][0] ),
    .S0(_120_),
    .S1(_121_),
    .X(_122_));
 sky130_fd_sc_hd__nand2_4 _421_ (.A(_272_),
    .B(_278_),
    .Y(_123_));
 sky130_fd_sc_hd__buf_4 _422_ (.A(_116_),
    .X(_124_));
 sky130_fd_sc_hd__nand2_4 _423_ (.A(_124_),
    .B(_278_),
    .Y(_125_));
 sky130_fd_sc_hd__buf_4 _424_ (.A(_120_),
    .X(_126_));
 sky130_fd_sc_hd__mux4_1 _425_ (.A0(\b_to_a_mem[2][0] ),
    .A1(\b_to_a_mem[3][0] ),
    .A2(\b_to_a_mem[6][0] ),
    .A3(\b_to_a_mem[7][0] ),
    .S0(_126_),
    .S1(_117_),
    .X(_127_));
 sky130_fd_sc_hd__o22ai_1 _426_ (.A1(_122_),
    .A2(_123_),
    .B1(_125_),
    .B2(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__mux4_1 _427_ (.A0(\b_to_a_mem[8][0] ),
    .A1(\b_to_a_mem[9][0] ),
    .A2(\b_to_a_mem[10][0] ),
    .A3(\b_to_a_mem[11][0] ),
    .S0(_120_),
    .S1(_116_),
    .X(_129_));
 sky130_fd_sc_hd__nand2_4 _428_ (.A(_288_),
    .B(\a_rd_ptr[3] ),
    .Y(_130_));
 sky130_fd_sc_hd__nand2_4 _429_ (.A(_117_),
    .B(\a_rd_ptr[3] ),
    .Y(_131_));
 sky130_fd_sc_hd__mux4_1 _430_ (.A0(\b_to_a_mem[12][0] ),
    .A1(\b_to_a_mem[13][0] ),
    .A2(\b_to_a_mem[14][0] ),
    .A3(\b_to_a_mem[15][0] ),
    .S0(_126_),
    .S1(_124_),
    .X(_132_));
 sky130_fd_sc_hd__o22ai_1 _431_ (.A1(_129_),
    .A2(_130_),
    .B1(_131_),
    .B2(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__nor2_1 _432_ (.A(_128_),
    .B(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__o21ai_4 _433_ (.A1(_081_),
    .A2(_096_),
    .B1(net2),
    .Y(_135_));
 sky130_fd_sc_hd__mux2_1 _434_ (.A0(_134_),
    .A1(net26),
    .S(_135_),
    .X(_038_));
 sky130_fd_sc_hd__buf_4 _435_ (.A(_120_),
    .X(_136_));
 sky130_fd_sc_hd__mux4_1 _436_ (.A0(\b_to_a_mem[2][1] ),
    .A1(\b_to_a_mem[3][1] ),
    .A2(\b_to_a_mem[6][1] ),
    .A3(\b_to_a_mem[7][1] ),
    .S0(_136_),
    .S1(_121_),
    .X(_137_));
 sky130_fd_sc_hd__clkbuf_8 _437_ (.A(_120_),
    .X(_138_));
 sky130_fd_sc_hd__mux4_1 _438_ (.A0(\b_to_a_mem[0][1] ),
    .A1(\b_to_a_mem[1][1] ),
    .A2(\b_to_a_mem[4][1] ),
    .A3(\b_to_a_mem[5][1] ),
    .S0(_138_),
    .S1(_117_),
    .X(_139_));
 sky130_fd_sc_hd__o22ai_1 _439_ (.A1(_125_),
    .A2(_137_),
    .B1(_139_),
    .B2(_123_),
    .Y(_140_));
 sky130_fd_sc_hd__mux4_1 _440_ (.A0(\b_to_a_mem[12][1] ),
    .A1(\b_to_a_mem[13][1] ),
    .A2(\b_to_a_mem[14][1] ),
    .A3(\b_to_a_mem[15][1] ),
    .S0(_138_),
    .S1(_116_),
    .X(_141_));
 sky130_fd_sc_hd__mux4_1 _441_ (.A0(\b_to_a_mem[8][1] ),
    .A1(\b_to_a_mem[9][1] ),
    .A2(\b_to_a_mem[10][1] ),
    .A3(\b_to_a_mem[11][1] ),
    .S0(_126_),
    .S1(_124_),
    .X(_142_));
 sky130_fd_sc_hd__o22ai_2 _442_ (.A1(_131_),
    .A2(_141_),
    .B1(_142_),
    .B2(_130_),
    .Y(_143_));
 sky130_fd_sc_hd__nor2_1 _443_ (.A(_140_),
    .B(_143_),
    .Y(_144_));
 sky130_fd_sc_hd__mux2_1 _444_ (.A0(_144_),
    .A1(net27),
    .S(_135_),
    .X(_039_));
 sky130_fd_sc_hd__mux4_1 _445_ (.A0(\b_to_a_mem[2][2] ),
    .A1(\b_to_a_mem[3][2] ),
    .A2(\b_to_a_mem[6][2] ),
    .A3(\b_to_a_mem[7][2] ),
    .S0(_136_),
    .S1(_121_),
    .X(_145_));
 sky130_fd_sc_hd__mux4_1 _446_ (.A0(\b_to_a_mem[0][2] ),
    .A1(\b_to_a_mem[1][2] ),
    .A2(\b_to_a_mem[4][2] ),
    .A3(\b_to_a_mem[5][2] ),
    .S0(_138_),
    .S1(_117_),
    .X(_146_));
 sky130_fd_sc_hd__o22ai_1 _447_ (.A1(_125_),
    .A2(_145_),
    .B1(_146_),
    .B2(_123_),
    .Y(_147_));
 sky130_fd_sc_hd__mux4_1 _448_ (.A0(\b_to_a_mem[12][2] ),
    .A1(\b_to_a_mem[13][2] ),
    .A2(\b_to_a_mem[14][2] ),
    .A3(\b_to_a_mem[15][2] ),
    .S0(_138_),
    .S1(_116_),
    .X(_148_));
 sky130_fd_sc_hd__mux4_1 _449_ (.A0(\b_to_a_mem[8][2] ),
    .A1(\b_to_a_mem[9][2] ),
    .A2(\b_to_a_mem[10][2] ),
    .A3(\b_to_a_mem[11][2] ),
    .S0(_126_),
    .S1(_124_),
    .X(_149_));
 sky130_fd_sc_hd__o22ai_2 _450_ (.A1(_131_),
    .A2(_148_),
    .B1(_149_),
    .B2(_130_),
    .Y(_150_));
 sky130_fd_sc_hd__nor2_1 _451_ (.A(_147_),
    .B(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__mux2_1 _452_ (.A0(_151_),
    .A1(net28),
    .S(_135_),
    .X(_040_));
 sky130_fd_sc_hd__mux4_2 _453_ (.A0(\b_to_a_mem[2][3] ),
    .A1(\b_to_a_mem[3][3] ),
    .A2(\b_to_a_mem[6][3] ),
    .A3(\b_to_a_mem[7][3] ),
    .S0(_136_),
    .S1(_121_),
    .X(_152_));
 sky130_fd_sc_hd__mux4_1 _454_ (.A0(\b_to_a_mem[0][3] ),
    .A1(\b_to_a_mem[1][3] ),
    .A2(\b_to_a_mem[4][3] ),
    .A3(\b_to_a_mem[5][3] ),
    .S0(_136_),
    .S1(_117_),
    .X(_153_));
 sky130_fd_sc_hd__o22ai_4 _455_ (.A1(_125_),
    .A2(_152_),
    .B1(_153_),
    .B2(_123_),
    .Y(_154_));
 sky130_fd_sc_hd__mux4_1 _456_ (.A0(\b_to_a_mem[12][3] ),
    .A1(\b_to_a_mem[13][3] ),
    .A2(\b_to_a_mem[14][3] ),
    .A3(\b_to_a_mem[15][3] ),
    .S0(_138_),
    .S1(_116_),
    .X(_155_));
 sky130_fd_sc_hd__mux4_1 _457_ (.A0(\b_to_a_mem[8][3] ),
    .A1(\b_to_a_mem[9][3] ),
    .A2(\b_to_a_mem[10][3] ),
    .A3(\b_to_a_mem[11][3] ),
    .S0(_126_),
    .S1(_124_),
    .X(_156_));
 sky130_fd_sc_hd__o22ai_1 _458_ (.A1(_131_),
    .A2(_155_),
    .B1(_156_),
    .B2(_130_),
    .Y(_157_));
 sky130_fd_sc_hd__nor2_1 _459_ (.A(_154_),
    .B(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__mux2_1 _460_ (.A0(_158_),
    .A1(net29),
    .S(_135_),
    .X(_041_));
 sky130_fd_sc_hd__mux4_1 _461_ (.A0(\b_to_a_mem[2][4] ),
    .A1(\b_to_a_mem[3][4] ),
    .A2(\b_to_a_mem[6][4] ),
    .A3(\b_to_a_mem[7][4] ),
    .S0(_136_),
    .S1(_121_),
    .X(_159_));
 sky130_fd_sc_hd__mux4_1 _462_ (.A0(\b_to_a_mem[0][4] ),
    .A1(\b_to_a_mem[1][4] ),
    .A2(\b_to_a_mem[4][4] ),
    .A3(\b_to_a_mem[5][4] ),
    .S0(_136_),
    .S1(_117_),
    .X(_160_));
 sky130_fd_sc_hd__o22ai_2 _463_ (.A1(_125_),
    .A2(_159_),
    .B1(_160_),
    .B2(_123_),
    .Y(_161_));
 sky130_fd_sc_hd__mux4_1 _464_ (.A0(\b_to_a_mem[12][4] ),
    .A1(\b_to_a_mem[13][4] ),
    .A2(\b_to_a_mem[14][4] ),
    .A3(\b_to_a_mem[15][4] ),
    .S0(_138_),
    .S1(_116_),
    .X(_162_));
 sky130_fd_sc_hd__mux4_1 _465_ (.A0(\b_to_a_mem[8][4] ),
    .A1(\b_to_a_mem[9][4] ),
    .A2(\b_to_a_mem[10][4] ),
    .A3(\b_to_a_mem[11][4] ),
    .S0(_126_),
    .S1(_124_),
    .X(_163_));
 sky130_fd_sc_hd__o22ai_1 _466_ (.A1(_131_),
    .A2(_162_),
    .B1(_163_),
    .B2(_130_),
    .Y(_164_));
 sky130_fd_sc_hd__nor2_1 _467_ (.A(_161_),
    .B(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__mux2_1 _468_ (.A0(_165_),
    .A1(net30),
    .S(_135_),
    .X(_042_));
 sky130_fd_sc_hd__mux4_1 _469_ (.A0(\b_to_a_mem[2][5] ),
    .A1(\b_to_a_mem[3][5] ),
    .A2(\b_to_a_mem[6][5] ),
    .A3(\b_to_a_mem[7][5] ),
    .S0(_136_),
    .S1(_121_),
    .X(_166_));
 sky130_fd_sc_hd__mux4_1 _470_ (.A0(\b_to_a_mem[0][5] ),
    .A1(\b_to_a_mem[1][5] ),
    .A2(\b_to_a_mem[4][5] ),
    .A3(\b_to_a_mem[5][5] ),
    .S0(_136_),
    .S1(_117_),
    .X(_167_));
 sky130_fd_sc_hd__o22ai_2 _471_ (.A1(_125_),
    .A2(_166_),
    .B1(_167_),
    .B2(_123_),
    .Y(_168_));
 sky130_fd_sc_hd__mux4_1 _472_ (.A0(\b_to_a_mem[12][5] ),
    .A1(\b_to_a_mem[13][5] ),
    .A2(\b_to_a_mem[14][5] ),
    .A3(\b_to_a_mem[15][5] ),
    .S0(_138_),
    .S1(_116_),
    .X(_169_));
 sky130_fd_sc_hd__mux4_1 _473_ (.A0(\b_to_a_mem[8][5] ),
    .A1(\b_to_a_mem[9][5] ),
    .A2(\b_to_a_mem[10][5] ),
    .A3(\b_to_a_mem[11][5] ),
    .S0(_126_),
    .S1(_124_),
    .X(_170_));
 sky130_fd_sc_hd__o22ai_1 _474_ (.A1(_131_),
    .A2(_169_),
    .B1(_170_),
    .B2(_130_),
    .Y(_171_));
 sky130_fd_sc_hd__nor2_1 _475_ (.A(_168_),
    .B(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__mux2_1 _476_ (.A0(_172_),
    .A1(net31),
    .S(_135_),
    .X(_043_));
 sky130_fd_sc_hd__mux4_1 _477_ (.A0(\b_to_a_mem[2][6] ),
    .A1(\b_to_a_mem[3][6] ),
    .A2(\b_to_a_mem[6][6] ),
    .A3(\b_to_a_mem[7][6] ),
    .S0(_120_),
    .S1(_121_),
    .X(_173_));
 sky130_fd_sc_hd__mux4_1 _478_ (.A0(\b_to_a_mem[0][6] ),
    .A1(\b_to_a_mem[1][6] ),
    .A2(\b_to_a_mem[4][6] ),
    .A3(\b_to_a_mem[5][6] ),
    .S0(_136_),
    .S1(_121_),
    .X(_174_));
 sky130_fd_sc_hd__o22ai_2 _479_ (.A1(_125_),
    .A2(_173_),
    .B1(_174_),
    .B2(_123_),
    .Y(_175_));
 sky130_fd_sc_hd__mux4_1 _480_ (.A0(\b_to_a_mem[12][6] ),
    .A1(\b_to_a_mem[13][6] ),
    .A2(\b_to_a_mem[14][6] ),
    .A3(\b_to_a_mem[15][6] ),
    .S0(_138_),
    .S1(_116_),
    .X(_176_));
 sky130_fd_sc_hd__mux4_1 _481_ (.A0(\b_to_a_mem[8][6] ),
    .A1(\b_to_a_mem[9][6] ),
    .A2(\b_to_a_mem[10][6] ),
    .A3(\b_to_a_mem[11][6] ),
    .S0(_126_),
    .S1(_124_),
    .X(_177_));
 sky130_fd_sc_hd__o22ai_1 _482_ (.A1(_131_),
    .A2(_176_),
    .B1(_177_),
    .B2(_130_),
    .Y(_178_));
 sky130_fd_sc_hd__nor2_1 _483_ (.A(_175_),
    .B(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__mux2_1 _484_ (.A0(_179_),
    .A1(net32),
    .S(_135_),
    .X(_044_));
 sky130_fd_sc_hd__mux4_1 _485_ (.A0(\b_to_a_mem[2][7] ),
    .A1(\b_to_a_mem[3][7] ),
    .A2(\b_to_a_mem[6][7] ),
    .A3(\b_to_a_mem[7][7] ),
    .S0(_120_),
    .S1(_121_),
    .X(_180_));
 sky130_fd_sc_hd__mux4_1 _486_ (.A0(\b_to_a_mem[0][7] ),
    .A1(\b_to_a_mem[1][7] ),
    .A2(\b_to_a_mem[4][7] ),
    .A3(\b_to_a_mem[5][7] ),
    .S0(_136_),
    .S1(_121_),
    .X(_181_));
 sky130_fd_sc_hd__o22ai_2 _487_ (.A1(_125_),
    .A2(_180_),
    .B1(_181_),
    .B2(_123_),
    .Y(_182_));
 sky130_fd_sc_hd__mux4_1 _488_ (.A0(\b_to_a_mem[12][7] ),
    .A1(\b_to_a_mem[13][7] ),
    .A2(\b_to_a_mem[14][7] ),
    .A3(\b_to_a_mem[15][7] ),
    .S0(_138_),
    .S1(_116_),
    .X(_183_));
 sky130_fd_sc_hd__mux4_1 _489_ (.A0(\b_to_a_mem[8][7] ),
    .A1(\b_to_a_mem[9][7] ),
    .A2(\b_to_a_mem[10][7] ),
    .A3(\b_to_a_mem[11][7] ),
    .S0(_138_),
    .S1(_124_),
    .X(_184_));
 sky130_fd_sc_hd__o22ai_2 _490_ (.A1(_131_),
    .A2(_183_),
    .B1(_184_),
    .B2(_130_),
    .Y(_185_));
 sky130_fd_sc_hd__nor2_1 _491_ (.A(_182_),
    .B(_185_),
    .Y(_186_));
 sky130_fd_sc_hd__mux2_1 _492_ (.A0(_186_),
    .A1(net33),
    .S(_135_),
    .X(_045_));
 sky130_fd_sc_hd__xnor2_1 _493_ (.A(_126_),
    .B(_135_),
    .Y(_046_));
 sky130_fd_sc_hd__mux2_1 _494_ (.A0(_037_),
    .A1(_124_),
    .S(_135_),
    .X(_047_));
 sky130_fd_sc_hd__o211ai_1 _495_ (.A1(net55),
    .A2(_096_),
    .B1(net2),
    .C1(_303_),
    .Y(_187_));
 sky130_fd_sc_hd__xnor2_1 _496_ (.A(_117_),
    .B(_187_),
    .Y(_048_));
 sky130_fd_sc_hd__nand2_1 _497_ (.A(net2),
    .B(_126_),
    .Y(_188_));
 sky130_fd_sc_hd__nor3_1 _498_ (.A(_272_),
    .B(_288_),
    .C(_188_),
    .Y(_189_));
 sky130_fd_sc_hd__o21ai_0 _499_ (.A1(net55),
    .A2(_096_),
    .B1(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__xnor2_1 _500_ (.A(\a_rd_ptr[3] ),
    .B(_190_),
    .Y(_049_));
 sky130_fd_sc_hd__and4_1 _501_ (.A(net2),
    .B(_117_),
    .C(\a_rd_ptr[3] ),
    .D(_303_),
    .X(_191_));
 sky130_fd_sc_hd__o21ai_1 _502_ (.A1(net55),
    .A2(_096_),
    .B1(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__xnor2_1 _503_ (.A(\a_rd_ptr[4] ),
    .B(_192_),
    .Y(_050_));
 sky130_fd_sc_hd__xnor2_1 _504_ (.A(_032_),
    .B(_102_),
    .Y(_051_));
 sky130_fd_sc_hd__mux2_1 _505_ (.A0(\a_wr_ptr[1] ),
    .A1(_033_),
    .S(_099_),
    .X(_052_));
 sky130_fd_sc_hd__xor2_1 _506_ (.A(\a_wr_ptr[2] ),
    .B(_101_),
    .X(_053_));
 sky130_fd_sc_hd__nand4_1 _507_ (.A(net11),
    .B(\a_wr_ptr[2] ),
    .C(\a_wr_ptr[1] ),
    .D(\a_wr_ptr[0] ),
    .Y(_193_));
 sky130_fd_sc_hd__a21oi_1 _508_ (.A1(net38),
    .A2(_092_),
    .B1(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__xor2_1 _509_ (.A(\a_wr_ptr[3] ),
    .B(_194_),
    .X(_054_));
 sky130_fd_sc_hd__xor2_1 _510_ (.A(\a_wr_ptr[4] ),
    .B(_006_),
    .X(_055_));
 sky130_fd_sc_hd__clkbuf_4 _511_ (.A(\b_rd_ptr[0] ),
    .X(_195_));
 sky130_fd_sc_hd__buf_4 _512_ (.A(\b_rd_ptr[2] ),
    .X(_196_));
 sky130_fd_sc_hd__mux4_1 _513_ (.A0(\a_to_b_mem[0][0] ),
    .A1(\a_to_b_mem[1][0] ),
    .A2(\a_to_b_mem[4][0] ),
    .A3(\a_to_b_mem[5][0] ),
    .S0(_195_),
    .S1(_196_),
    .X(_197_));
 sky130_fd_sc_hd__nand2_4 _514_ (.A(_275_),
    .B(_283_),
    .Y(_198_));
 sky130_fd_sc_hd__buf_4 _515_ (.A(_118_),
    .X(_199_));
 sky130_fd_sc_hd__nand2_4 _516_ (.A(_199_),
    .B(_283_),
    .Y(_200_));
 sky130_fd_sc_hd__buf_6 _517_ (.A(_195_),
    .X(_201_));
 sky130_fd_sc_hd__mux4_1 _518_ (.A0(\a_to_b_mem[2][0] ),
    .A1(\a_to_b_mem[3][0] ),
    .A2(\a_to_b_mem[6][0] ),
    .A3(\a_to_b_mem[7][0] ),
    .S0(_201_),
    .S1(_119_),
    .X(_202_));
 sky130_fd_sc_hd__o22ai_1 _519_ (.A1(_197_),
    .A2(_198_),
    .B1(_200_),
    .B2(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__mux4_1 _520_ (.A0(\a_to_b_mem[8][0] ),
    .A1(\a_to_b_mem[9][0] ),
    .A2(\a_to_b_mem[10][0] ),
    .A3(\a_to_b_mem[11][0] ),
    .S0(_195_),
    .S1(_118_),
    .X(_204_));
 sky130_fd_sc_hd__nand2_8 _521_ (.A(_291_),
    .B(\b_rd_ptr[3] ),
    .Y(_205_));
 sky130_fd_sc_hd__nand2_8 _522_ (.A(_119_),
    .B(\b_rd_ptr[3] ),
    .Y(_206_));
 sky130_fd_sc_hd__mux4_1 _523_ (.A0(\a_to_b_mem[12][0] ),
    .A1(\a_to_b_mem[13][0] ),
    .A2(\a_to_b_mem[14][0] ),
    .A3(\a_to_b_mem[15][0] ),
    .S0(_201_),
    .S1(_199_),
    .X(_207_));
 sky130_fd_sc_hd__o22ai_1 _524_ (.A1(_204_),
    .A2(_205_),
    .B1(_206_),
    .B2(_207_),
    .Y(_208_));
 sky130_fd_sc_hd__nor2_1 _525_ (.A(_203_),
    .B(_208_),
    .Y(_209_));
 sky130_fd_sc_hd__o21ai_4 _526_ (.A1(_089_),
    .A2(_097_),
    .B1(net12),
    .Y(_210_));
 sky130_fd_sc_hd__mux2_1 _527_ (.A0(_209_),
    .A1(net43),
    .S(_210_),
    .X(_056_));
 sky130_fd_sc_hd__buf_4 _528_ (.A(_195_),
    .X(_211_));
 sky130_fd_sc_hd__mux4_1 _529_ (.A0(\a_to_b_mem[2][1] ),
    .A1(\a_to_b_mem[3][1] ),
    .A2(\a_to_b_mem[6][1] ),
    .A3(\a_to_b_mem[7][1] ),
    .S0(_211_),
    .S1(_196_),
    .X(_212_));
 sky130_fd_sc_hd__clkbuf_8 _530_ (.A(_195_),
    .X(_213_));
 sky130_fd_sc_hd__mux4_1 _531_ (.A0(\a_to_b_mem[0][1] ),
    .A1(\a_to_b_mem[1][1] ),
    .A2(\a_to_b_mem[4][1] ),
    .A3(\a_to_b_mem[5][1] ),
    .S0(_213_),
    .S1(_119_),
    .X(_214_));
 sky130_fd_sc_hd__o22ai_1 _532_ (.A1(_200_),
    .A2(_212_),
    .B1(_214_),
    .B2(_198_),
    .Y(_215_));
 sky130_fd_sc_hd__mux4_1 _533_ (.A0(\a_to_b_mem[12][1] ),
    .A1(\a_to_b_mem[13][1] ),
    .A2(\a_to_b_mem[14][1] ),
    .A3(\a_to_b_mem[15][1] ),
    .S0(_213_),
    .S1(_118_),
    .X(_216_));
 sky130_fd_sc_hd__mux4_2 _534_ (.A0(\a_to_b_mem[8][1] ),
    .A1(\a_to_b_mem[9][1] ),
    .A2(\a_to_b_mem[10][1] ),
    .A3(\a_to_b_mem[11][1] ),
    .S0(_201_),
    .S1(_199_),
    .X(_217_));
 sky130_fd_sc_hd__o22ai_2 _535_ (.A1(_206_),
    .A2(_216_),
    .B1(_217_),
    .B2(_205_),
    .Y(_218_));
 sky130_fd_sc_hd__nor2_1 _536_ (.A(_215_),
    .B(_218_),
    .Y(_219_));
 sky130_fd_sc_hd__mux2_1 _537_ (.A0(_219_),
    .A1(net44),
    .S(_210_),
    .X(_057_));
 sky130_fd_sc_hd__mux4_1 _538_ (.A0(\a_to_b_mem[2][2] ),
    .A1(\a_to_b_mem[3][2] ),
    .A2(\a_to_b_mem[6][2] ),
    .A3(\a_to_b_mem[7][2] ),
    .S0(_211_),
    .S1(_196_),
    .X(_220_));
 sky130_fd_sc_hd__mux4_1 _539_ (.A0(\a_to_b_mem[0][2] ),
    .A1(\a_to_b_mem[1][2] ),
    .A2(\a_to_b_mem[4][2] ),
    .A3(\a_to_b_mem[5][2] ),
    .S0(_213_),
    .S1(_119_),
    .X(_221_));
 sky130_fd_sc_hd__o22ai_1 _540_ (.A1(_200_),
    .A2(_220_),
    .B1(_221_),
    .B2(_198_),
    .Y(_222_));
 sky130_fd_sc_hd__mux4_1 _541_ (.A0(\a_to_b_mem[12][2] ),
    .A1(\a_to_b_mem[13][2] ),
    .A2(\a_to_b_mem[14][2] ),
    .A3(\a_to_b_mem[15][2] ),
    .S0(_213_),
    .S1(_118_),
    .X(_223_));
 sky130_fd_sc_hd__mux4_1 _542_ (.A0(\a_to_b_mem[8][2] ),
    .A1(\a_to_b_mem[9][2] ),
    .A2(\a_to_b_mem[10][2] ),
    .A3(\a_to_b_mem[11][2] ),
    .S0(_201_),
    .S1(_199_),
    .X(_224_));
 sky130_fd_sc_hd__o22ai_2 _543_ (.A1(_206_),
    .A2(_223_),
    .B1(_224_),
    .B2(_205_),
    .Y(_225_));
 sky130_fd_sc_hd__nor2_1 _544_ (.A(_222_),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__mux2_1 _545_ (.A0(_226_),
    .A1(net45),
    .S(_210_),
    .X(_058_));
 sky130_fd_sc_hd__mux4_1 _546_ (.A0(\a_to_b_mem[2][3] ),
    .A1(\a_to_b_mem[3][3] ),
    .A2(\a_to_b_mem[6][3] ),
    .A3(\a_to_b_mem[7][3] ),
    .S0(_211_),
    .S1(_196_),
    .X(_227_));
 sky130_fd_sc_hd__mux4_1 _547_ (.A0(\a_to_b_mem[0][3] ),
    .A1(\a_to_b_mem[1][3] ),
    .A2(\a_to_b_mem[4][3] ),
    .A3(\a_to_b_mem[5][3] ),
    .S0(_211_),
    .S1(_119_),
    .X(_228_));
 sky130_fd_sc_hd__o22ai_1 _548_ (.A1(_200_),
    .A2(_227_),
    .B1(_228_),
    .B2(_198_),
    .Y(_229_));
 sky130_fd_sc_hd__mux4_1 _549_ (.A0(\a_to_b_mem[12][3] ),
    .A1(\a_to_b_mem[13][3] ),
    .A2(\a_to_b_mem[14][3] ),
    .A3(\a_to_b_mem[15][3] ),
    .S0(_213_),
    .S1(_118_),
    .X(_230_));
 sky130_fd_sc_hd__mux4_1 _550_ (.A0(\a_to_b_mem[8][3] ),
    .A1(\a_to_b_mem[9][3] ),
    .A2(\a_to_b_mem[10][3] ),
    .A3(\a_to_b_mem[11][3] ),
    .S0(_201_),
    .S1(_199_),
    .X(_231_));
 sky130_fd_sc_hd__o22ai_1 _551_ (.A1(_206_),
    .A2(_230_),
    .B1(_231_),
    .B2(_205_),
    .Y(_232_));
 sky130_fd_sc_hd__nor2_1 _552_ (.A(_229_),
    .B(_232_),
    .Y(_233_));
 sky130_fd_sc_hd__mux2_1 _553_ (.A0(_233_),
    .A1(net46),
    .S(_210_),
    .X(_059_));
 sky130_fd_sc_hd__mux4_1 _554_ (.A0(\a_to_b_mem[2][4] ),
    .A1(\a_to_b_mem[3][4] ),
    .A2(\a_to_b_mem[6][4] ),
    .A3(\a_to_b_mem[7][4] ),
    .S0(_211_),
    .S1(_196_),
    .X(_234_));
 sky130_fd_sc_hd__mux4_1 _555_ (.A0(\a_to_b_mem[0][4] ),
    .A1(\a_to_b_mem[1][4] ),
    .A2(\a_to_b_mem[4][4] ),
    .A3(\a_to_b_mem[5][4] ),
    .S0(_211_),
    .S1(_119_),
    .X(_235_));
 sky130_fd_sc_hd__o22ai_1 _556_ (.A1(_200_),
    .A2(_234_),
    .B1(_235_),
    .B2(_198_),
    .Y(_236_));
 sky130_fd_sc_hd__mux4_2 _557_ (.A0(\a_to_b_mem[12][4] ),
    .A1(\a_to_b_mem[13][4] ),
    .A2(\a_to_b_mem[14][4] ),
    .A3(\a_to_b_mem[15][4] ),
    .S0(_213_),
    .S1(_118_),
    .X(_237_));
 sky130_fd_sc_hd__mux4_2 _558_ (.A0(\a_to_b_mem[8][4] ),
    .A1(\a_to_b_mem[9][4] ),
    .A2(\a_to_b_mem[10][4] ),
    .A3(\a_to_b_mem[11][4] ),
    .S0(_201_),
    .S1(_199_),
    .X(_238_));
 sky130_fd_sc_hd__o22ai_4 _559_ (.A1(_206_),
    .A2(_237_),
    .B1(_238_),
    .B2(_205_),
    .Y(_239_));
 sky130_fd_sc_hd__nor2_1 _560_ (.A(_236_),
    .B(_239_),
    .Y(_240_));
 sky130_fd_sc_hd__mux2_1 _561_ (.A0(_240_),
    .A1(net47),
    .S(_210_),
    .X(_060_));
 sky130_fd_sc_hd__mux4_1 _562_ (.A0(\a_to_b_mem[2][5] ),
    .A1(\a_to_b_mem[3][5] ),
    .A2(\a_to_b_mem[6][5] ),
    .A3(\a_to_b_mem[7][5] ),
    .S0(_211_),
    .S1(_196_),
    .X(_241_));
 sky130_fd_sc_hd__mux4_1 _563_ (.A0(\a_to_b_mem[0][5] ),
    .A1(\a_to_b_mem[1][5] ),
    .A2(\a_to_b_mem[4][5] ),
    .A3(\a_to_b_mem[5][5] ),
    .S0(_211_),
    .S1(_119_),
    .X(_242_));
 sky130_fd_sc_hd__o22ai_1 _564_ (.A1(_200_),
    .A2(_241_),
    .B1(_242_),
    .B2(_198_),
    .Y(_243_));
 sky130_fd_sc_hd__mux4_1 _565_ (.A0(\a_to_b_mem[12][5] ),
    .A1(\a_to_b_mem[13][5] ),
    .A2(\a_to_b_mem[14][5] ),
    .A3(\a_to_b_mem[15][5] ),
    .S0(_213_),
    .S1(_118_),
    .X(_244_));
 sky130_fd_sc_hd__mux4_1 _566_ (.A0(\a_to_b_mem[8][5] ),
    .A1(\a_to_b_mem[9][5] ),
    .A2(\a_to_b_mem[10][5] ),
    .A3(\a_to_b_mem[11][5] ),
    .S0(_201_),
    .S1(_199_),
    .X(_245_));
 sky130_fd_sc_hd__o22ai_1 _567_ (.A1(_206_),
    .A2(_244_),
    .B1(_245_),
    .B2(_205_),
    .Y(_246_));
 sky130_fd_sc_hd__nor2_1 _568_ (.A(_243_),
    .B(_246_),
    .Y(_247_));
 sky130_fd_sc_hd__mux2_1 _569_ (.A0(_247_),
    .A1(net48),
    .S(_210_),
    .X(_061_));
 sky130_fd_sc_hd__mux4_1 _570_ (.A0(\a_to_b_mem[2][6] ),
    .A1(\a_to_b_mem[3][6] ),
    .A2(\a_to_b_mem[6][6] ),
    .A3(\a_to_b_mem[7][6] ),
    .S0(_195_),
    .S1(_196_),
    .X(_248_));
 sky130_fd_sc_hd__mux4_1 _571_ (.A0(\a_to_b_mem[0][6] ),
    .A1(\a_to_b_mem[1][6] ),
    .A2(\a_to_b_mem[4][6] ),
    .A3(\a_to_b_mem[5][6] ),
    .S0(_211_),
    .S1(_196_),
    .X(_249_));
 sky130_fd_sc_hd__o22ai_1 _572_ (.A1(_200_),
    .A2(_248_),
    .B1(_249_),
    .B2(_198_),
    .Y(_250_));
 sky130_fd_sc_hd__mux4_1 _573_ (.A0(\a_to_b_mem[12][6] ),
    .A1(\a_to_b_mem[13][6] ),
    .A2(\a_to_b_mem[14][6] ),
    .A3(\a_to_b_mem[15][6] ),
    .S0(_213_),
    .S1(_118_),
    .X(_251_));
 sky130_fd_sc_hd__mux4_2 _574_ (.A0(\a_to_b_mem[8][6] ),
    .A1(\a_to_b_mem[9][6] ),
    .A2(\a_to_b_mem[10][6] ),
    .A3(\a_to_b_mem[11][6] ),
    .S0(_201_),
    .S1(_199_),
    .X(_252_));
 sky130_fd_sc_hd__o22ai_4 _575_ (.A1(_206_),
    .A2(_251_),
    .B1(_252_),
    .B2(_205_),
    .Y(_253_));
 sky130_fd_sc_hd__nor2_1 _576_ (.A(_250_),
    .B(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__mux2_1 _577_ (.A0(_254_),
    .A1(net49),
    .S(_210_),
    .X(_062_));
 sky130_fd_sc_hd__mux4_1 _578_ (.A0(\a_to_b_mem[2][7] ),
    .A1(\a_to_b_mem[3][7] ),
    .A2(\a_to_b_mem[6][7] ),
    .A3(\a_to_b_mem[7][7] ),
    .S0(_195_),
    .S1(_196_),
    .X(_255_));
 sky130_fd_sc_hd__mux4_1 _579_ (.A0(\a_to_b_mem[0][7] ),
    .A1(\a_to_b_mem[1][7] ),
    .A2(\a_to_b_mem[4][7] ),
    .A3(\a_to_b_mem[5][7] ),
    .S0(_211_),
    .S1(_196_),
    .X(_256_));
 sky130_fd_sc_hd__o22ai_1 _580_ (.A1(_200_),
    .A2(_255_),
    .B1(_256_),
    .B2(_198_),
    .Y(_257_));
 sky130_fd_sc_hd__mux4_1 _581_ (.A0(\a_to_b_mem[12][7] ),
    .A1(\a_to_b_mem[13][7] ),
    .A2(\a_to_b_mem[14][7] ),
    .A3(\a_to_b_mem[15][7] ),
    .S0(_213_),
    .S1(_118_),
    .X(_258_));
 sky130_fd_sc_hd__mux4_1 _582_ (.A0(\a_to_b_mem[8][7] ),
    .A1(\a_to_b_mem[9][7] ),
    .A2(\a_to_b_mem[10][7] ),
    .A3(\a_to_b_mem[11][7] ),
    .S0(_213_),
    .S1(_199_),
    .X(_259_));
 sky130_fd_sc_hd__o22ai_4 _583_ (.A1(_206_),
    .A2(_258_),
    .B1(_259_),
    .B2(_205_),
    .Y(_260_));
 sky130_fd_sc_hd__nor2_1 _584_ (.A(_257_),
    .B(_260_),
    .Y(_261_));
 sky130_fd_sc_hd__mux2_1 _585_ (.A0(_261_),
    .A1(net50),
    .S(_210_),
    .X(_063_));
 sky130_fd_sc_hd__xnor2_1 _586_ (.A(_201_),
    .B(_210_),
    .Y(_064_));
 sky130_fd_sc_hd__mux2_1 _587_ (.A0(_034_),
    .A1(_199_),
    .S(_210_),
    .X(_065_));
 sky130_fd_sc_hd__o211ai_1 _588_ (.A1(net38),
    .A2(_097_),
    .B1(net12),
    .C1(_294_),
    .Y(_262_));
 sky130_fd_sc_hd__xnor2_1 _589_ (.A(_119_),
    .B(_262_),
    .Y(_066_));
 sky130_fd_sc_hd__nand2_1 _590_ (.A(net12),
    .B(_201_),
    .Y(_263_));
 sky130_fd_sc_hd__nor3_1 _591_ (.A(_275_),
    .B(_291_),
    .C(_263_),
    .Y(_264_));
 sky130_fd_sc_hd__o21ai_0 _592_ (.A1(net38),
    .A2(_097_),
    .B1(_264_),
    .Y(_265_));
 sky130_fd_sc_hd__xnor2_1 _593_ (.A(\b_rd_ptr[3] ),
    .B(_265_),
    .Y(_067_));
 sky130_fd_sc_hd__and4_1 _594_ (.A(net12),
    .B(_119_),
    .C(\b_rd_ptr[3] ),
    .D(_294_),
    .X(_266_));
 sky130_fd_sc_hd__o21ai_0 _595_ (.A1(net38),
    .A2(_097_),
    .B1(_266_),
    .Y(_267_));
 sky130_fd_sc_hd__xnor2_1 _596_ (.A(\b_rd_ptr[4] ),
    .B(_267_),
    .Y(_068_));
 sky130_fd_sc_hd__xnor2_1 _597_ (.A(_035_),
    .B(_111_),
    .Y(_069_));
 sky130_fd_sc_hd__mux2_1 _598_ (.A0(\b_wr_ptr[1] ),
    .A1(_036_),
    .S(_108_),
    .X(_070_));
 sky130_fd_sc_hd__xor2_1 _599_ (.A(\b_wr_ptr[2] ),
    .B(_110_),
    .X(_071_));
 sky130_fd_sc_hd__nand4_1 _600_ (.A(net21),
    .B(\b_wr_ptr[2] ),
    .C(\b_wr_ptr[1] ),
    .D(\b_wr_ptr[0] ),
    .Y(_268_));
 sky130_fd_sc_hd__a21oi_1 _601_ (.A1(net55),
    .A2(_095_),
    .B1(_268_),
    .Y(_269_));
 sky130_fd_sc_hd__xor2_1 _602_ (.A(\b_wr_ptr[3] ),
    .B(_269_),
    .X(_072_));
 sky130_fd_sc_hd__xor2_1 _603_ (.A(\b_wr_ptr[4] ),
    .B(_022_),
    .X(_073_));
 sky130_fd_sc_hd__xor2_1 _604_ (.A(_315_),
    .B(net52),
    .X(_270_));
 sky130_fd_sc_hd__nor4_1 _605_ (.A(net53),
    .B(net54),
    .C(net55),
    .D(_270_),
    .Y(net22));
 sky130_fd_sc_hd__a31o_1 _606_ (.A1(net52),
    .A2(net53),
    .A3(net54),
    .B1(net55),
    .X(net23));
 sky130_fd_sc_hd__xor2_1 _607_ (.A(_313_),
    .B(net35),
    .X(_271_));
 sky130_fd_sc_hd__nor4_1 _608_ (.A(net37),
    .B(net36),
    .C(net38),
    .D(_271_),
    .Y(net39));
 sky130_fd_sc_hd__a31o_1 _609_ (.A1(net35),
    .A2(net37),
    .A3(net36),
    .B1(net38),
    .X(net40));
 sky130_fd_sc_hd__fa_2 _610_ (.A(_272_),
    .B(\b_wr_ptr[1] ),
    .CIN(_273_),
    .COUT(_274_),
    .SUM(net52));
 sky130_fd_sc_hd__fa_4 _611_ (.A(\a_wr_ptr[1] ),
    .B(_275_),
    .CIN(_276_),
    .COUT(_277_),
    .SUM(net35));
 sky130_fd_sc_hd__ha_1 _612_ (.A(_278_),
    .B(\b_wr_ptr[3] ),
    .COUT(_279_),
    .SUM(_280_));
 sky130_fd_sc_hd__ha_1 _613_ (.A(_272_),
    .B(\b_wr_ptr[1] ),
    .COUT(_281_),
    .SUM(_282_));
 sky130_fd_sc_hd__ha_1 _614_ (.A(\a_wr_ptr[3] ),
    .B(_283_),
    .COUT(_284_),
    .SUM(_285_));
 sky130_fd_sc_hd__ha_1 _615_ (.A(\a_wr_ptr[1] ),
    .B(_275_),
    .COUT(_286_),
    .SUM(_287_));
 sky130_fd_sc_hd__ha_1 _616_ (.A(_288_),
    .B(\b_wr_ptr[2] ),
    .COUT(_289_),
    .SUM(_290_));
 sky130_fd_sc_hd__ha_2 _617_ (.A(\a_wr_ptr[2] ),
    .B(_291_),
    .COUT(_292_),
    .SUM(_293_));
 sky130_fd_sc_hd__ha_1 _618_ (.A(\b_rd_ptr[0] ),
    .B(\b_rd_ptr[1] ),
    .COUT(_294_),
    .SUM(_034_));
 sky130_fd_sc_hd__ha_1 _619_ (.A(_035_),
    .B(_295_),
    .COUT(_296_),
    .SUM(_036_));
 sky130_fd_sc_hd__ha_1 _620_ (.A(_035_),
    .B(\b_wr_ptr[1] ),
    .COUT(_297_),
    .SUM(_298_));
 sky130_fd_sc_hd__ha_1 _621_ (.A(\b_wr_ptr[0] ),
    .B(_295_),
    .COUT(_299_),
    .SUM(_300_));
 sky130_fd_sc_hd__ha_1 _622_ (.A(\b_wr_ptr[0] ),
    .B(\b_wr_ptr[1] ),
    .COUT(_301_),
    .SUM(_302_));
 sky130_fd_sc_hd__ha_1 _623_ (.A(\a_rd_ptr[0] ),
    .B(\a_rd_ptr[1] ),
    .COUT(_303_),
    .SUM(_037_));
 sky130_fd_sc_hd__ha_1 _624_ (.A(_032_),
    .B(_304_),
    .COUT(_305_),
    .SUM(_033_));
 sky130_fd_sc_hd__ha_1 _625_ (.A(_032_),
    .B(\a_wr_ptr[1] ),
    .COUT(_306_),
    .SUM(_307_));
 sky130_fd_sc_hd__ha_1 _626_ (.A(\a_wr_ptr[0] ),
    .B(_304_),
    .COUT(_308_),
    .SUM(_309_));
 sky130_fd_sc_hd__ha_1 _627_ (.A(\a_wr_ptr[0] ),
    .B(\a_wr_ptr[1] ),
    .COUT(_310_),
    .SUM(_311_));
 sky130_fd_sc_hd__ha_1 _628_ (.A(_032_),
    .B(\b_rd_ptr[0] ),
    .COUT(_312_),
    .SUM(_313_));
 sky130_fd_sc_hd__ha_1 _629_ (.A(\a_rd_ptr[0] ),
    .B(_035_),
    .COUT(_314_),
    .SUM(_315_));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_data_reg[0]$_DFFE_PN0P_  (.D(_038_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_data_reg[1]$_DFFE_PN0P_  (.D(_039_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_data_reg[2]$_DFFE_PN0P_  (.D(_040_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_data_reg[3]$_DFFE_PN0P_  (.D(_041_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_data_reg[4]$_DFFE_PN0P_  (.D(_042_),
    .Q(net30),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_data_reg[5]$_DFFE_PN0P_  (.D(_043_),
    .Q(net31),
    .RESET_B(net1),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_data_reg[6]$_DFFE_PN0P_  (.D(_044_),
    .Q(net32),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_data_reg[7]$_DFFE_PN0P_  (.D(_045_),
    .Q(net33),
    .RESET_B(net1),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_ptr[0]$_DFFE_PN0P_  (.D(_046_),
    .Q(\a_rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_ptr[1]$_DFFE_PN0P_  (.D(_047_),
    .Q(\a_rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_ptr[2]$_DFFE_PN0P_  (.D(_048_),
    .Q(\a_rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_4 \a_rd_ptr[3]$_DFFE_PN0P_  (.D(_049_),
    .Q(\a_rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_rd_ptr[4]$_DFFE_PN0P_  (.D(_050_),
    .Q(\a_rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[0][0]$_DFFE_PP_  (.D(net3),
    .DE(_000_),
    .Q(\a_to_b_mem[0][0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[0][1]$_DFFE_PP_  (.D(net4),
    .DE(_000_),
    .Q(\a_to_b_mem[0][1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[0][2]$_DFFE_PP_  (.D(net5),
    .DE(_000_),
    .Q(\a_to_b_mem[0][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[0][3]$_DFFE_PP_  (.D(net6),
    .DE(_000_),
    .Q(\a_to_b_mem[0][3] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[0][4]$_DFFE_PP_  (.D(net7),
    .DE(_000_),
    .Q(\a_to_b_mem[0][4] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[0][5]$_DFFE_PP_  (.D(net8),
    .DE(_000_),
    .Q(\a_to_b_mem[0][5] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[0][6]$_DFFE_PP_  (.D(net9),
    .DE(_000_),
    .Q(\a_to_b_mem[0][6] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[0][7]$_DFFE_PP_  (.D(net10),
    .DE(_000_),
    .Q(\a_to_b_mem[0][7] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[10][0]$_DFFE_PP_  (.D(net3),
    .DE(_001_),
    .Q(\a_to_b_mem[10][0] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[10][1]$_DFFE_PP_  (.D(net4),
    .DE(_001_),
    .Q(\a_to_b_mem[10][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[10][2]$_DFFE_PP_  (.D(net5),
    .DE(_001_),
    .Q(\a_to_b_mem[10][2] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[10][3]$_DFFE_PP_  (.D(net6),
    .DE(_001_),
    .Q(\a_to_b_mem[10][3] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[10][4]$_DFFE_PP_  (.D(net7),
    .DE(_001_),
    .Q(\a_to_b_mem[10][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[10][5]$_DFFE_PP_  (.D(net8),
    .DE(_001_),
    .Q(\a_to_b_mem[10][5] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[10][6]$_DFFE_PP_  (.D(net9),
    .DE(_001_),
    .Q(\a_to_b_mem[10][6] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[10][7]$_DFFE_PP_  (.D(net10),
    .DE(_001_),
    .Q(\a_to_b_mem[10][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[11][0]$_DFFE_PP_  (.D(net3),
    .DE(_002_),
    .Q(\a_to_b_mem[11][0] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[11][1]$_DFFE_PP_  (.D(net4),
    .DE(_002_),
    .Q(\a_to_b_mem[11][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[11][2]$_DFFE_PP_  (.D(net5),
    .DE(_002_),
    .Q(\a_to_b_mem[11][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[11][3]$_DFFE_PP_  (.D(net6),
    .DE(_002_),
    .Q(\a_to_b_mem[11][3] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[11][4]$_DFFE_PP_  (.D(net7),
    .DE(_002_),
    .Q(\a_to_b_mem[11][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[11][5]$_DFFE_PP_  (.D(net8),
    .DE(_002_),
    .Q(\a_to_b_mem[11][5] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[11][6]$_DFFE_PP_  (.D(net9),
    .DE(_002_),
    .Q(\a_to_b_mem[11][6] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[11][7]$_DFFE_PP_  (.D(net10),
    .DE(_002_),
    .Q(\a_to_b_mem[11][7] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[12][0]$_DFFE_PP_  (.D(net3),
    .DE(_003_),
    .Q(\a_to_b_mem[12][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[12][1]$_DFFE_PP_  (.D(net4),
    .DE(_003_),
    .Q(\a_to_b_mem[12][1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[12][2]$_DFFE_PP_  (.D(net5),
    .DE(_003_),
    .Q(\a_to_b_mem[12][2] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[12][3]$_DFFE_PP_  (.D(net6),
    .DE(_003_),
    .Q(\a_to_b_mem[12][3] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[12][4]$_DFFE_PP_  (.D(net7),
    .DE(_003_),
    .Q(\a_to_b_mem[12][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[12][5]$_DFFE_PP_  (.D(net8),
    .DE(_003_),
    .Q(\a_to_b_mem[12][5] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[12][6]$_DFFE_PP_  (.D(net9),
    .DE(_003_),
    .Q(\a_to_b_mem[12][6] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[12][7]$_DFFE_PP_  (.D(net10),
    .DE(_003_),
    .Q(\a_to_b_mem[12][7] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[13][0]$_DFFE_PP_  (.D(net3),
    .DE(_004_),
    .Q(\a_to_b_mem[13][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[13][1]$_DFFE_PP_  (.D(net4),
    .DE(_004_),
    .Q(\a_to_b_mem[13][1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[13][2]$_DFFE_PP_  (.D(net5),
    .DE(_004_),
    .Q(\a_to_b_mem[13][2] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[13][3]$_DFFE_PP_  (.D(net6),
    .DE(_004_),
    .Q(\a_to_b_mem[13][3] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[13][4]$_DFFE_PP_  (.D(net7),
    .DE(_004_),
    .Q(\a_to_b_mem[13][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[13][5]$_DFFE_PP_  (.D(net8),
    .DE(_004_),
    .Q(\a_to_b_mem[13][5] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[13][6]$_DFFE_PP_  (.D(net9),
    .DE(_004_),
    .Q(\a_to_b_mem[13][6] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[13][7]$_DFFE_PP_  (.D(net10),
    .DE(_004_),
    .Q(\a_to_b_mem[13][7] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[14][0]$_DFFE_PP_  (.D(net3),
    .DE(_005_),
    .Q(\a_to_b_mem[14][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[14][1]$_DFFE_PP_  (.D(net4),
    .DE(_005_),
    .Q(\a_to_b_mem[14][1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[14][2]$_DFFE_PP_  (.D(net5),
    .DE(_005_),
    .Q(\a_to_b_mem[14][2] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[14][3]$_DFFE_PP_  (.D(net6),
    .DE(_005_),
    .Q(\a_to_b_mem[14][3] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[14][4]$_DFFE_PP_  (.D(net7),
    .DE(_005_),
    .Q(\a_to_b_mem[14][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[14][5]$_DFFE_PP_  (.D(net8),
    .DE(_005_),
    .Q(\a_to_b_mem[14][5] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[14][6]$_DFFE_PP_  (.D(net9),
    .DE(_005_),
    .Q(\a_to_b_mem[14][6] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[14][7]$_DFFE_PP_  (.D(net10),
    .DE(_005_),
    .Q(\a_to_b_mem[14][7] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[15][0]$_DFFE_PP_  (.D(net3),
    .DE(_006_),
    .Q(\a_to_b_mem[15][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[15][1]$_DFFE_PP_  (.D(net4),
    .DE(_006_),
    .Q(\a_to_b_mem[15][1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[15][2]$_DFFE_PP_  (.D(net5),
    .DE(_006_),
    .Q(\a_to_b_mem[15][2] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[15][3]$_DFFE_PP_  (.D(net6),
    .DE(_006_),
    .Q(\a_to_b_mem[15][3] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[15][4]$_DFFE_PP_  (.D(net7),
    .DE(_006_),
    .Q(\a_to_b_mem[15][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[15][5]$_DFFE_PP_  (.D(net8),
    .DE(_006_),
    .Q(\a_to_b_mem[15][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[15][6]$_DFFE_PP_  (.D(net9),
    .DE(_006_),
    .Q(\a_to_b_mem[15][6] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[15][7]$_DFFE_PP_  (.D(net10),
    .DE(_006_),
    .Q(\a_to_b_mem[15][7] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[1][0]$_DFFE_PP_  (.D(net3),
    .DE(_007_),
    .Q(\a_to_b_mem[1][0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[1][1]$_DFFE_PP_  (.D(net4),
    .DE(_007_),
    .Q(\a_to_b_mem[1][1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[1][2]$_DFFE_PP_  (.D(net5),
    .DE(_007_),
    .Q(\a_to_b_mem[1][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[1][3]$_DFFE_PP_  (.D(net6),
    .DE(_007_),
    .Q(\a_to_b_mem[1][3] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[1][4]$_DFFE_PP_  (.D(net7),
    .DE(_007_),
    .Q(\a_to_b_mem[1][4] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[1][5]$_DFFE_PP_  (.D(net8),
    .DE(_007_),
    .Q(\a_to_b_mem[1][5] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[1][6]$_DFFE_PP_  (.D(net9),
    .DE(_007_),
    .Q(\a_to_b_mem[1][6] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[1][7]$_DFFE_PP_  (.D(net10),
    .DE(_007_),
    .Q(\a_to_b_mem[1][7] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[2][0]$_DFFE_PP_  (.D(net3),
    .DE(_008_),
    .Q(\a_to_b_mem[2][0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[2][1]$_DFFE_PP_  (.D(net4),
    .DE(_008_),
    .Q(\a_to_b_mem[2][1] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[2][2]$_DFFE_PP_  (.D(net5),
    .DE(_008_),
    .Q(\a_to_b_mem[2][2] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[2][3]$_DFFE_PP_  (.D(net6),
    .DE(_008_),
    .Q(\a_to_b_mem[2][3] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[2][4]$_DFFE_PP_  (.D(net7),
    .DE(_008_),
    .Q(\a_to_b_mem[2][4] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[2][5]$_DFFE_PP_  (.D(net8),
    .DE(_008_),
    .Q(\a_to_b_mem[2][5] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[2][6]$_DFFE_PP_  (.D(net9),
    .DE(_008_),
    .Q(\a_to_b_mem[2][6] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[2][7]$_DFFE_PP_  (.D(net10),
    .DE(_008_),
    .Q(\a_to_b_mem[2][7] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[3][0]$_DFFE_PP_  (.D(net3),
    .DE(_009_),
    .Q(\a_to_b_mem[3][0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[3][1]$_DFFE_PP_  (.D(net4),
    .DE(_009_),
    .Q(\a_to_b_mem[3][1] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[3][2]$_DFFE_PP_  (.D(net5),
    .DE(_009_),
    .Q(\a_to_b_mem[3][2] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[3][3]$_DFFE_PP_  (.D(net6),
    .DE(_009_),
    .Q(\a_to_b_mem[3][3] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[3][4]$_DFFE_PP_  (.D(net7),
    .DE(_009_),
    .Q(\a_to_b_mem[3][4] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[3][5]$_DFFE_PP_  (.D(net8),
    .DE(_009_),
    .Q(\a_to_b_mem[3][5] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[3][6]$_DFFE_PP_  (.D(net9),
    .DE(_009_),
    .Q(\a_to_b_mem[3][6] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[3][7]$_DFFE_PP_  (.D(net10),
    .DE(_009_),
    .Q(\a_to_b_mem[3][7] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[4][0]$_DFFE_PP_  (.D(net3),
    .DE(_010_),
    .Q(\a_to_b_mem[4][0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[4][1]$_DFFE_PP_  (.D(net4),
    .DE(_010_),
    .Q(\a_to_b_mem[4][1] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[4][2]$_DFFE_PP_  (.D(net5),
    .DE(_010_),
    .Q(\a_to_b_mem[4][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[4][3]$_DFFE_PP_  (.D(net6),
    .DE(_010_),
    .Q(\a_to_b_mem[4][3] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[4][4]$_DFFE_PP_  (.D(net7),
    .DE(_010_),
    .Q(\a_to_b_mem[4][4] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[4][5]$_DFFE_PP_  (.D(net8),
    .DE(_010_),
    .Q(\a_to_b_mem[4][5] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[4][6]$_DFFE_PP_  (.D(net9),
    .DE(_010_),
    .Q(\a_to_b_mem[4][6] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[4][7]$_DFFE_PP_  (.D(net10),
    .DE(_010_),
    .Q(\a_to_b_mem[4][7] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[5][0]$_DFFE_PP_  (.D(net3),
    .DE(_011_),
    .Q(\a_to_b_mem[5][0] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[5][1]$_DFFE_PP_  (.D(net4),
    .DE(_011_),
    .Q(\a_to_b_mem[5][1] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[5][2]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\a_to_b_mem[5][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[5][3]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\a_to_b_mem[5][3] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[5][4]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\a_to_b_mem[5][4] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[5][5]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\a_to_b_mem[5][5] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[5][6]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\a_to_b_mem[5][6] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[5][7]$_DFFE_PP_  (.D(net10),
    .DE(_011_),
    .Q(\a_to_b_mem[5][7] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[6][0]$_DFFE_PP_  (.D(net3),
    .DE(_012_),
    .Q(\a_to_b_mem[6][0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[6][1]$_DFFE_PP_  (.D(net4),
    .DE(_012_),
    .Q(\a_to_b_mem[6][1] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[6][2]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\a_to_b_mem[6][2] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[6][3]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\a_to_b_mem[6][3] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[6][4]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\a_to_b_mem[6][4] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[6][5]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\a_to_b_mem[6][5] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[6][6]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\a_to_b_mem[6][6] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[6][7]$_DFFE_PP_  (.D(net10),
    .DE(_012_),
    .Q(\a_to_b_mem[6][7] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[7][0]$_DFFE_PP_  (.D(net3),
    .DE(_013_),
    .Q(\a_to_b_mem[7][0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[7][1]$_DFFE_PP_  (.D(net4),
    .DE(_013_),
    .Q(\a_to_b_mem[7][1] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[7][2]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\a_to_b_mem[7][2] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[7][3]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\a_to_b_mem[7][3] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[7][4]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\a_to_b_mem[7][4] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[7][5]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\a_to_b_mem[7][5] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[7][6]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\a_to_b_mem[7][6] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[7][7]$_DFFE_PP_  (.D(net10),
    .DE(_013_),
    .Q(\a_to_b_mem[7][7] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[8][0]$_DFFE_PP_  (.D(net3),
    .DE(_014_),
    .Q(\a_to_b_mem[8][0] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[8][1]$_DFFE_PP_  (.D(net4),
    .DE(_014_),
    .Q(\a_to_b_mem[8][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[8][2]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\a_to_b_mem[8][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[8][3]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\a_to_b_mem[8][3] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[8][4]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\a_to_b_mem[8][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[8][5]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\a_to_b_mem[8][5] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[8][6]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\a_to_b_mem[8][6] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[8][7]$_DFFE_PP_  (.D(net10),
    .DE(_014_),
    .Q(\a_to_b_mem[8][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[9][0]$_DFFE_PP_  (.D(net3),
    .DE(_015_),
    .Q(\a_to_b_mem[9][0] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[9][1]$_DFFE_PP_  (.D(net4),
    .DE(_015_),
    .Q(\a_to_b_mem[9][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[9][2]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\a_to_b_mem[9][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[9][3]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\a_to_b_mem[9][3] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[9][4]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\a_to_b_mem[9][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[9][5]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\a_to_b_mem[9][5] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[9][6]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\a_to_b_mem[9][6] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \a_to_b_mem[9][7]$_DFFE_PP_  (.D(net10),
    .DE(_015_),
    .Q(\a_to_b_mem[9][7] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_wr_ptr[0]$_DFFE_PN0P_  (.D(_051_),
    .Q(\a_wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \a_wr_ptr[1]$_DFFE_PN0P_  (.D(_052_),
    .Q(\a_wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \a_wr_ptr[2]$_DFFE_PN0P_  (.D(_053_),
    .Q(\a_wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \a_wr_ptr[3]$_DFFE_PN0P_  (.D(_054_),
    .Q(\a_wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_wr_ptr[4]$_DFFE_PN0P_  (.D(_055_),
    .Q(\a_wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_data_reg[0]$_DFFE_PN0P_  (.D(_056_),
    .Q(net43),
    .RESET_B(net1),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_data_reg[1]$_DFFE_PN0P_  (.D(_057_),
    .Q(net44),
    .RESET_B(net1),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_data_reg[2]$_DFFE_PN0P_  (.D(_058_),
    .Q(net45),
    .RESET_B(net1),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_data_reg[3]$_DFFE_PN0P_  (.D(_059_),
    .Q(net46),
    .RESET_B(net1),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_data_reg[4]$_DFFE_PN0P_  (.D(_060_),
    .Q(net47),
    .RESET_B(net1),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_data_reg[5]$_DFFE_PN0P_  (.D(_061_),
    .Q(net48),
    .RESET_B(net1),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_data_reg[6]$_DFFE_PN0P_  (.D(_062_),
    .Q(net49),
    .RESET_B(net1),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_data_reg[7]$_DFFE_PN0P_  (.D(_063_),
    .Q(net50),
    .RESET_B(net1),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_ptr[0]$_DFFE_PN0P_  (.D(_064_),
    .Q(\b_rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_ptr[1]$_DFFE_PN0P_  (.D(_065_),
    .Q(\b_rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_ptr[2]$_DFFE_PN0P_  (.D(_066_),
    .Q(\b_rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \b_rd_ptr[3]$_DFFE_PN0P_  (.D(_067_),
    .Q(\b_rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_rd_ptr[4]$_DFFE_PN0P_  (.D(_068_),
    .Q(\b_rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[0][0]$_DFFE_PP_  (.D(net13),
    .DE(_016_),
    .Q(\b_to_a_mem[0][0] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[0][1]$_DFFE_PP_  (.D(net14),
    .DE(_016_),
    .Q(\b_to_a_mem[0][1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[0][2]$_DFFE_PP_  (.D(net15),
    .DE(_016_),
    .Q(\b_to_a_mem[0][2] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[0][3]$_DFFE_PP_  (.D(net16),
    .DE(_016_),
    .Q(\b_to_a_mem[0][3] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[0][4]$_DFFE_PP_  (.D(net17),
    .DE(_016_),
    .Q(\b_to_a_mem[0][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[0][5]$_DFFE_PP_  (.D(net18),
    .DE(_016_),
    .Q(\b_to_a_mem[0][5] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[0][6]$_DFFE_PP_  (.D(net19),
    .DE(_016_),
    .Q(\b_to_a_mem[0][6] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[0][7]$_DFFE_PP_  (.D(net20),
    .DE(_016_),
    .Q(\b_to_a_mem[0][7] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[10][0]$_DFFE_PP_  (.D(net13),
    .DE(_017_),
    .Q(\b_to_a_mem[10][0] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[10][1]$_DFFE_PP_  (.D(net14),
    .DE(_017_),
    .Q(\b_to_a_mem[10][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[10][2]$_DFFE_PP_  (.D(net15),
    .DE(_017_),
    .Q(\b_to_a_mem[10][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[10][3]$_DFFE_PP_  (.D(net16),
    .DE(_017_),
    .Q(\b_to_a_mem[10][3] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[10][4]$_DFFE_PP_  (.D(net17),
    .DE(_017_),
    .Q(\b_to_a_mem[10][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[10][5]$_DFFE_PP_  (.D(net18),
    .DE(_017_),
    .Q(\b_to_a_mem[10][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[10][6]$_DFFE_PP_  (.D(net19),
    .DE(_017_),
    .Q(\b_to_a_mem[10][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[10][7]$_DFFE_PP_  (.D(net20),
    .DE(_017_),
    .Q(\b_to_a_mem[10][7] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[11][0]$_DFFE_PP_  (.D(net13),
    .DE(_018_),
    .Q(\b_to_a_mem[11][0] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[11][1]$_DFFE_PP_  (.D(net14),
    .DE(_018_),
    .Q(\b_to_a_mem[11][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[11][2]$_DFFE_PP_  (.D(net15),
    .DE(_018_),
    .Q(\b_to_a_mem[11][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[11][3]$_DFFE_PP_  (.D(net16),
    .DE(_018_),
    .Q(\b_to_a_mem[11][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[11][4]$_DFFE_PP_  (.D(net17),
    .DE(_018_),
    .Q(\b_to_a_mem[11][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[11][5]$_DFFE_PP_  (.D(net18),
    .DE(_018_),
    .Q(\b_to_a_mem[11][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[11][6]$_DFFE_PP_  (.D(net19),
    .DE(_018_),
    .Q(\b_to_a_mem[11][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[11][7]$_DFFE_PP_  (.D(net20),
    .DE(_018_),
    .Q(\b_to_a_mem[11][7] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[12][0]$_DFFE_PP_  (.D(net13),
    .DE(_019_),
    .Q(\b_to_a_mem[12][0] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[12][1]$_DFFE_PP_  (.D(net14),
    .DE(_019_),
    .Q(\b_to_a_mem[12][1] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[12][2]$_DFFE_PP_  (.D(net15),
    .DE(_019_),
    .Q(\b_to_a_mem[12][2] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[12][3]$_DFFE_PP_  (.D(net16),
    .DE(_019_),
    .Q(\b_to_a_mem[12][3] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[12][4]$_DFFE_PP_  (.D(net17),
    .DE(_019_),
    .Q(\b_to_a_mem[12][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[12][5]$_DFFE_PP_  (.D(net18),
    .DE(_019_),
    .Q(\b_to_a_mem[12][5] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[12][6]$_DFFE_PP_  (.D(net19),
    .DE(_019_),
    .Q(\b_to_a_mem[12][6] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[12][7]$_DFFE_PP_  (.D(net20),
    .DE(_019_),
    .Q(\b_to_a_mem[12][7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[13][0]$_DFFE_PP_  (.D(net13),
    .DE(_020_),
    .Q(\b_to_a_mem[13][0] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[13][1]$_DFFE_PP_  (.D(net14),
    .DE(_020_),
    .Q(\b_to_a_mem[13][1] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[13][2]$_DFFE_PP_  (.D(net15),
    .DE(_020_),
    .Q(\b_to_a_mem[13][2] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[13][3]$_DFFE_PP_  (.D(net16),
    .DE(_020_),
    .Q(\b_to_a_mem[13][3] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[13][4]$_DFFE_PP_  (.D(net17),
    .DE(_020_),
    .Q(\b_to_a_mem[13][4] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[13][5]$_DFFE_PP_  (.D(net18),
    .DE(_020_),
    .Q(\b_to_a_mem[13][5] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[13][6]$_DFFE_PP_  (.D(net19),
    .DE(_020_),
    .Q(\b_to_a_mem[13][6] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[13][7]$_DFFE_PP_  (.D(net20),
    .DE(_020_),
    .Q(\b_to_a_mem[13][7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[14][0]$_DFFE_PP_  (.D(net13),
    .DE(_021_),
    .Q(\b_to_a_mem[14][0] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[14][1]$_DFFE_PP_  (.D(net14),
    .DE(_021_),
    .Q(\b_to_a_mem[14][1] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[14][2]$_DFFE_PP_  (.D(net15),
    .DE(_021_),
    .Q(\b_to_a_mem[14][2] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[14][3]$_DFFE_PP_  (.D(net16),
    .DE(_021_),
    .Q(\b_to_a_mem[14][3] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[14][4]$_DFFE_PP_  (.D(net17),
    .DE(_021_),
    .Q(\b_to_a_mem[14][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[14][5]$_DFFE_PP_  (.D(net18),
    .DE(_021_),
    .Q(\b_to_a_mem[14][5] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[14][6]$_DFFE_PP_  (.D(net19),
    .DE(_021_),
    .Q(\b_to_a_mem[14][6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[14][7]$_DFFE_PP_  (.D(net20),
    .DE(_021_),
    .Q(\b_to_a_mem[14][7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[15][0]$_DFFE_PP_  (.D(net13),
    .DE(_022_),
    .Q(\b_to_a_mem[15][0] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[15][1]$_DFFE_PP_  (.D(net14),
    .DE(_022_),
    .Q(\b_to_a_mem[15][1] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[15][2]$_DFFE_PP_  (.D(net15),
    .DE(_022_),
    .Q(\b_to_a_mem[15][2] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[15][3]$_DFFE_PP_  (.D(net16),
    .DE(_022_),
    .Q(\b_to_a_mem[15][3] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[15][4]$_DFFE_PP_  (.D(net17),
    .DE(_022_),
    .Q(\b_to_a_mem[15][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[15][5]$_DFFE_PP_  (.D(net18),
    .DE(_022_),
    .Q(\b_to_a_mem[15][5] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[15][6]$_DFFE_PP_  (.D(net19),
    .DE(_022_),
    .Q(\b_to_a_mem[15][6] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[15][7]$_DFFE_PP_  (.D(net20),
    .DE(_022_),
    .Q(\b_to_a_mem[15][7] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[1][0]$_DFFE_PP_  (.D(net13),
    .DE(_023_),
    .Q(\b_to_a_mem[1][0] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[1][1]$_DFFE_PP_  (.D(net14),
    .DE(_023_),
    .Q(\b_to_a_mem[1][1] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[1][2]$_DFFE_PP_  (.D(net15),
    .DE(_023_),
    .Q(\b_to_a_mem[1][2] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[1][3]$_DFFE_PP_  (.D(net16),
    .DE(_023_),
    .Q(\b_to_a_mem[1][3] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[1][4]$_DFFE_PP_  (.D(net17),
    .DE(_023_),
    .Q(\b_to_a_mem[1][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[1][5]$_DFFE_PP_  (.D(net18),
    .DE(_023_),
    .Q(\b_to_a_mem[1][5] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[1][6]$_DFFE_PP_  (.D(net19),
    .DE(_023_),
    .Q(\b_to_a_mem[1][6] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[1][7]$_DFFE_PP_  (.D(net20),
    .DE(_023_),
    .Q(\b_to_a_mem[1][7] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[2][0]$_DFFE_PP_  (.D(net13),
    .DE(_024_),
    .Q(\b_to_a_mem[2][0] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[2][1]$_DFFE_PP_  (.D(net14),
    .DE(_024_),
    .Q(\b_to_a_mem[2][1] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[2][2]$_DFFE_PP_  (.D(net15),
    .DE(_024_),
    .Q(\b_to_a_mem[2][2] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[2][3]$_DFFE_PP_  (.D(net16),
    .DE(_024_),
    .Q(\b_to_a_mem[2][3] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[2][4]$_DFFE_PP_  (.D(net17),
    .DE(_024_),
    .Q(\b_to_a_mem[2][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[2][5]$_DFFE_PP_  (.D(net18),
    .DE(_024_),
    .Q(\b_to_a_mem[2][5] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[2][6]$_DFFE_PP_  (.D(net19),
    .DE(_024_),
    .Q(\b_to_a_mem[2][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[2][7]$_DFFE_PP_  (.D(net20),
    .DE(_024_),
    .Q(\b_to_a_mem[2][7] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[3][0]$_DFFE_PP_  (.D(net13),
    .DE(_025_),
    .Q(\b_to_a_mem[3][0] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[3][1]$_DFFE_PP_  (.D(net14),
    .DE(_025_),
    .Q(\b_to_a_mem[3][1] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[3][2]$_DFFE_PP_  (.D(net15),
    .DE(_025_),
    .Q(\b_to_a_mem[3][2] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[3][3]$_DFFE_PP_  (.D(net16),
    .DE(_025_),
    .Q(\b_to_a_mem[3][3] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[3][4]$_DFFE_PP_  (.D(net17),
    .DE(_025_),
    .Q(\b_to_a_mem[3][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[3][5]$_DFFE_PP_  (.D(net18),
    .DE(_025_),
    .Q(\b_to_a_mem[3][5] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[3][6]$_DFFE_PP_  (.D(net19),
    .DE(_025_),
    .Q(\b_to_a_mem[3][6] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[3][7]$_DFFE_PP_  (.D(net20),
    .DE(_025_),
    .Q(\b_to_a_mem[3][7] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[4][0]$_DFFE_PP_  (.D(net13),
    .DE(_026_),
    .Q(\b_to_a_mem[4][0] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[4][1]$_DFFE_PP_  (.D(net14),
    .DE(_026_),
    .Q(\b_to_a_mem[4][1] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[4][2]$_DFFE_PP_  (.D(net15),
    .DE(_026_),
    .Q(\b_to_a_mem[4][2] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[4][3]$_DFFE_PP_  (.D(net16),
    .DE(_026_),
    .Q(\b_to_a_mem[4][3] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[4][4]$_DFFE_PP_  (.D(net17),
    .DE(_026_),
    .Q(\b_to_a_mem[4][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[4][5]$_DFFE_PP_  (.D(net18),
    .DE(_026_),
    .Q(\b_to_a_mem[4][5] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[4][6]$_DFFE_PP_  (.D(net19),
    .DE(_026_),
    .Q(\b_to_a_mem[4][6] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[4][7]$_DFFE_PP_  (.D(net20),
    .DE(_026_),
    .Q(\b_to_a_mem[4][7] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[5][0]$_DFFE_PP_  (.D(net13),
    .DE(_027_),
    .Q(\b_to_a_mem[5][0] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[5][1]$_DFFE_PP_  (.D(net14),
    .DE(_027_),
    .Q(\b_to_a_mem[5][1] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[5][2]$_DFFE_PP_  (.D(net15),
    .DE(_027_),
    .Q(\b_to_a_mem[5][2] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[5][3]$_DFFE_PP_  (.D(net16),
    .DE(_027_),
    .Q(\b_to_a_mem[5][3] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[5][4]$_DFFE_PP_  (.D(net17),
    .DE(_027_),
    .Q(\b_to_a_mem[5][4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[5][5]$_DFFE_PP_  (.D(net18),
    .DE(_027_),
    .Q(\b_to_a_mem[5][5] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[5][6]$_DFFE_PP_  (.D(net19),
    .DE(_027_),
    .Q(\b_to_a_mem[5][6] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[5][7]$_DFFE_PP_  (.D(net20),
    .DE(_027_),
    .Q(\b_to_a_mem[5][7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[6][0]$_DFFE_PP_  (.D(net13),
    .DE(_028_),
    .Q(\b_to_a_mem[6][0] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[6][1]$_DFFE_PP_  (.D(net14),
    .DE(_028_),
    .Q(\b_to_a_mem[6][1] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[6][2]$_DFFE_PP_  (.D(net15),
    .DE(_028_),
    .Q(\b_to_a_mem[6][2] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[6][3]$_DFFE_PP_  (.D(net16),
    .DE(_028_),
    .Q(\b_to_a_mem[6][3] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[6][4]$_DFFE_PP_  (.D(net17),
    .DE(_028_),
    .Q(\b_to_a_mem[6][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[6][5]$_DFFE_PP_  (.D(net18),
    .DE(_028_),
    .Q(\b_to_a_mem[6][5] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[6][6]$_DFFE_PP_  (.D(net19),
    .DE(_028_),
    .Q(\b_to_a_mem[6][6] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[6][7]$_DFFE_PP_  (.D(net20),
    .DE(_028_),
    .Q(\b_to_a_mem[6][7] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[7][0]$_DFFE_PP_  (.D(net13),
    .DE(_029_),
    .Q(\b_to_a_mem[7][0] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[7][1]$_DFFE_PP_  (.D(net14),
    .DE(_029_),
    .Q(\b_to_a_mem[7][1] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[7][2]$_DFFE_PP_  (.D(net15),
    .DE(_029_),
    .Q(\b_to_a_mem[7][2] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[7][3]$_DFFE_PP_  (.D(net16),
    .DE(_029_),
    .Q(\b_to_a_mem[7][3] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[7][4]$_DFFE_PP_  (.D(net17),
    .DE(_029_),
    .Q(\b_to_a_mem[7][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[7][5]$_DFFE_PP_  (.D(net18),
    .DE(_029_),
    .Q(\b_to_a_mem[7][5] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[7][6]$_DFFE_PP_  (.D(net19),
    .DE(_029_),
    .Q(\b_to_a_mem[7][6] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[7][7]$_DFFE_PP_  (.D(net20),
    .DE(_029_),
    .Q(\b_to_a_mem[7][7] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[8][0]$_DFFE_PP_  (.D(net13),
    .DE(_030_),
    .Q(\b_to_a_mem[8][0] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[8][1]$_DFFE_PP_  (.D(net14),
    .DE(_030_),
    .Q(\b_to_a_mem[8][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[8][2]$_DFFE_PP_  (.D(net15),
    .DE(_030_),
    .Q(\b_to_a_mem[8][2] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[8][3]$_DFFE_PP_  (.D(net16),
    .DE(_030_),
    .Q(\b_to_a_mem[8][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[8][4]$_DFFE_PP_  (.D(net17),
    .DE(_030_),
    .Q(\b_to_a_mem[8][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[8][5]$_DFFE_PP_  (.D(net18),
    .DE(_030_),
    .Q(\b_to_a_mem[8][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[8][6]$_DFFE_PP_  (.D(net19),
    .DE(_030_),
    .Q(\b_to_a_mem[8][6] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[8][7]$_DFFE_PP_  (.D(net20),
    .DE(_030_),
    .Q(\b_to_a_mem[8][7] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[9][0]$_DFFE_PP_  (.D(net13),
    .DE(_031_),
    .Q(\b_to_a_mem[9][0] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[9][1]$_DFFE_PP_  (.D(net14),
    .DE(_031_),
    .Q(\b_to_a_mem[9][1] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[9][2]$_DFFE_PP_  (.D(net15),
    .DE(_031_),
    .Q(\b_to_a_mem[9][2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[9][3]$_DFFE_PP_  (.D(net16),
    .DE(_031_),
    .Q(\b_to_a_mem[9][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[9][4]$_DFFE_PP_  (.D(net17),
    .DE(_031_),
    .Q(\b_to_a_mem[9][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[9][5]$_DFFE_PP_  (.D(net18),
    .DE(_031_),
    .Q(\b_to_a_mem[9][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[9][6]$_DFFE_PP_  (.D(net19),
    .DE(_031_),
    .Q(\b_to_a_mem[9][6] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \b_to_a_mem[9][7]$_DFFE_PP_  (.D(net20),
    .DE(_031_),
    .Q(\b_to_a_mem[9][7] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_wr_ptr[0]$_DFFE_PN0P_  (.D(_069_),
    .Q(\b_wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \b_wr_ptr[1]$_DFFE_PN0P_  (.D(_070_),
    .Q(\b_wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \b_wr_ptr[2]$_DFFE_PN0P_  (.D(_071_),
    .Q(\b_wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \b_wr_ptr[3]$_DFFE_PN0P_  (.D(_072_),
    .Q(\b_wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_wr_ptr[4]$_DFFE_PN0P_  (.D(_073_),
    .Q(\b_wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__buf_12 hold1 (.A(net56),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_274 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(a_rd_en),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(net69),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_8 input3 (.A(net58),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input4 (.A(net67),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input5 (.A(net64),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input6 (.A(net57),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input7 (.A(a_wr_data[5]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input8 (.A(net68),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input9 (.A(net60),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(a_wr_en),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(b_rd_en),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input12 (.A(net59),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input13 (.A(net62),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input14 (.A(b_wr_data[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input15 (.A(net65),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input16 (.A(b_wr_data[4]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input17 (.A(net66),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input18 (.A(net63),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input19 (.A(net61),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(b_wr_en),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(a_almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(a_almost_full));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(a_empty));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(a_full));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(a_rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(a_rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(a_rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(a_rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(a_rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(a_rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(a_rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(a_rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(a_to_b_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(a_to_b_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net36),
    .X(a_to_b_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net37),
    .X(a_to_b_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net38),
    .X(a_to_b_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net39),
    .X(b_almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net40),
    .X(b_almost_full));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net41),
    .X(b_empty));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net42),
    .X(b_full));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net43),
    .X(b_rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net44),
    .X(b_rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net45),
    .X(b_rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net46),
    .X(b_rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net47),
    .X(b_rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net48),
    .X(b_rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net49),
    .X(b_rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net50),
    .X(b_rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net51),
    .X(b_to_a_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net52),
    .X(b_to_a_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net53),
    .X(b_to_a_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net54),
    .X(b_to_a_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net55),
    .X(b_to_a_count[4]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload1 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload2 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinv_2 clkload3 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload4 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload5 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__bufinv_16 clkload6 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkinv_2 clkload7 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkinv_2 clkload8 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload9 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__bufinv_16 clkload10 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload11 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload12 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkinv_4 clkload13 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__bufinv_16 clkload15 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__bufinv_16 clkload16 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_1 clkload17 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload18 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinv_2 clkload19 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload20 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_2 clkload21 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinv_2 clkload22 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkinv_1 clkload23 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(a_wr_data[4]),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(a_wr_data[1]),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(b_wr_data[0]),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(a_wr_data[7]),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(b_wr_data[7]),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(b_wr_data[1]),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(b_wr_data[6]),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(a_wr_data[3]),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(b_wr_data[3]),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(b_wr_data[5]),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(a_wr_data[2]),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(a_wr_data[6]),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(a_wr_data[0]),
    .X(net69));
 sky130_fd_sc_hd__fill_4 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_299 ();
endmodule
