module cordic (clk,
    done,
    rst_n,
    start,
    x_in,
    x_out,
    y_in,
    y_out,
    z_in,
    z_out);
 input clk;
 output done;
 input rst_n;
 input start;
 input [15:0] x_in;
 output [15:0] x_out;
 input [15:0] y_in;
 output [15:0] y_out;
 input [15:0] z_in;
 output [15:0] z_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire \iteration[0] ;
 wire \iteration[1] ;
 wire \iteration[2] ;
 wire \iteration[3] ;
 wire \next_state[1] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \x[0] ;
 wire \x[10] ;
 wire \x[11] ;
 wire \x[12] ;
 wire \x[13] ;
 wire \x[14] ;
 wire \x[15] ;
 wire \x[1] ;
 wire \x[2] ;
 wire \x[3] ;
 wire \x[4] ;
 wire \x[5] ;
 wire \x[6] ;
 wire \x[7] ;
 wire \x[8] ;
 wire \x[9] ;
 wire \y[0] ;
 wire \y[10] ;
 wire \y[11] ;
 wire \y[12] ;
 wire \y[13] ;
 wire \y[14] ;
 wire \y[15] ;
 wire \y[1] ;
 wire \y[2] ;
 wire \y[3] ;
 wire \y[4] ;
 wire \y[5] ;
 wire \y[6] ;
 wire \y[7] ;
 wire \y[8] ;
 wire \y[9] ;
 wire \z[0] ;
 wire \z[10] ;
 wire \z[11] ;
 wire \z[12] ;
 wire \z[13] ;
 wire \z[14] ;
 wire \z[15] ;
 wire \z[1] ;
 wire \z[2] ;
 wire \z[3] ;
 wire \z[4] ;
 wire \z[5] ;
 wire \z[6] ;
 wire \z[7] ;
 wire \z[8] ;
 wire \z[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;

 sky130_fd_sc_hd__buf_6 _0918_ (.A(\iteration[1] ),
    .X(_0266_));
 sky130_fd_sc_hd__buf_4 _0919_ (.A(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__buf_4 _0920_ (.A(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__clkinvlp_4 _0921_ (.A(_0268_),
    .Y(_0764_));
 sky130_fd_sc_hd__buf_6 _0922_ (.A(\iteration[3] ),
    .X(_0269_));
 sky130_fd_sc_hd__clkbuf_4 _0923_ (.A(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__buf_4 _0924_ (.A(\iteration[2] ),
    .X(_0271_));
 sky130_fd_sc_hd__buf_4 _0925_ (.A(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_1 _0926_ (.A(_0272_),
    .B(_0268_),
    .Y(_0273_));
 sky130_fd_sc_hd__and2_0 _0927_ (.A(_0272_),
    .B(_0775_),
    .X(_0274_));
 sky130_fd_sc_hd__nand2b_1 _0928_ (.A_N(_0766_),
    .B(_0269_),
    .Y(_0275_));
 sky130_fd_sc_hd__o31ai_2 _0929_ (.A1(_0270_),
    .A2(_0273_),
    .A3(_0274_),
    .B1(_0275_),
    .Y(_0746_));
 sky130_fd_sc_hd__inv_1 _0930_ (.A(_0746_),
    .Y(_0749_));
 sky130_fd_sc_hd__buf_8 _0931_ (.A(\iteration[0] ),
    .X(_0276_));
 sky130_fd_sc_hd__buf_6 _0932_ (.A(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__buf_4 _0933_ (.A(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__clkinv_4 _0934_ (.A(_0278_),
    .Y(_0763_));
 sky130_fd_sc_hd__buf_4 _0935_ (.A(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__a211oi_1 _0936_ (.A1(_0279_),
    .A2(_0268_),
    .B1(_0273_),
    .C1(_0270_),
    .Y(_0280_));
 sky130_fd_sc_hd__a21oi_1 _0937_ (.A1(_0270_),
    .A2(_0771_),
    .B1(_0280_),
    .Y(_0748_));
 sky130_fd_sc_hd__clkbuf_4 _0938_ (.A(_0270_),
    .X(_0281_));
 sky130_fd_sc_hd__nand2_1 _0939_ (.A(_0269_),
    .B(_0763_),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_1 _0940_ (.A(\iteration[3] ),
    .Y(_0283_));
 sky130_fd_sc_hd__buf_4 _0941_ (.A(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__buf_4 _0942_ (.A(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__buf_4 _0943_ (.A(_0271_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2i_1 _0944_ (.A0(_0771_),
    .A1(_0767_),
    .S(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__nand2_1 _0945_ (.A(_0285_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__o32ai_4 _0946_ (.A1(_0771_),
    .A2(_0767_),
    .A3(_0282_),
    .B1(_0288_),
    .B2(_0773_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand2_1 _0947_ (.A(_0750_),
    .B(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__clkinv_2 _0948_ (.A(_0271_),
    .Y(_0291_));
 sky130_fd_sc_hd__buf_4 _0949_ (.A(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__nand2_1 _0950_ (.A(_0292_),
    .B(_0766_),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2_1 _0951_ (.A(_0286_),
    .B(_0771_),
    .Y(_0294_));
 sky130_fd_sc_hd__nor2_1 _0952_ (.A(_0285_),
    .B(_0767_),
    .Y(_0295_));
 sky130_fd_sc_hd__a31oi_2 _0953_ (.A1(_0285_),
    .A2(_0293_),
    .A3(_0294_),
    .B1(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__mux2i_1 _0954_ (.A0(_0268_),
    .A1(_0779_),
    .S(_0286_),
    .Y(_0297_));
 sky130_fd_sc_hd__nor2_1 _0955_ (.A(_0270_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__a21oi_2 _0956_ (.A1(_0270_),
    .A2(_0775_),
    .B1(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__nor3b_2 _0957_ (.A(_0290_),
    .B(_0296_),
    .C_N(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__buf_4 _0958_ (.A(\z[15] ),
    .X(_0301_));
 sky130_fd_sc_hd__buf_4 _0959_ (.A(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__a21oi_1 _0960_ (.A1(_0281_),
    .A2(_0300_),
    .B1(_0302_),
    .Y(_0808_));
 sky130_fd_sc_hd__mux4_4 _0961_ (.A0(\x[12] ),
    .A1(\x[13] ),
    .A2(\x[14] ),
    .A3(\x[15] ),
    .S0(_0276_),
    .S1(_0266_),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_4 _0962_ (.A(_0266_),
    .X(_0304_));
 sky130_fd_sc_hd__mux4_1 _0963_ (.A0(\x[4] ),
    .A1(\x[5] ),
    .A2(\x[6] ),
    .A3(\x[7] ),
    .S0(_0276_),
    .S1(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _0964_ (.A0(_0303_),
    .A1(_0305_),
    .S(_0283_),
    .X(_0306_));
 sky130_fd_sc_hd__buf_4 _0965_ (.A(_0266_),
    .X(_0307_));
 sky130_fd_sc_hd__mux4_1 _0966_ (.A0(\x[0] ),
    .A1(\x[1] ),
    .A2(\x[2] ),
    .A3(\x[3] ),
    .S0(_0277_),
    .S1(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__nor2_2 _0967_ (.A(_0271_),
    .B(_0269_),
    .Y(_0309_));
 sky130_fd_sc_hd__nor2b_2 _0968_ (.A(_0271_),
    .B_N(\iteration[3] ),
    .Y(_0310_));
 sky130_fd_sc_hd__mux4_2 _0969_ (.A0(\x[8] ),
    .A1(\x[9] ),
    .A2(\x[10] ),
    .A3(\x[11] ),
    .S0(_0276_),
    .S1(_0266_),
    .X(_0311_));
 sky130_fd_sc_hd__a22o_1 _0970_ (.A1(_0308_),
    .A2(_0309_),
    .B1(_0310_),
    .B2(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__a21oi_4 _0971_ (.A1(_0272_),
    .A2(_0306_),
    .B1(_0312_),
    .Y(_0816_));
 sky130_fd_sc_hd__inv_1 _0972_ (.A(_0816_),
    .Y(_0812_));
 sky130_fd_sc_hd__clkbuf_4 _0973_ (.A(_0286_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2i_2 _0974_ (.A0(\x[14] ),
    .A1(\x[15] ),
    .S(_0276_),
    .Y(_0314_));
 sky130_fd_sc_hd__or2_2 _0975_ (.A(_0266_),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2i_4 _0976_ (.A0(\x[7] ),
    .A1(\x[9] ),
    .S(_0266_),
    .Y(_0316_));
 sky130_fd_sc_hd__nor2b_4 _0977_ (.A(\iteration[3] ),
    .B_N(_0277_),
    .Y(_0317_));
 sky130_fd_sc_hd__mux2_1 _0978_ (.A0(\x[6] ),
    .A1(\x[8] ),
    .S(_0266_),
    .X(_0318_));
 sky130_fd_sc_hd__nor3_1 _0979_ (.A(\iteration[3] ),
    .B(_0277_),
    .C(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__a221oi_4 _0980_ (.A1(\iteration[3] ),
    .A2(_0315_),
    .B1(_0316_),
    .B2(_0317_),
    .C1(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__mux4_4 _0981_ (.A0(\x[10] ),
    .A1(\x[11] ),
    .A2(\x[12] ),
    .A3(\x[13] ),
    .S0(_0276_),
    .S1(_0266_),
    .X(_0321_));
 sky130_fd_sc_hd__nand2_1 _0982_ (.A(_0281_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__mux4_1 _0983_ (.A0(\x[2] ),
    .A1(\x[3] ),
    .A2(\x[4] ),
    .A3(\x[5] ),
    .S0(_0276_),
    .S1(_0304_),
    .X(_0323_));
 sky130_fd_sc_hd__nand2_1 _0984_ (.A(_0285_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21oi_1 _0985_ (.A1(_0322_),
    .A2(_0324_),
    .B1(_0313_),
    .Y(_0325_));
 sky130_fd_sc_hd__a21oi_1 _0986_ (.A1(_0313_),
    .A2(_0320_),
    .B1(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__buf_4 _0987_ (.A(_0301_),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_1 _0988_ (.A(_0327_),
    .B(_0817_),
    .Y(_0328_));
 sky130_fd_sc_hd__xor2_1 _0989_ (.A(_0326_),
    .B(_0328_),
    .X(_0821_));
 sky130_fd_sc_hd__mux4_4 _0990_ (.A0(\x[11] ),
    .A1(\x[12] ),
    .A2(\x[13] ),
    .A3(\x[14] ),
    .S0(_0276_),
    .S1(_0307_),
    .X(_0329_));
 sky130_fd_sc_hd__mux4_1 _0991_ (.A0(\x[3] ),
    .A1(\x[4] ),
    .A2(\x[5] ),
    .A3(\x[6] ),
    .S0(_0277_),
    .S1(_0267_),
    .X(_0330_));
 sky130_fd_sc_hd__a22oi_2 _0992_ (.A1(_0310_),
    .A2(_0329_),
    .B1(_0330_),
    .B2(_0309_),
    .Y(_0331_));
 sky130_fd_sc_hd__nand2b_1 _0993_ (.A_N(_0304_),
    .B(\x[15] ),
    .Y(_0332_));
 sky130_fd_sc_hd__a21oi_1 _0994_ (.A1(_0269_),
    .A2(_0332_),
    .B1(_0278_),
    .Y(_0333_));
 sky130_fd_sc_hd__mux2i_1 _0995_ (.A0(\x[8] ),
    .A1(\x[10] ),
    .S(_0307_),
    .Y(_0334_));
 sky130_fd_sc_hd__nor2_1 _0996_ (.A(_0269_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nor2_4 _0997_ (.A(_0269_),
    .B(_0277_),
    .Y(_0336_));
 sky130_fd_sc_hd__a21oi_1 _0998_ (.A1(_0316_),
    .A2(_0336_),
    .B1(_0291_),
    .Y(_0337_));
 sky130_fd_sc_hd__o21ai_2 _0999_ (.A1(_0333_),
    .A2(_0335_),
    .B1(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_2 _1000_ (.A(_0331_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(\x[13] ),
    .A1(\x[15] ),
    .S(\iteration[1] ),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(\x[5] ),
    .A1(\x[7] ),
    .S(net104),
    .X(_0341_));
 sky130_fd_sc_hd__nor2b_1 _1003_ (.A(_0266_),
    .B_N(\x[14] ),
    .Y(_0342_));
 sky130_fd_sc_hd__mux4_1 _1004_ (.A0(_0340_),
    .A1(_0341_),
    .A2(_0342_),
    .A3(_0318_),
    .S0(_0283_),
    .S1(_0278_),
    .X(_0343_));
 sky130_fd_sc_hd__mux4_1 _1005_ (.A0(\x[9] ),
    .A1(\x[10] ),
    .A2(\x[11] ),
    .A3(\x[12] ),
    .S0(_0277_),
    .S1(_0307_),
    .X(_0344_));
 sky130_fd_sc_hd__mux4_1 _1006_ (.A0(\x[1] ),
    .A1(\x[2] ),
    .A2(\x[3] ),
    .A3(\x[4] ),
    .S0(_0277_),
    .S1(_0307_),
    .X(_0345_));
 sky130_fd_sc_hd__a22o_1 _1007_ (.A1(_0310_),
    .A2(_0344_),
    .B1(_0345_),
    .B2(_0309_),
    .X(_0346_));
 sky130_fd_sc_hd__a21oi_2 _1008_ (.A1(_0272_),
    .A2(_0343_),
    .B1(_0346_),
    .Y(_0815_));
 sky130_fd_sc_hd__buf_4 _1009_ (.A(_0301_),
    .X(_0347_));
 sky130_fd_sc_hd__a31oi_1 _1010_ (.A1(_0816_),
    .A2(_0326_),
    .A3(_0815_),
    .B1(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__xnor2_1 _1011_ (.A(_0339_),
    .B(_0348_),
    .Y(_0824_));
 sky130_fd_sc_hd__inv_1 _1012_ (.A(_0813_),
    .Y(_0737_));
 sky130_fd_sc_hd__buf_4 _1013_ (.A(_0301_),
    .X(_0349_));
 sky130_fd_sc_hd__a41oi_1 _1014_ (.A1(_0817_),
    .A2(_0326_),
    .A3(_0331_),
    .A4(_0338_),
    .B1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__and3_1 _1015_ (.A(_0271_),
    .B(_0284_),
    .C(_0311_),
    .X(_0351_));
 sky130_fd_sc_hd__a21oi_1 _1016_ (.A1(_0292_),
    .A2(_0306_),
    .B1(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__xor2_1 _1017_ (.A(_0350_),
    .B(_0352_),
    .X(_0827_));
 sky130_fd_sc_hd__nand2_2 _1018_ (.A(_0271_),
    .B(_0284_),
    .Y(_0353_));
 sky130_fd_sc_hd__mux2i_1 _1019_ (.A0(\x[9] ),
    .A1(\x[11] ),
    .S(_0307_),
    .Y(_0354_));
 sky130_fd_sc_hd__mux2i_1 _1020_ (.A0(\x[10] ),
    .A1(\x[12] ),
    .S(_0307_),
    .Y(_0355_));
 sky130_fd_sc_hd__mux2_2 _1021_ (.A0(_0354_),
    .A1(_0355_),
    .S(_0277_),
    .X(_0356_));
 sky130_fd_sc_hd__nand2_1 _1022_ (.A(_0291_),
    .B(_0343_),
    .Y(_0357_));
 sky130_fd_sc_hd__o21ai_2 _1023_ (.A1(_0353_),
    .A2(_0356_),
    .B1(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_1 _1024_ (.A(_0816_),
    .B(_0815_),
    .Y(_0359_));
 sky130_fd_sc_hd__o21ai_0 _1025_ (.A1(_0305_),
    .A2(_0323_),
    .B1(_0309_),
    .Y(_0360_));
 sky130_fd_sc_hd__o21ai_0 _1026_ (.A1(_0303_),
    .A2(_0321_),
    .B1(_0310_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_1 _1027_ (.A(_0360_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__a211o_1 _1028_ (.A1(_0271_),
    .A2(_0320_),
    .B1(_0351_),
    .C1(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__clkinv_4 _1029_ (.A(_0301_),
    .Y(_0364_));
 sky130_fd_sc_hd__o31ai_1 _1030_ (.A1(_0339_),
    .A2(_0359_),
    .A3(_0363_),
    .B1(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__xor2_1 _1031_ (.A(_0358_),
    .B(_0365_),
    .X(_0830_));
 sky130_fd_sc_hd__nor2_4 _1032_ (.A(_0291_),
    .B(_0269_),
    .Y(_0366_));
 sky130_fd_sc_hd__a22oi_2 _1033_ (.A1(_0292_),
    .A2(_0320_),
    .B1(_0321_),
    .B2(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__or4b_1 _1034_ (.A(_0339_),
    .B(_0358_),
    .C(_0363_),
    .D_N(_0817_),
    .X(_0368_));
 sky130_fd_sc_hd__nand2_1 _1035_ (.A(_0364_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__xnor2_1 _1036_ (.A(_0367_),
    .B(_0369_),
    .Y(_0833_));
 sky130_fd_sc_hd__a21oi_1 _1037_ (.A1(_0316_),
    .A2(_0336_),
    .B1(_0272_),
    .Y(_0370_));
 sky130_fd_sc_hd__o21ai_1 _1038_ (.A1(_0333_),
    .A2(_0335_),
    .B1(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_1 _1039_ (.A(_0366_),
    .B(_0329_),
    .Y(_0372_));
 sky130_fd_sc_hd__nand2_2 _1040_ (.A(_0371_),
    .B(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__a2111o_1 _1041_ (.A1(_0366_),
    .A2(_0321_),
    .B1(_0351_),
    .C1(_0362_),
    .D1(_0320_),
    .X(_0374_));
 sky130_fd_sc_hd__nor4_4 _1042_ (.A(_0339_),
    .B(_0359_),
    .C(_0358_),
    .D(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__nor2_1 _1043_ (.A(_0302_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__xnor2_1 _1044_ (.A(_0373_),
    .B(_0376_),
    .Y(_0836_));
 sky130_fd_sc_hd__buf_4 _1045_ (.A(_0309_),
    .X(_0377_));
 sky130_fd_sc_hd__a22oi_2 _1046_ (.A1(net101),
    .A2(_0366_),
    .B1(_0311_),
    .B2(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__inv_1 _1047_ (.A(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2b_1 _1048_ (.A_N(_0368_),
    .B(_0367_),
    .Y(_0380_));
 sky130_fd_sc_hd__nor2_1 _1049_ (.A(_0373_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__nor2_1 _1050_ (.A(_0302_),
    .B(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__xnor2_1 _1051_ (.A(_0379_),
    .B(_0382_),
    .Y(_0839_));
 sky130_fd_sc_hd__mux2i_1 _1052_ (.A0(_0340_),
    .A1(_0342_),
    .S(_0278_),
    .Y(_0383_));
 sky130_fd_sc_hd__mux2i_2 _1053_ (.A0(_0383_),
    .A1(_0356_),
    .S(_0291_),
    .Y(_0384_));
 sky130_fd_sc_hd__and2_1 _1054_ (.A(_0285_),
    .B(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_1 _1055_ (.A(_0373_),
    .B(_0379_),
    .Y(_0386_));
 sky130_fd_sc_hd__a21oi_1 _1056_ (.A1(_0375_),
    .A2(_0386_),
    .B1(_0327_),
    .Y(_0387_));
 sky130_fd_sc_hd__xnor2_1 _1057_ (.A(_0385_),
    .B(_0387_),
    .Y(_0842_));
 sky130_fd_sc_hd__nor2_1 _1058_ (.A(_0268_),
    .B(_0314_),
    .Y(_0388_));
 sky130_fd_sc_hd__mux2i_1 _1059_ (.A0(_0388_),
    .A1(_0321_),
    .S(_0292_),
    .Y(_0389_));
 sky130_fd_sc_hd__nor2_1 _1060_ (.A(_0270_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__o41a_1 _1061_ (.A1(_0373_),
    .A2(_0379_),
    .A3(_0380_),
    .A4(_0385_),
    .B1(_0364_),
    .X(_0391_));
 sky130_fd_sc_hd__xnor2_1 _1062_ (.A(_0390_),
    .B(_0391_),
    .Y(_0845_));
 sky130_fd_sc_hd__nand2_1 _1063_ (.A(_0292_),
    .B(_0329_),
    .Y(_0392_));
 sky130_fd_sc_hd__nor2_1 _1064_ (.A(_0279_),
    .B(_0268_),
    .Y(_0393_));
 sky130_fd_sc_hd__nand3_2 _1065_ (.A(_0286_),
    .B(\x[15] ),
    .C(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__a21o_2 _1066_ (.A1(_0392_),
    .A2(_0394_),
    .B1(_0270_),
    .X(_0395_));
 sky130_fd_sc_hd__nor4_2 _1067_ (.A(_0373_),
    .B(_0379_),
    .C(_0385_),
    .D(_0390_),
    .Y(_0396_));
 sky130_fd_sc_hd__a21oi_1 _1068_ (.A1(_0375_),
    .A2(_0396_),
    .B1(_0301_),
    .Y(_0397_));
 sky130_fd_sc_hd__xor2_1 _1069_ (.A(_0395_),
    .B(_0397_),
    .X(_0848_));
 sky130_fd_sc_hd__nand2_1 _1070_ (.A(_0395_),
    .B(_0396_),
    .Y(_0398_));
 sky130_fd_sc_hd__nor2_2 _1071_ (.A(_0380_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__nor2_1 _1072_ (.A(_0347_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__buf_2 _1073_ (.A(_0377_),
    .X(_0401_));
 sky130_fd_sc_hd__nand2_1 _1074_ (.A(net102),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__xor2_1 _1075_ (.A(_0400_),
    .B(_0402_),
    .X(_0851_));
 sky130_fd_sc_hd__nand2_1 _1076_ (.A(_0763_),
    .B(_0340_),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _1077_ (.A(_0279_),
    .B(_0342_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand2_1 _1078_ (.A(_0403_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__nand2_1 _1079_ (.A(_0364_),
    .B(net102),
    .Y(_0406_));
 sky130_fd_sc_hd__nor2b_1 _1080_ (.A(net102),
    .B_N(_0395_),
    .Y(_0407_));
 sky130_fd_sc_hd__o21ai_0 _1081_ (.A1(_0349_),
    .A2(_0407_),
    .B1(_0405_),
    .Y(_0408_));
 sky130_fd_sc_hd__o22ai_1 _1082_ (.A1(_0405_),
    .A2(_0406_),
    .B1(_0408_),
    .B2(_0397_),
    .Y(_0409_));
 sky130_fd_sc_hd__nor2_1 _1083_ (.A(_0349_),
    .B(_0395_),
    .Y(_0410_));
 sky130_fd_sc_hd__nor2_1 _1084_ (.A(_0397_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__a21oi_1 _1085_ (.A1(_0401_),
    .A2(_0405_),
    .B1(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__a21oi_1 _1086_ (.A1(_0401_),
    .A2(_0409_),
    .B1(_0412_),
    .Y(_0854_));
 sky130_fd_sc_hd__nor2_1 _1087_ (.A(net102),
    .B(_0405_),
    .Y(_0413_));
 sky130_fd_sc_hd__a21oi_1 _1088_ (.A1(_0399_),
    .A2(_0413_),
    .B1(_0349_),
    .Y(_0414_));
 sky130_fd_sc_hd__o21ai_0 _1089_ (.A1(_0301_),
    .A2(_0413_),
    .B1(_0315_),
    .Y(_0415_));
 sky130_fd_sc_hd__a2bb2oi_1 _1090_ (.A1_N(_0349_),
    .A2_N(_0399_),
    .B1(_0415_),
    .B2(_0401_),
    .Y(_0416_));
 sky130_fd_sc_hd__a31o_1 _1091_ (.A1(_0401_),
    .A2(_0388_),
    .A3(_0414_),
    .B1(_0416_),
    .X(_0857_));
 sky130_fd_sc_hd__clkbuf_4 _1092_ (.A(_0313_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2i_4 _1093_ (.A0(\y[1] ),
    .A1(\y[3] ),
    .S(_0267_),
    .Y(_0418_));
 sky130_fd_sc_hd__mux2i_2 _1094_ (.A0(\y[0] ),
    .A1(\y[2] ),
    .S(_0268_),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _1095_ (.A(_0269_),
    .B(_0278_),
    .Y(_0420_));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(\y[9] ),
    .A1(\y[11] ),
    .S(_0304_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_2 _1097_ (.A0(\y[8] ),
    .A1(\y[10] ),
    .S(_0304_),
    .X(_0422_));
 sky130_fd_sc_hd__o22ai_2 _1098_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0422_),
    .B2(_0282_),
    .Y(_0423_));
 sky130_fd_sc_hd__a221oi_4 _1099_ (.A1(_0317_),
    .A2(_0418_),
    .B1(_0419_),
    .B2(_0336_),
    .C1(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__clkbuf_4 _1100_ (.A(\y[15] ),
    .X(_0425_));
 sky130_fd_sc_hd__mux4_4 _1101_ (.A0(\y[12] ),
    .A1(\y[13] ),
    .A2(\y[14] ),
    .A3(_0425_),
    .S0(_0276_),
    .S1(_0304_),
    .X(_0426_));
 sky130_fd_sc_hd__mux4_2 _1102_ (.A0(\y[4] ),
    .A1(\y[5] ),
    .A2(\y[6] ),
    .A3(\y[7] ),
    .S0(_0276_),
    .S1(_0307_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2i_4 _1103_ (.A0(_0426_),
    .A1(_0427_),
    .S(_0284_),
    .Y(_0428_));
 sky130_fd_sc_hd__nand2_1 _1104_ (.A(_0417_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__o21ai_2 _1105_ (.A1(_0417_),
    .A2(_0424_),
    .B1(_0429_),
    .Y(_0863_));
 sky130_fd_sc_hd__inv_1 _1106_ (.A(_0863_),
    .Y(_0860_));
 sky130_fd_sc_hd__mux2i_1 _1107_ (.A0(\y[13] ),
    .A1(_0425_),
    .S(_0307_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand3b_1 _1108_ (.A_N(_0267_),
    .B(\y[14] ),
    .C(_0278_),
    .Y(_0431_));
 sky130_fd_sc_hd__o21ai_2 _1109_ (.A1(_0278_),
    .A2(_0430_),
    .B1(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__mux2i_1 _1110_ (.A0(\y[5] ),
    .A1(\y[7] ),
    .S(_0267_),
    .Y(_0433_));
 sky130_fd_sc_hd__mux2i_2 _1111_ (.A0(\y[6] ),
    .A1(\y[8] ),
    .S(_0267_),
    .Y(_0434_));
 sky130_fd_sc_hd__a22oi_2 _1112_ (.A1(_0336_),
    .A2(_0433_),
    .B1(_0434_),
    .B2(_0317_),
    .Y(_0435_));
 sky130_fd_sc_hd__o21ai_2 _1113_ (.A1(_0284_),
    .A2(_0432_),
    .B1(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__mux2_1 _1114_ (.A0(\y[2] ),
    .A1(\y[4] ),
    .S(_0304_),
    .X(_0437_));
 sky130_fd_sc_hd__nand2_1 _1115_ (.A(_0763_),
    .B(_0418_),
    .Y(_0438_));
 sky130_fd_sc_hd__o21ai_1 _1116_ (.A1(_0763_),
    .A2(_0437_),
    .B1(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__mux2_2 _1117_ (.A0(\y[10] ),
    .A1(\y[12] ),
    .S(_0304_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _1118_ (.A0(_0421_),
    .A1(_0440_),
    .S(_0278_),
    .X(_0441_));
 sky130_fd_sc_hd__nor2_1 _1119_ (.A(_0284_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__a21oi_2 _1120_ (.A1(_0284_),
    .A2(_0439_),
    .B1(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nor2_1 _1121_ (.A(_0417_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__a21oi_1 _1122_ (.A1(_0417_),
    .A2(_0436_),
    .B1(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__mux2_1 _1123_ (.A0(_0866_),
    .A1(_0445_),
    .S(_0349_),
    .X(_0867_));
 sky130_fd_sc_hd__inv_1 _1124_ (.A(_0867_),
    .Y(_0743_));
 sky130_fd_sc_hd__inv_1 _1125_ (.A(\x[1] ),
    .Y(_0741_));
 sky130_fd_sc_hd__inv_1 _1126_ (.A(_0861_),
    .Y(_0742_));
 sky130_fd_sc_hd__inv_1 _1127_ (.A(\y[0] ),
    .Y(_0811_));
 sky130_fd_sc_hd__mux2_1 _1128_ (.A0(_0432_),
    .A1(_0441_),
    .S(_0292_),
    .X(_0446_));
 sky130_fd_sc_hd__nand2_1 _1129_ (.A(_0285_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__mux2_2 _1130_ (.A0(\y[11] ),
    .A1(\y[13] ),
    .S(_0304_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _1131_ (.A0(\y[3] ),
    .A1(\y[5] ),
    .S(_0307_),
    .X(_0449_));
 sky130_fd_sc_hd__mux4_4 _1132_ (.A0(_0440_),
    .A1(_0437_),
    .A2(_0448_),
    .A3(_0449_),
    .S0(_0284_),
    .S1(_0279_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2i_1 _1133_ (.A0(\y[14] ),
    .A1(_0425_),
    .S(_0277_),
    .Y(_0451_));
 sky130_fd_sc_hd__nor2_1 _1134_ (.A(_0267_),
    .B(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__mux2i_2 _1135_ (.A0(\y[7] ),
    .A1(\y[9] ),
    .S(_0267_),
    .Y(_0453_));
 sky130_fd_sc_hd__a22oi_2 _1136_ (.A1(_0336_),
    .A2(_0434_),
    .B1(_0453_),
    .B2(_0317_),
    .Y(_0454_));
 sky130_fd_sc_hd__o21ai_2 _1137_ (.A1(_0284_),
    .A2(_0452_),
    .B1(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__nand4_1 _1138_ (.A(_0313_),
    .B(_0428_),
    .C(_0436_),
    .D(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__o41ai_4 _1139_ (.A1(_0286_),
    .A2(_0424_),
    .A3(_0443_),
    .A4(_0450_),
    .B1(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _1140_ (.A(_0292_),
    .B(_0285_),
    .Y(_0458_));
 sky130_fd_sc_hd__mux2i_4 _1141_ (.A0(_0421_),
    .A1(_0422_),
    .S(_0763_),
    .Y(_0459_));
 sky130_fd_sc_hd__nand2_1 _1142_ (.A(_0366_),
    .B(_0426_),
    .Y(_0460_));
 sky130_fd_sc_hd__o21ai_2 _1143_ (.A1(_0458_),
    .A2(_0459_),
    .B1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nand2b_1 _1144_ (.A_N(_0267_),
    .B(_0425_),
    .Y(_0462_));
 sky130_fd_sc_hd__a21oi_1 _1145_ (.A1(_0269_),
    .A2(_0462_),
    .B1(_0279_),
    .Y(_0463_));
 sky130_fd_sc_hd__and2_0 _1146_ (.A(_0284_),
    .B(_0422_),
    .X(_0464_));
 sky130_fd_sc_hd__nand2_1 _1147_ (.A(_0336_),
    .B(_0453_),
    .Y(_0465_));
 sky130_fd_sc_hd__o21ai_0 _1148_ (.A1(_0463_),
    .A2(_0464_),
    .B1(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__mux2_1 _1149_ (.A0(\y[12] ),
    .A1(\y[14] ),
    .S(_0304_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_2 _1150_ (.A0(_0467_),
    .A1(_0448_),
    .S(_0763_),
    .X(_0468_));
 sky130_fd_sc_hd__nand2_1 _1151_ (.A(_0366_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__o21ai_1 _1152_ (.A1(_0272_),
    .A2(_0466_),
    .B1(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__mux2i_4 _1153_ (.A0(_0440_),
    .A1(_0448_),
    .S(_0279_),
    .Y(_0471_));
 sky130_fd_sc_hd__o22ai_2 _1154_ (.A1(_0286_),
    .A2(_0455_),
    .B1(_0471_),
    .B2(_0353_),
    .Y(_0472_));
 sky130_fd_sc_hd__o22a_1 _1155_ (.A1(_0272_),
    .A2(_0428_),
    .B1(_0459_),
    .B2(_0353_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2i_1 _1156_ (.A0(\y[4] ),
    .A1(\y[6] ),
    .S(_0267_),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_1 _1157_ (.A(_0279_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__o211ai_4 _1158_ (.A1(_0279_),
    .A2(_0449_),
    .B1(_0475_),
    .C1(_0377_),
    .Y(_0476_));
 sky130_fd_sc_hd__o211ai_2 _1159_ (.A1(_0463_),
    .A2(_0464_),
    .B1(_0465_),
    .C1(_0272_),
    .Y(_0477_));
 sky130_fd_sc_hd__nand2_1 _1160_ (.A(_0310_),
    .B(_0468_),
    .Y(_0478_));
 sky130_fd_sc_hd__nand4_1 _1161_ (.A(_0473_),
    .B(_0476_),
    .C(_0477_),
    .D(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand2_1 _1162_ (.A(_0366_),
    .B(_0441_),
    .Y(_0480_));
 sky130_fd_sc_hd__o21ai_2 _1163_ (.A1(_0272_),
    .A2(_0436_),
    .B1(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__nor4_2 _1164_ (.A(_0470_),
    .B(_0472_),
    .C(_0479_),
    .D(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__and2b_1 _1165_ (.A_N(_0461_),
    .B(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__a21oi_1 _1166_ (.A1(_0457_),
    .A2(_0483_),
    .B1(_0327_),
    .Y(_0484_));
 sky130_fd_sc_hd__xnor2_1 _1167_ (.A(_0447_),
    .B(_0484_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand2_1 _1168_ (.A(_0377_),
    .B(_0426_),
    .Y(_0485_));
 sky130_fd_sc_hd__nor2_1 _1169_ (.A(_0286_),
    .B(_0450_),
    .Y(_0486_));
 sky130_fd_sc_hd__a21oi_1 _1170_ (.A1(_0286_),
    .A2(_0455_),
    .B1(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__nor2b_2 _1171_ (.A(_0487_),
    .B_N(_0865_),
    .Y(_0488_));
 sky130_fd_sc_hd__and3_1 _1172_ (.A(_0447_),
    .B(_0483_),
    .C(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nor2b_1 _1173_ (.A(_0278_),
    .B_N(\y[14] ),
    .Y(_0490_));
 sky130_fd_sc_hd__o21ai_0 _1174_ (.A1(_0425_),
    .A2(_0490_),
    .B1(_0764_),
    .Y(_0491_));
 sky130_fd_sc_hd__mux2i_1 _1175_ (.A0(_0467_),
    .A1(_0440_),
    .S(_0763_),
    .Y(_0492_));
 sky130_fd_sc_hd__nor2_1 _1176_ (.A(_0272_),
    .B(_0448_),
    .Y(_0493_));
 sky130_fd_sc_hd__a221o_2 _1177_ (.A1(_0286_),
    .A2(_0491_),
    .B1(_0492_),
    .B2(_0493_),
    .C1(_0270_),
    .X(_0494_));
 sky130_fd_sc_hd__a21oi_1 _1178_ (.A1(_0489_),
    .A2(_0494_),
    .B1(_0327_),
    .Y(_0495_));
 sky130_fd_sc_hd__xnor2_1 _1179_ (.A(_0485_),
    .B(_0495_),
    .Y(_0900_));
 sky130_fd_sc_hd__nand2_1 _1180_ (.A(_0377_),
    .B(_0432_),
    .Y(_0496_));
 sky130_fd_sc_hd__and3_1 _1181_ (.A(_0447_),
    .B(_0457_),
    .C(_0483_),
    .X(_0497_));
 sky130_fd_sc_hd__a31oi_1 _1182_ (.A1(_0485_),
    .A2(_0494_),
    .A3(_0497_),
    .B1(_0347_),
    .Y(_0498_));
 sky130_fd_sc_hd__xnor2_1 _1183_ (.A(_0496_),
    .B(_0498_),
    .Y(_0903_));
 sky130_fd_sc_hd__inv_1 _1184_ (.A(\state[0] ),
    .Y(_0909_));
 sky130_fd_sc_hd__nor2_1 _1185_ (.A(_0302_),
    .B(_0751_),
    .Y(_0499_));
 sky130_fd_sc_hd__a21oi_1 _1186_ (.A1(_0302_),
    .A2(_0748_),
    .B1(_0499_),
    .Y(_0734_));
 sky130_fd_sc_hd__a21boi_1 _1187_ (.A1(_0285_),
    .A2(_0773_),
    .B1_N(_0420_),
    .Y(_0500_));
 sky130_fd_sc_hd__nor2_1 _1188_ (.A(_0302_),
    .B(_0750_),
    .Y(_0501_));
 sky130_fd_sc_hd__xnor2_1 _1189_ (.A(_0500_),
    .B(_0501_),
    .Y(_0754_));
 sky130_fd_sc_hd__o21ai_0 _1190_ (.A1(_0771_),
    .A2(_0767_),
    .B1(_0288_),
    .Y(_0502_));
 sky130_fd_sc_hd__and2_0 _1191_ (.A(_0749_),
    .B(_0748_),
    .X(_0503_));
 sky130_fd_sc_hd__a21oi_1 _1192_ (.A1(_0500_),
    .A2(_0503_),
    .B1(_0327_),
    .Y(_0504_));
 sky130_fd_sc_hd__xnor2_1 _1193_ (.A(_0502_),
    .B(_0504_),
    .Y(_0757_));
 sky130_fd_sc_hd__a21oi_1 _1194_ (.A1(_0750_),
    .A2(_0289_),
    .B1(_0327_),
    .Y(_0505_));
 sky130_fd_sc_hd__xnor2_1 _1195_ (.A(_0299_),
    .B(_0505_),
    .Y(_0760_));
 sky130_fd_sc_hd__a31oi_1 _1196_ (.A1(_0289_),
    .A2(_0299_),
    .A3(_0503_),
    .B1(_0347_),
    .Y(_0506_));
 sky130_fd_sc_hd__xor2_1 _1197_ (.A(_0296_),
    .B(_0506_),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_1 _1198_ (.A(_0313_),
    .B(_0279_),
    .Y(_0507_));
 sky130_fd_sc_hd__a21oi_1 _1199_ (.A1(_0293_),
    .A2(_0507_),
    .B1(_0270_),
    .Y(_0508_));
 sky130_fd_sc_hd__nor2_1 _1200_ (.A(_0327_),
    .B(_0300_),
    .Y(_0509_));
 sky130_fd_sc_hd__xor2_1 _1201_ (.A(_0508_),
    .B(_0509_),
    .X(_0784_));
 sky130_fd_sc_hd__nor2_1 _1202_ (.A(_0296_),
    .B(_0508_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand4_1 _1203_ (.A(_0289_),
    .B(_0299_),
    .C(_0503_),
    .D(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__and2_0 _1204_ (.A(_0364_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__nand2_1 _1205_ (.A(_0417_),
    .B(_0763_),
    .Y(_0513_));
 sky130_fd_sc_hd__a21oi_1 _1206_ (.A1(_0293_),
    .A2(_0513_),
    .B1(_0281_),
    .Y(_0514_));
 sky130_fd_sc_hd__xor2_1 _1207_ (.A(_0512_),
    .B(_0514_),
    .X(_0787_));
 sky130_fd_sc_hd__o21ai_0 _1208_ (.A1(_0313_),
    .A2(_0766_),
    .B1(_0285_),
    .Y(_0515_));
 sky130_fd_sc_hd__a21oi_2 _1209_ (.A1(_0300_),
    .A2(_0515_),
    .B1(_0349_),
    .Y(_0516_));
 sky130_fd_sc_hd__mux2i_1 _1210_ (.A0(_0268_),
    .A1(_0773_),
    .S(_0417_),
    .Y(_0517_));
 sky130_fd_sc_hd__nor2_1 _1211_ (.A(_0281_),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__xor2_1 _1212_ (.A(_0516_),
    .B(_0518_),
    .X(_0790_));
 sky130_fd_sc_hd__mux2i_1 _1213_ (.A0(_0773_),
    .A1(_0765_),
    .S(_0417_),
    .Y(_0519_));
 sky130_fd_sc_hd__nor2_1 _1214_ (.A(_0281_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__xor2_1 _1215_ (.A(_0512_),
    .B(_0520_),
    .X(_0793_));
 sky130_fd_sc_hd__nand2_1 _1216_ (.A(_0777_),
    .B(_0401_),
    .Y(_0521_));
 sky130_fd_sc_hd__xnor2_1 _1217_ (.A(_0516_),
    .B(_0521_),
    .Y(_0796_));
 sky130_fd_sc_hd__inv_1 _1218_ (.A(_0765_),
    .Y(_0522_));
 sky130_fd_sc_hd__nor3_1 _1219_ (.A(_0313_),
    .B(_0268_),
    .C(_0777_),
    .Y(_0523_));
 sky130_fd_sc_hd__a21oi_1 _1220_ (.A1(_0313_),
    .A2(_0522_),
    .B1(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__nor2_1 _1221_ (.A(_0773_),
    .B(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__nor2_1 _1222_ (.A(_0281_),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__nor2_1 _1223_ (.A(_0511_),
    .B(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__nor2_1 _1224_ (.A(_0349_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand2_1 _1225_ (.A(_0769_),
    .B(_0401_),
    .Y(_0529_));
 sky130_fd_sc_hd__xnor2_1 _1226_ (.A(_0528_),
    .B(_0529_),
    .Y(_0799_));
 sky130_fd_sc_hd__nand2_1 _1227_ (.A(_0773_),
    .B(_0401_),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_1 _1228_ (.A(_0769_),
    .Y(_0531_));
 sky130_fd_sc_hd__a21oi_1 _1229_ (.A1(_0364_),
    .A2(_0531_),
    .B1(_0458_),
    .Y(_0532_));
 sky130_fd_sc_hd__nor2_1 _1230_ (.A(_0526_),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__a21oi_1 _1231_ (.A1(_0347_),
    .A2(_0530_),
    .B1(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__o22a_1 _1232_ (.A1(_0302_),
    .A2(_0530_),
    .B1(_0534_),
    .B2(_0516_),
    .X(_0802_));
 sky130_fd_sc_hd__a21oi_1 _1233_ (.A1(_0531_),
    .A2(_0527_),
    .B1(_0302_),
    .Y(_0535_));
 sky130_fd_sc_hd__o21ai_0 _1234_ (.A1(_0349_),
    .A2(_0531_),
    .B1(_0522_),
    .Y(_0536_));
 sky130_fd_sc_hd__a21oi_1 _1235_ (.A1(_0401_),
    .A2(_0536_),
    .B1(_0528_),
    .Y(_0537_));
 sky130_fd_sc_hd__a31oi_1 _1236_ (.A1(_0765_),
    .A2(_0401_),
    .A3(_0535_),
    .B1(_0537_),
    .Y(_0805_));
 sky130_fd_sc_hd__nor2_1 _1237_ (.A(_0364_),
    .B(_0815_),
    .Y(_0538_));
 sky130_fd_sc_hd__a21oi_2 _1238_ (.A1(_0364_),
    .A2(_0818_),
    .B1(_0538_),
    .Y(_0738_));
 sky130_fd_sc_hd__inv_1 _1239_ (.A(_0445_),
    .Y(_0864_));
 sky130_fd_sc_hd__nor2_1 _1240_ (.A(_0327_),
    .B(_0865_),
    .Y(_0539_));
 sky130_fd_sc_hd__xor2_1 _1241_ (.A(_0487_),
    .B(_0539_),
    .X(_0870_));
 sky130_fd_sc_hd__nand3_1 _1242_ (.A(_0476_),
    .B(_0477_),
    .C(_0478_),
    .Y(_0540_));
 sky130_fd_sc_hd__inv_1 _1243_ (.A(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__nor2_1 _1244_ (.A(_0302_),
    .B(_0457_),
    .Y(_0542_));
 sky130_fd_sc_hd__xnor2_1 _1245_ (.A(_0541_),
    .B(_0542_),
    .Y(_0873_));
 sky130_fd_sc_hd__a21oi_1 _1246_ (.A1(_0541_),
    .A2(_0488_),
    .B1(_0327_),
    .Y(_0543_));
 sky130_fd_sc_hd__xnor2_1 _1247_ (.A(_0473_),
    .B(_0543_),
    .Y(_0876_));
 sky130_fd_sc_hd__a31oi_1 _1248_ (.A1(_0457_),
    .A2(_0473_),
    .A3(_0541_),
    .B1(_0347_),
    .Y(_0544_));
 sky130_fd_sc_hd__xor2_1 _1249_ (.A(_0481_),
    .B(_0544_),
    .X(_0879_));
 sky130_fd_sc_hd__nor2_1 _1250_ (.A(_0479_),
    .B(_0481_),
    .Y(_0545_));
 sky130_fd_sc_hd__a21oi_1 _1251_ (.A1(_0545_),
    .A2(_0488_),
    .B1(_0347_),
    .Y(_0546_));
 sky130_fd_sc_hd__xor2_1 _1252_ (.A(_0472_),
    .B(_0546_),
    .X(_0882_));
 sky130_fd_sc_hd__nor3_1 _1253_ (.A(_0472_),
    .B(_0479_),
    .C(_0481_),
    .Y(_0547_));
 sky130_fd_sc_hd__a21oi_1 _1254_ (.A1(_0457_),
    .A2(_0547_),
    .B1(_0347_),
    .Y(_0548_));
 sky130_fd_sc_hd__xor2_1 _1255_ (.A(_0470_),
    .B(_0548_),
    .X(_0885_));
 sky130_fd_sc_hd__a21oi_1 _1256_ (.A1(_0482_),
    .A2(_0488_),
    .B1(_0347_),
    .Y(_0549_));
 sky130_fd_sc_hd__xor2_1 _1257_ (.A(_0461_),
    .B(_0549_),
    .X(_0888_));
 sky130_fd_sc_hd__nand2_1 _1258_ (.A(_0313_),
    .B(_0452_),
    .Y(_0550_));
 sky130_fd_sc_hd__o21ai_0 _1259_ (.A1(_0313_),
    .A2(_0471_),
    .B1(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _1260_ (.A(_0285_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__nor2_1 _1261_ (.A(_0327_),
    .B(_0489_),
    .Y(_0553_));
 sky130_fd_sc_hd__xnor2_1 _1262_ (.A(_0552_),
    .B(_0553_),
    .Y(_0894_));
 sky130_fd_sc_hd__a21oi_1 _1263_ (.A1(_0497_),
    .A2(_0552_),
    .B1(_0347_),
    .Y(_0554_));
 sky130_fd_sc_hd__and2_0 _1264_ (.A(_0292_),
    .B(_0468_),
    .X(_0555_));
 sky130_fd_sc_hd__a31oi_1 _1265_ (.A1(_0417_),
    .A2(_0425_),
    .A3(_0393_),
    .B1(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nor2_1 _1266_ (.A(_0281_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__xor2_1 _1267_ (.A(_0554_),
    .B(_0557_),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_1 _1268_ (.A(_0377_),
    .B(_0452_),
    .Y(_0558_));
 sky130_fd_sc_hd__a41oi_1 _1269_ (.A1(_0485_),
    .A2(_0489_),
    .A3(_0494_),
    .A4(_0496_),
    .B1(_0349_),
    .Y(_0559_));
 sky130_fd_sc_hd__xnor2_1 _1270_ (.A(_0558_),
    .B(_0559_),
    .Y(_0906_));
 sky130_fd_sc_hd__inv_1 _1271_ (.A(\state[1] ),
    .Y(_0910_));
 sky130_fd_sc_hd__clkbuf_4 _1272_ (.A(\next_state[1] ),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_4 _1273_ (.A(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__buf_4 _1274_ (.A(_0914_),
    .X(_0562_));
 sky130_fd_sc_hd__nand2_2 _1275_ (.A(_0562_),
    .B(\next_state[1] ),
    .Y(_0563_));
 sky130_fd_sc_hd__mux2i_1 _1276_ (.A0(_0561_),
    .A1(_0563_),
    .S(_0763_),
    .Y(_0001_));
 sky130_fd_sc_hd__buf_4 _1277_ (.A(_0562_),
    .X(_0564_));
 sky130_fd_sc_hd__clkbuf_4 _1278_ (.A(_0560_),
    .X(_0565_));
 sky130_fd_sc_hd__nand3_1 _1279_ (.A(_0564_),
    .B(_0766_),
    .C(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__o21ai_0 _1280_ (.A1(_0764_),
    .A2(_0561_),
    .B1(_0566_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand2_1 _1281_ (.A(_0292_),
    .B(_0779_),
    .Y(_0567_));
 sky130_fd_sc_hd__inv_2 _1282_ (.A(_0914_),
    .Y(_0568_));
 sky130_fd_sc_hd__buf_4 _1283_ (.A(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_4 _1284_ (.A(\next_state[1] ),
    .X(_0570_));
 sky130_fd_sc_hd__o21ai_0 _1285_ (.A1(_0779_),
    .A2(_0569_),
    .B1(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__nand2_1 _1286_ (.A(_0417_),
    .B(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__o21ai_0 _1287_ (.A1(_0563_),
    .A2(_0567_),
    .B1(_0572_),
    .Y(_0003_));
 sky130_fd_sc_hd__nand3_1 _1288_ (.A(_0417_),
    .B(_0279_),
    .C(_0268_),
    .Y(_0573_));
 sky130_fd_sc_hd__buf_4 _1289_ (.A(_0560_),
    .X(_0574_));
 sky130_fd_sc_hd__nand2_1 _1290_ (.A(_0564_),
    .B(_0573_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _1291_ (.A(_0574_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_1 _1292_ (.A(_0281_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__o31ai_1 _1293_ (.A1(_0281_),
    .A2(_0563_),
    .A3(_0573_),
    .B1(_0577_),
    .Y(_0004_));
 sky130_fd_sc_hd__buf_4 _1294_ (.A(_0562_),
    .X(_0578_));
 sky130_fd_sc_hd__nor2b_1 _1295_ (.A(net2),
    .B_N(_0911_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand3_1 _1296_ (.A(_0292_),
    .B(_0281_),
    .C(_0779_),
    .Y(_0580_));
 sky130_fd_sc_hd__a21oi_1 _1297_ (.A1(_0578_),
    .A2(_0580_),
    .B1(_0579_),
    .Y(_0581_));
 sky130_fd_sc_hd__o32a_1 _1298_ (.A1(_0578_),
    .A2(_0912_),
    .A3(_0579_),
    .B1(_0581_),
    .B2(\state[0] ),
    .X(_0005_));
 sky130_fd_sc_hd__buf_4 _1299_ (.A(_0560_),
    .X(_0582_));
 sky130_fd_sc_hd__nand2_1 _1300_ (.A(_0582_),
    .B(_0581_),
    .Y(_0583_));
 sky130_fd_sc_hd__o21ai_0 _1301_ (.A1(_0910_),
    .A2(_0581_),
    .B1(_0583_),
    .Y(_0006_));
 sky130_fd_sc_hd__buf_2 _1302_ (.A(_0570_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2i_1 _1303_ (.A0(net3),
    .A1(_0862_),
    .S(_0564_),
    .Y(_0585_));
 sky130_fd_sc_hd__nor2_1 _1304_ (.A(\x[0] ),
    .B(_0582_),
    .Y(_0586_));
 sky130_fd_sc_hd__a21oi_1 _1305_ (.A1(_0584_),
    .A2(_0585_),
    .B1(_0586_),
    .Y(_0007_));
 sky130_fd_sc_hd__nor2b_1 _1306_ (.A(_0744_),
    .B_N(_0872_),
    .Y(_0587_));
 sky130_fd_sc_hd__o21a_1 _1307_ (.A1(_0871_),
    .A2(_0587_),
    .B1(_0875_),
    .X(_0588_));
 sky130_fd_sc_hd__o21ai_1 _1308_ (.A1(_0874_),
    .A2(_0588_),
    .B1(_0878_),
    .Y(_0589_));
 sky130_fd_sc_hd__nor3_1 _1309_ (.A(_0877_),
    .B(_0880_),
    .C(_0883_),
    .Y(_0590_));
 sky130_fd_sc_hd__o21a_1 _1310_ (.A1(_0881_),
    .A2(_0880_),
    .B1(_0884_),
    .X(_0591_));
 sky130_fd_sc_hd__o21ai_0 _1311_ (.A1(_0883_),
    .A2(_0591_),
    .B1(_0887_),
    .Y(_0592_));
 sky130_fd_sc_hd__a21oi_1 _1312_ (.A1(_0589_),
    .A2(_0590_),
    .B1(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__o21a_1 _1313_ (.A1(_0890_),
    .A2(_0889_),
    .B1(_0893_),
    .X(_0594_));
 sky130_fd_sc_hd__o31ai_2 _1314_ (.A1(_0886_),
    .A2(_0889_),
    .A3(_0593_),
    .B1(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2b_1 _1315_ (.A_N(_0892_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__xor2_1 _1316_ (.A(_0896_),
    .B(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__buf_6 _1317_ (.A(_0562_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2i_1 _1318_ (.A0(net4),
    .A1(_0597_),
    .S(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__nor2_1 _1319_ (.A(\x[10] ),
    .B(_0582_),
    .Y(_0600_));
 sky130_fd_sc_hd__a21oi_1 _1320_ (.A1(_0584_),
    .A2(_0599_),
    .B1(_0600_),
    .Y(_0008_));
 sky130_fd_sc_hd__nand2b_1 _1321_ (.A_N(_0878_),
    .B(_0590_),
    .Y(_0601_));
 sky130_fd_sc_hd__a211oi_2 _1322_ (.A1(_0861_),
    .A2(_0869_),
    .B1(_0868_),
    .C1(_0871_),
    .Y(_0602_));
 sky130_fd_sc_hd__o21ai_0 _1323_ (.A1(_0872_),
    .A2(_0871_),
    .B1(_0875_),
    .Y(_0603_));
 sky130_fd_sc_hd__nor4_1 _1324_ (.A(_0874_),
    .B(_0877_),
    .C(_0880_),
    .D(_0883_),
    .Y(_0604_));
 sky130_fd_sc_hd__o21ai_0 _1325_ (.A1(_0602_),
    .A2(_0603_),
    .B1(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__nand3b_1 _1326_ (.A_N(_0592_),
    .B(_0601_),
    .C(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__nor3_1 _1327_ (.A(_0886_),
    .B(_0889_),
    .C(_0892_),
    .Y(_0607_));
 sky130_fd_sc_hd__nor2_1 _1328_ (.A(_0892_),
    .B(_0594_),
    .Y(_0608_));
 sky130_fd_sc_hd__a21oi_2 _1329_ (.A1(_0606_),
    .A2(_0607_),
    .B1(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__a21oi_1 _1330_ (.A1(_0896_),
    .A2(_0609_),
    .B1(_0895_),
    .Y(_0610_));
 sky130_fd_sc_hd__xnor2_1 _1331_ (.A(_0899_),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__mux2i_1 _1332_ (.A0(net5),
    .A1(_0611_),
    .S(_0598_),
    .Y(_0612_));
 sky130_fd_sc_hd__nor2_1 _1333_ (.A(\x[11] ),
    .B(_0582_),
    .Y(_0613_));
 sky130_fd_sc_hd__a21oi_1 _1334_ (.A1(_0584_),
    .A2(_0612_),
    .B1(_0613_),
    .Y(_0009_));
 sky130_fd_sc_hd__nor3_1 _1335_ (.A(_0892_),
    .B(_0895_),
    .C(_0898_),
    .Y(_0614_));
 sky130_fd_sc_hd__or2_0 _1336_ (.A(_0896_),
    .B(_0895_),
    .X(_0615_));
 sky130_fd_sc_hd__a21oi_1 _1337_ (.A1(_0899_),
    .A2(_0615_),
    .B1(_0898_),
    .Y(_0616_));
 sky130_fd_sc_hd__a21oi_1 _1338_ (.A1(_0595_),
    .A2(_0614_),
    .B1(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__xor2_1 _1339_ (.A(_0902_),
    .B(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2i_1 _1340_ (.A0(net6),
    .A1(_0618_),
    .S(_0598_),
    .Y(_0619_));
 sky130_fd_sc_hd__nor2_1 _1341_ (.A(\x[12] ),
    .B(_0582_),
    .Y(_0620_));
 sky130_fd_sc_hd__a21oi_1 _1342_ (.A1(_0584_),
    .A2(_0619_),
    .B1(_0620_),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_1 _1343_ (.A(_0902_),
    .B(_0898_),
    .Y(_0621_));
 sky130_fd_sc_hd__nand3_1 _1344_ (.A(_0899_),
    .B(_0902_),
    .C(_0895_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_1 _1345_ (.A(_0621_),
    .B(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__a41o_1 _1346_ (.A1(_0896_),
    .A2(_0899_),
    .A3(_0902_),
    .A4(_0609_),
    .B1(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__nor2_1 _1347_ (.A(_0901_),
    .B(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__xnor2_1 _1348_ (.A(_0905_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__mux2i_1 _1349_ (.A0(net7),
    .A1(_0626_),
    .S(_0598_),
    .Y(_0627_));
 sky130_fd_sc_hd__nor2_1 _1350_ (.A(\x[13] ),
    .B(_0582_),
    .Y(_0628_));
 sky130_fd_sc_hd__a21oi_1 _1351_ (.A1(_0584_),
    .A2(_0627_),
    .B1(_0628_),
    .Y(_0011_));
 sky130_fd_sc_hd__nand2b_1 _1352_ (.A_N(_0570_),
    .B(\x[14] ),
    .Y(_0629_));
 sky130_fd_sc_hd__nand3b_1 _1353_ (.A_N(_0908_),
    .B(_0560_),
    .C(_0562_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand3_1 _1354_ (.A(_0578_),
    .B(_0908_),
    .C(\next_state[1] ),
    .Y(_0631_));
 sky130_fd_sc_hd__a21o_1 _1355_ (.A1(_0905_),
    .A2(_0901_),
    .B1(_0904_),
    .X(_0632_));
 sky130_fd_sc_hd__a31oi_1 _1356_ (.A1(_0902_),
    .A2(_0905_),
    .A3(_0617_),
    .B1(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__mux2_1 _1357_ (.A0(_0630_),
    .A1(_0631_),
    .S(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__nand3_1 _1358_ (.A(_0569_),
    .B(net8),
    .C(_0565_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand3_1 _1359_ (.A(_0629_),
    .B(_0634_),
    .C(_0635_),
    .Y(_0012_));
 sky130_fd_sc_hd__nand4_1 _1360_ (.A(_0485_),
    .B(_0494_),
    .C(_0496_),
    .D(_0558_),
    .Y(_0636_));
 sky130_fd_sc_hd__nor3b_1 _1361_ (.A(_0636_),
    .B(_0461_),
    .C_N(_0447_),
    .Y(_0637_));
 sky130_fd_sc_hd__a31oi_1 _1362_ (.A1(_0457_),
    .A2(_0482_),
    .A3(_0637_),
    .B1(_0301_),
    .Y(_0638_));
 sky130_fd_sc_hd__inv_1 _1363_ (.A(\x[15] ),
    .Y(_0639_));
 sky130_fd_sc_hd__nand3_1 _1364_ (.A(_0425_),
    .B(_0377_),
    .C(_0393_),
    .Y(_0640_));
 sky130_fd_sc_hd__xnor2_1 _1365_ (.A(_0639_),
    .B(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__xnor2_1 _1366_ (.A(_0638_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nor4_1 _1367_ (.A(_0907_),
    .B(_0901_),
    .C(_0904_),
    .D(_0624_),
    .Y(_0643_));
 sky130_fd_sc_hd__nor3_1 _1368_ (.A(_0907_),
    .B(_0905_),
    .C(_0904_),
    .Y(_0644_));
 sky130_fd_sc_hd__nor2_1 _1369_ (.A(_0907_),
    .B(_0908_),
    .Y(_0645_));
 sky130_fd_sc_hd__nor3_1 _1370_ (.A(_0645_),
    .B(_0644_),
    .C(_0643_),
    .Y(_0646_));
 sky130_fd_sc_hd__nor2_1 _1371_ (.A(_0563_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand3_1 _1372_ (.A(_0568_),
    .B(net9),
    .C(_0560_),
    .Y(_0648_));
 sky130_fd_sc_hd__o21ai_0 _1373_ (.A1(_0639_),
    .A2(_0560_),
    .B1(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__nor3b_1 _1374_ (.A(_0563_),
    .B(_0642_),
    .C_N(_0646_),
    .Y(_0650_));
 sky130_fd_sc_hd__a211o_1 _1375_ (.A1(_0642_),
    .A2(_0647_),
    .B1(_0649_),
    .C1(_0650_),
    .X(_0013_));
 sky130_fd_sc_hd__nand2_1 _1376_ (.A(_0564_),
    .B(_0745_),
    .Y(_0651_));
 sky130_fd_sc_hd__o211ai_1 _1377_ (.A1(_0564_),
    .A2(net10),
    .B1(_0574_),
    .C1(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__o21ai_0 _1378_ (.A1(_0741_),
    .A2(_0582_),
    .B1(_0652_),
    .Y(_0014_));
 sky130_fd_sc_hd__nor2b_1 _1379_ (.A(_0872_),
    .B_N(_0744_),
    .Y(_0653_));
 sky130_fd_sc_hd__nor3_1 _1380_ (.A(_0569_),
    .B(_0587_),
    .C(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__a21oi_1 _1381_ (.A1(_0569_),
    .A2(net11),
    .B1(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__nor2_1 _1382_ (.A(\x[2] ),
    .B(_0582_),
    .Y(_0656_));
 sky130_fd_sc_hd__a21oi_1 _1383_ (.A1(_0584_),
    .A2(_0655_),
    .B1(_0656_),
    .Y(_0015_));
 sky130_fd_sc_hd__nor2_1 _1384_ (.A(_0602_),
    .B(_0603_),
    .Y(_0657_));
 sky130_fd_sc_hd__a21o_1 _1385_ (.A1(_0861_),
    .A2(_0869_),
    .B1(_0868_),
    .X(_0658_));
 sky130_fd_sc_hd__a211oi_1 _1386_ (.A1(_0872_),
    .A2(_0658_),
    .B1(_0871_),
    .C1(_0875_),
    .Y(_0659_));
 sky130_fd_sc_hd__nor3_1 _1387_ (.A(_0568_),
    .B(_0657_),
    .C(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__a21oi_1 _1388_ (.A1(_0569_),
    .A2(net12),
    .B1(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__buf_4 _1389_ (.A(_0560_),
    .X(_0662_));
 sky130_fd_sc_hd__nor2_1 _1390_ (.A(\x[3] ),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__a21oi_1 _1391_ (.A1(_0584_),
    .A2(_0661_),
    .B1(_0663_),
    .Y(_0016_));
 sky130_fd_sc_hd__or3_1 _1392_ (.A(_0878_),
    .B(_0874_),
    .C(_0588_),
    .X(_0664_));
 sky130_fd_sc_hd__nor2b_1 _1393_ (.A(_0562_),
    .B_N(net13),
    .Y(_0665_));
 sky130_fd_sc_hd__a31oi_1 _1394_ (.A1(_0564_),
    .A2(_0589_),
    .A3(_0664_),
    .B1(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__nor2_1 _1395_ (.A(\x[4] ),
    .B(_0662_),
    .Y(_0667_));
 sky130_fd_sc_hd__a21oi_1 _1396_ (.A1(_0584_),
    .A2(_0666_),
    .B1(_0667_),
    .Y(_0017_));
 sky130_fd_sc_hd__o21a_1 _1397_ (.A1(_0874_),
    .A2(_0657_),
    .B1(_0878_),
    .X(_0668_));
 sky130_fd_sc_hd__nor2_1 _1398_ (.A(_0877_),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__xnor2_1 _1399_ (.A(_0881_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__mux2i_1 _1400_ (.A0(net14),
    .A1(_0670_),
    .S(_0598_),
    .Y(_0671_));
 sky130_fd_sc_hd__nor2_1 _1401_ (.A(\x[5] ),
    .B(_0662_),
    .Y(_0672_));
 sky130_fd_sc_hd__a21oi_1 _1402_ (.A1(_0584_),
    .A2(_0671_),
    .B1(_0672_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2b_1 _1403_ (.A_N(_0877_),
    .B(_0589_),
    .Y(_0673_));
 sky130_fd_sc_hd__a21oi_1 _1404_ (.A1(_0881_),
    .A2(_0673_),
    .B1(_0880_),
    .Y(_0674_));
 sky130_fd_sc_hd__xnor2_1 _1405_ (.A(_0884_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__mux2i_1 _1406_ (.A0(net15),
    .A1(_0675_),
    .S(_0598_),
    .Y(_0676_));
 sky130_fd_sc_hd__nor2_1 _1407_ (.A(\x[6] ),
    .B(_0662_),
    .Y(_0677_));
 sky130_fd_sc_hd__a21oi_1 _1408_ (.A1(_0584_),
    .A2(_0676_),
    .B1(_0677_),
    .Y(_0019_));
 sky130_fd_sc_hd__buf_4 _1409_ (.A(_0570_),
    .X(_0678_));
 sky130_fd_sc_hd__o21ai_0 _1410_ (.A1(_0877_),
    .A2(_0668_),
    .B1(_0881_),
    .Y(_0679_));
 sky130_fd_sc_hd__nand2b_1 _1411_ (.A_N(_0880_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__a211o_1 _1412_ (.A1(_0884_),
    .A2(_0680_),
    .B1(_0883_),
    .C1(_0887_),
    .X(_0681_));
 sky130_fd_sc_hd__nor2b_1 _1413_ (.A(_0562_),
    .B_N(net16),
    .Y(_0682_));
 sky130_fd_sc_hd__a31oi_1 _1414_ (.A1(_0564_),
    .A2(_0606_),
    .A3(_0681_),
    .B1(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__nor2_1 _1415_ (.A(\x[7] ),
    .B(_0662_),
    .Y(_0684_));
 sky130_fd_sc_hd__a21oi_1 _1416_ (.A1(_0678_),
    .A2(_0683_),
    .B1(_0684_),
    .Y(_0020_));
 sky130_fd_sc_hd__nor2_1 _1417_ (.A(_0886_),
    .B(_0593_),
    .Y(_0685_));
 sky130_fd_sc_hd__xnor2_1 _1418_ (.A(_0890_),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__mux2i_1 _1419_ (.A0(net17),
    .A1(_0686_),
    .S(_0598_),
    .Y(_0687_));
 sky130_fd_sc_hd__nor2_1 _1420_ (.A(\x[8] ),
    .B(_0662_),
    .Y(_0688_));
 sky130_fd_sc_hd__a21oi_1 _1421_ (.A1(_0678_),
    .A2(_0687_),
    .B1(_0688_),
    .Y(_0021_));
 sky130_fd_sc_hd__nand2b_1 _1422_ (.A_N(_0886_),
    .B(_0606_),
    .Y(_0689_));
 sky130_fd_sc_hd__a21oi_1 _1423_ (.A1(_0890_),
    .A2(_0689_),
    .B1(_0889_),
    .Y(_0690_));
 sky130_fd_sc_hd__xnor2_1 _1424_ (.A(_0893_),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__mux2i_1 _1425_ (.A0(net18),
    .A1(_0691_),
    .S(_0598_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor2_1 _1426_ (.A(\x[9] ),
    .B(_0662_),
    .Y(_0693_));
 sky130_fd_sc_hd__a21oi_1 _1427_ (.A1(_0678_),
    .A2(_0692_),
    .B1(_0693_),
    .Y(_0022_));
 sky130_fd_sc_hd__clkbuf_4 _1428_ (.A(_0916_),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_4 _1429_ (.A(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _1430_ (.A0(net52),
    .A1(\x[0] ),
    .S(_0695_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _1431_ (.A0(net53),
    .A1(\x[10] ),
    .S(_0695_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(net54),
    .A1(\x[11] ),
    .S(_0695_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1433_ (.A0(net55),
    .A1(\x[12] ),
    .S(_0695_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _1434_ (.A0(net56),
    .A1(\x[13] ),
    .S(_0695_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1435_ (.A0(net57),
    .A1(\x[14] ),
    .S(_0695_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1436_ (.A0(net58),
    .A1(\x[15] ),
    .S(_0695_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1437_ (.A0(net59),
    .A1(\x[1] ),
    .S(_0695_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(net60),
    .A1(\x[2] ),
    .S(_0695_),
    .X(_0031_));
 sky130_fd_sc_hd__buf_4 _1439_ (.A(_0916_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(net61),
    .A1(\x[3] ),
    .S(_0696_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1441_ (.A0(net62),
    .A1(\x[4] ),
    .S(_0696_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _1442_ (.A0(net63),
    .A1(\x[5] ),
    .S(_0696_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _1443_ (.A0(net64),
    .A1(\x[6] ),
    .S(_0696_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(net65),
    .A1(\x[7] ),
    .S(_0696_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _1445_ (.A0(net66),
    .A1(\x[8] ),
    .S(_0696_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _1446_ (.A0(net67),
    .A1(\x[9] ),
    .S(_0696_),
    .X(_0038_));
 sky130_fd_sc_hd__nand2_1 _1447_ (.A(_0564_),
    .B(_0814_),
    .Y(_0697_));
 sky130_fd_sc_hd__o211ai_1 _1448_ (.A1(_0564_),
    .A2(net19),
    .B1(_0574_),
    .C1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__o21ai_0 _1449_ (.A1(_0811_),
    .A2(_0582_),
    .B1(_0698_),
    .Y(_0039_));
 sky130_fd_sc_hd__o21a_1 _1450_ (.A1(_0832_),
    .A2(_0831_),
    .B1(_0835_),
    .X(_0699_));
 sky130_fd_sc_hd__o21ai_0 _1451_ (.A1(_0834_),
    .A2(_0699_),
    .B1(_0838_),
    .Y(_0700_));
 sky130_fd_sc_hd__a21o_1 _1452_ (.A1(_0739_),
    .A2(_0823_),
    .B1(_0822_),
    .X(_0701_));
 sky130_fd_sc_hd__a21o_1 _1453_ (.A1(_0826_),
    .A2(_0701_),
    .B1(_0825_),
    .X(_0702_));
 sky130_fd_sc_hd__or3_1 _1454_ (.A(_0828_),
    .B(_0831_),
    .C(_0834_),
    .X(_0703_));
 sky130_fd_sc_hd__a21oi_1 _1455_ (.A1(_0829_),
    .A2(_0702_),
    .B1(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__nor2_1 _1456_ (.A(_0837_),
    .B(_0840_),
    .Y(_0705_));
 sky130_fd_sc_hd__o21ai_1 _1457_ (.A1(_0700_),
    .A2(_0704_),
    .B1(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__o21a_1 _1458_ (.A1(_0841_),
    .A2(_0840_),
    .B1(_0844_),
    .X(_0707_));
 sky130_fd_sc_hd__a21oi_1 _1459_ (.A1(_0706_),
    .A2(_0707_),
    .B1(_0843_),
    .Y(_0708_));
 sky130_fd_sc_hd__xnor2_1 _1460_ (.A(_0847_),
    .B(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__mux2i_1 _1461_ (.A0(net20),
    .A1(_0709_),
    .S(_0598_),
    .Y(_0710_));
 sky130_fd_sc_hd__nor2_1 _1462_ (.A(\y[10] ),
    .B(_0662_),
    .Y(_0711_));
 sky130_fd_sc_hd__a21oi_1 _1463_ (.A1(_0678_),
    .A2(_0710_),
    .B1(_0711_),
    .Y(_0040_));
 sky130_fd_sc_hd__nor2_1 _1464_ (.A(_0829_),
    .B(_0703_),
    .Y(_0712_));
 sky130_fd_sc_hd__nand2b_1 _1465_ (.A_N(_0813_),
    .B(_0820_),
    .Y(_0713_));
 sky130_fd_sc_hd__nor2_1 _1466_ (.A(_0819_),
    .B(_0822_),
    .Y(_0714_));
 sky130_fd_sc_hd__o21ai_0 _1467_ (.A1(_0823_),
    .A2(_0822_),
    .B1(_0826_),
    .Y(_0715_));
 sky130_fd_sc_hd__a21oi_2 _1468_ (.A1(_0713_),
    .A2(_0714_),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__o21a_1 _1469_ (.A1(_0834_),
    .A2(_0699_),
    .B1(_0838_),
    .X(_0717_));
 sky130_fd_sc_hd__o31ai_1 _1470_ (.A1(_0825_),
    .A2(_0703_),
    .A3(_0716_),
    .B1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__nor3_1 _1471_ (.A(_0837_),
    .B(_0840_),
    .C(_0843_),
    .Y(_0719_));
 sky130_fd_sc_hd__o21ai_1 _1472_ (.A1(_0712_),
    .A2(_0718_),
    .B1(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__or2_0 _1473_ (.A(_0843_),
    .B(_0707_),
    .X(_0721_));
 sky130_fd_sc_hd__a31oi_1 _1474_ (.A1(_0847_),
    .A2(_0720_),
    .A3(_0721_),
    .B1(_0846_),
    .Y(_0722_));
 sky130_fd_sc_hd__xnor2_1 _1475_ (.A(_0850_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__mux2i_1 _1476_ (.A0(net21),
    .A1(_0723_),
    .S(_0598_),
    .Y(_0724_));
 sky130_fd_sc_hd__nor2_1 _1477_ (.A(\y[11] ),
    .B(_0662_),
    .Y(_0725_));
 sky130_fd_sc_hd__a21oi_1 _1478_ (.A1(_0678_),
    .A2(_0724_),
    .B1(_0725_),
    .Y(_0041_));
 sky130_fd_sc_hd__a2111oi_2 _1479_ (.A1(_0706_),
    .A2(_0707_),
    .B1(_0843_),
    .C1(_0846_),
    .D1(_0849_),
    .Y(_0726_));
 sky130_fd_sc_hd__or2_0 _1480_ (.A(_0847_),
    .B(_0846_),
    .X(_0727_));
 sky130_fd_sc_hd__a21oi_1 _1481_ (.A1(_0850_),
    .A2(_0727_),
    .B1(_0849_),
    .Y(_0728_));
 sky130_fd_sc_hd__nor2_1 _1482_ (.A(_0726_),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__xor2_1 _1483_ (.A(_0853_),
    .B(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__clkbuf_8 _1484_ (.A(_0562_),
    .X(_0731_));
 sky130_fd_sc_hd__mux2i_1 _1485_ (.A0(net22),
    .A1(_0730_),
    .S(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__nor2_1 _1486_ (.A(\y[12] ),
    .B(_0662_),
    .Y(_0103_));
 sky130_fd_sc_hd__a21oi_1 _1487_ (.A1(_0678_),
    .A2(_0732_),
    .B1(_0103_),
    .Y(_0042_));
 sky130_fd_sc_hd__and3_1 _1488_ (.A(_0847_),
    .B(_0850_),
    .C(_0853_),
    .X(_0104_));
 sky130_fd_sc_hd__nand2_1 _1489_ (.A(_0853_),
    .B(_0849_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand3_1 _1490_ (.A(_0850_),
    .B(_0853_),
    .C(_0846_),
    .Y(_0106_));
 sky130_fd_sc_hd__nand2_1 _1491_ (.A(_0105_),
    .B(_0106_),
    .Y(_0107_));
 sky130_fd_sc_hd__a31oi_2 _1492_ (.A1(_0720_),
    .A2(_0721_),
    .A3(_0104_),
    .B1(_0107_),
    .Y(_0108_));
 sky130_fd_sc_hd__nor2b_1 _1493_ (.A(_0852_),
    .B_N(_0108_),
    .Y(_0109_));
 sky130_fd_sc_hd__xnor2_1 _1494_ (.A(_0856_),
    .B(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__mux2i_1 _1495_ (.A0(net23),
    .A1(_0110_),
    .S(_0731_),
    .Y(_0111_));
 sky130_fd_sc_hd__buf_4 _1496_ (.A(_0560_),
    .X(_0112_));
 sky130_fd_sc_hd__nor2_1 _1497_ (.A(\y[13] ),
    .B(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hd__a21oi_1 _1498_ (.A1(_0678_),
    .A2(_0111_),
    .B1(_0113_),
    .Y(_0043_));
 sky130_fd_sc_hd__nand2_1 _1499_ (.A(_0853_),
    .B(_0856_),
    .Y(_0114_));
 sky130_fd_sc_hd__a21oi_1 _1500_ (.A1(_0856_),
    .A2(_0852_),
    .B1(_0855_),
    .Y(_0115_));
 sky130_fd_sc_hd__o31ai_1 _1501_ (.A1(_0726_),
    .A2(_0728_),
    .A3(_0114_),
    .B1(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__xor2_1 _1502_ (.A(_0859_),
    .B(_0116_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2i_1 _1503_ (.A0(net24),
    .A1(_0117_),
    .S(_0731_),
    .Y(_0118_));
 sky130_fd_sc_hd__nor2_1 _1504_ (.A(\y[14] ),
    .B(_0112_),
    .Y(_0119_));
 sky130_fd_sc_hd__a21oi_1 _1505_ (.A1(_0678_),
    .A2(_0118_),
    .B1(_0119_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand3_1 _1506_ (.A(\x[15] ),
    .B(_0377_),
    .C(_0393_),
    .Y(_0120_));
 sky130_fd_sc_hd__xor2_1 _1507_ (.A(_0425_),
    .B(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__o31ai_2 _1508_ (.A1(net102),
    .A2(_0388_),
    .A3(_0405_),
    .B1(_0377_),
    .Y(_0122_));
 sky130_fd_sc_hd__a41oi_4 _1509_ (.A1(_0375_),
    .A2(_0395_),
    .A3(_0396_),
    .A4(_0122_),
    .B1(_0301_),
    .Y(_0123_));
 sky130_fd_sc_hd__xnor2_1 _1510_ (.A(_0121_),
    .B(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__nor3_1 _1511_ (.A(_0852_),
    .B(_0855_),
    .C(_0858_),
    .Y(_0125_));
 sky130_fd_sc_hd__or2_0 _1512_ (.A(_0856_),
    .B(_0855_),
    .X(_0126_));
 sky130_fd_sc_hd__a21oi_1 _1513_ (.A1(_0859_),
    .A2(_0126_),
    .B1(_0858_),
    .Y(_0127_));
 sky130_fd_sc_hd__a21oi_2 _1514_ (.A1(_0108_),
    .A2(_0125_),
    .B1(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__or3_1 _1515_ (.A(_0563_),
    .B(_0124_),
    .C(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__nand4_1 _1516_ (.A(_0564_),
    .B(_0574_),
    .C(_0124_),
    .D(_0128_),
    .Y(_0130_));
 sky130_fd_sc_hd__nor2b_1 _1517_ (.A(\next_state[1] ),
    .B_N(_0425_),
    .Y(_0131_));
 sky130_fd_sc_hd__a31oi_1 _1518_ (.A1(_0569_),
    .A2(net25),
    .A3(_0570_),
    .B1(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__nand3_1 _1519_ (.A(_0129_),
    .B(_0130_),
    .C(_0132_),
    .Y(_0045_));
 sky130_fd_sc_hd__mux2i_1 _1520_ (.A0(net26),
    .A1(_0740_),
    .S(_0731_),
    .Y(_0133_));
 sky130_fd_sc_hd__nor2_1 _1521_ (.A(\y[1] ),
    .B(_0112_),
    .Y(_0134_));
 sky130_fd_sc_hd__a21oi_1 _1522_ (.A1(_0678_),
    .A2(_0133_),
    .B1(_0134_),
    .Y(_0046_));
 sky130_fd_sc_hd__xnor2_1 _1523_ (.A(_0739_),
    .B(_0823_),
    .Y(_0135_));
 sky130_fd_sc_hd__nor2_1 _1524_ (.A(_0578_),
    .B(net27),
    .Y(_0136_));
 sky130_fd_sc_hd__a21oi_1 _1525_ (.A1(_0578_),
    .A2(_0135_),
    .B1(_0136_),
    .Y(_0137_));
 sky130_fd_sc_hd__mux2_1 _1526_ (.A0(\y[2] ),
    .A1(_0137_),
    .S(_0570_),
    .X(_0047_));
 sky130_fd_sc_hd__nand2b_1 _1527_ (.A_N(_0819_),
    .B(_0713_),
    .Y(_0138_));
 sky130_fd_sc_hd__a211oi_1 _1528_ (.A1(_0823_),
    .A2(_0138_),
    .B1(_0822_),
    .C1(_0826_),
    .Y(_0139_));
 sky130_fd_sc_hd__nand2_1 _1529_ (.A(_0569_),
    .B(net28),
    .Y(_0140_));
 sky130_fd_sc_hd__o311ai_0 _1530_ (.A1(_0568_),
    .A2(_0716_),
    .A3(_0139_),
    .B1(_0140_),
    .C1(_0570_),
    .Y(_0141_));
 sky130_fd_sc_hd__o21a_1 _1531_ (.A1(\y[3] ),
    .A2(_0582_),
    .B1(_0141_),
    .X(_0048_));
 sky130_fd_sc_hd__xor2_1 _1532_ (.A(_0829_),
    .B(_0702_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2i_1 _1533_ (.A0(net29),
    .A1(_0142_),
    .S(_0731_),
    .Y(_0143_));
 sky130_fd_sc_hd__nor2_1 _1534_ (.A(\y[4] ),
    .B(_0112_),
    .Y(_0144_));
 sky130_fd_sc_hd__a21oi_1 _1535_ (.A1(_0678_),
    .A2(_0143_),
    .B1(_0144_),
    .Y(_0049_));
 sky130_fd_sc_hd__clkbuf_4 _1536_ (.A(_0570_),
    .X(_0145_));
 sky130_fd_sc_hd__o21ai_0 _1537_ (.A1(_0825_),
    .A2(_0716_),
    .B1(_0829_),
    .Y(_0146_));
 sky130_fd_sc_hd__nand2b_1 _1538_ (.A_N(_0828_),
    .B(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__xor2_1 _1539_ (.A(_0832_),
    .B(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2i_1 _1540_ (.A0(net30),
    .A1(_0148_),
    .S(_0731_),
    .Y(_0149_));
 sky130_fd_sc_hd__nor2_1 _1541_ (.A(\y[5] ),
    .B(_0112_),
    .Y(_0150_));
 sky130_fd_sc_hd__a21oi_1 _1542_ (.A1(_0145_),
    .A2(_0149_),
    .B1(_0150_),
    .Y(_0050_));
 sky130_fd_sc_hd__a21o_1 _1543_ (.A1(_0829_),
    .A2(_0702_),
    .B1(_0828_),
    .X(_0151_));
 sky130_fd_sc_hd__a21oi_1 _1544_ (.A1(_0832_),
    .A2(_0151_),
    .B1(_0831_),
    .Y(_0152_));
 sky130_fd_sc_hd__xnor2_1 _1545_ (.A(_0835_),
    .B(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__mux2i_1 _1546_ (.A0(net31),
    .A1(_0153_),
    .S(_0731_),
    .Y(_0154_));
 sky130_fd_sc_hd__nor2_1 _1547_ (.A(\y[6] ),
    .B(_0112_),
    .Y(_0155_));
 sky130_fd_sc_hd__a21oi_1 _1548_ (.A1(_0145_),
    .A2(_0154_),
    .B1(_0155_),
    .Y(_0051_));
 sky130_fd_sc_hd__a21o_1 _1549_ (.A1(_0832_),
    .A2(_0147_),
    .B1(_0831_),
    .X(_0156_));
 sky130_fd_sc_hd__a21oi_1 _1550_ (.A1(_0835_),
    .A2(_0156_),
    .B1(_0834_),
    .Y(_0157_));
 sky130_fd_sc_hd__xnor2_1 _1551_ (.A(_0838_),
    .B(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__mux2i_1 _1552_ (.A0(net32),
    .A1(_0158_),
    .S(_0731_),
    .Y(_0159_));
 sky130_fd_sc_hd__nor2_1 _1553_ (.A(\y[7] ),
    .B(_0112_),
    .Y(_0160_));
 sky130_fd_sc_hd__a21oi_1 _1554_ (.A1(_0145_),
    .A2(_0159_),
    .B1(_0160_),
    .Y(_0052_));
 sky130_fd_sc_hd__nor2_1 _1555_ (.A(_0700_),
    .B(_0704_),
    .Y(_0161_));
 sky130_fd_sc_hd__nor2_1 _1556_ (.A(_0837_),
    .B(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__xnor2_1 _1557_ (.A(_0841_),
    .B(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__mux2i_1 _1558_ (.A0(net33),
    .A1(_0163_),
    .S(_0731_),
    .Y(_0164_));
 sky130_fd_sc_hd__nor2_1 _1559_ (.A(\y[8] ),
    .B(_0112_),
    .Y(_0165_));
 sky130_fd_sc_hd__a21oi_1 _1560_ (.A1(_0145_),
    .A2(_0164_),
    .B1(_0165_),
    .Y(_0053_));
 sky130_fd_sc_hd__o21bai_1 _1561_ (.A1(_0712_),
    .A2(_0718_),
    .B1_N(_0837_),
    .Y(_0166_));
 sky130_fd_sc_hd__a21oi_1 _1562_ (.A1(_0841_),
    .A2(_0166_),
    .B1(_0840_),
    .Y(_0167_));
 sky130_fd_sc_hd__xnor2_1 _1563_ (.A(_0844_),
    .B(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__mux2i_1 _1564_ (.A0(net34),
    .A1(_0168_),
    .S(_0731_),
    .Y(_0169_));
 sky130_fd_sc_hd__nor2_1 _1565_ (.A(\y[9] ),
    .B(_0112_),
    .Y(_0170_));
 sky130_fd_sc_hd__a21oi_1 _1566_ (.A1(_0145_),
    .A2(_0169_),
    .B1(_0170_),
    .Y(_0054_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(net68),
    .A1(\y[0] ),
    .S(_0696_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1568_ (.A0(net69),
    .A1(\y[10] ),
    .S(_0696_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _1569_ (.A0(net70),
    .A1(\y[11] ),
    .S(_0696_),
    .X(_0057_));
 sky130_fd_sc_hd__clkbuf_4 _1570_ (.A(_0916_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _1571_ (.A0(net71),
    .A1(\y[12] ),
    .S(_0171_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _1572_ (.A0(net72),
    .A1(\y[13] ),
    .S(_0171_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _1573_ (.A0(net73),
    .A1(\y[14] ),
    .S(_0171_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1574_ (.A0(net74),
    .A1(_0425_),
    .S(_0171_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1575_ (.A0(net75),
    .A1(\y[1] ),
    .S(_0171_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1576_ (.A0(net76),
    .A1(\y[2] ),
    .S(_0171_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1577_ (.A0(net77),
    .A1(\y[3] ),
    .S(_0171_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1578_ (.A0(net78),
    .A1(\y[4] ),
    .S(_0171_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1579_ (.A0(net79),
    .A1(\y[5] ),
    .S(_0171_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1580_ (.A0(net80),
    .A1(\y[6] ),
    .S(_0171_),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_4 _1581_ (.A(_0916_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _1582_ (.A0(net81),
    .A1(\y[7] ),
    .S(_0172_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1583_ (.A0(net82),
    .A1(\y[8] ),
    .S(_0172_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1584_ (.A0(net83),
    .A1(\y[9] ),
    .S(_0172_),
    .X(_0070_));
 sky130_fd_sc_hd__buf_4 _1585_ (.A(_0562_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2i_1 _1586_ (.A0(net35),
    .A1(_0747_),
    .S(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__nor2_1 _1587_ (.A(_0565_),
    .B(\z[0] ),
    .Y(_0175_));
 sky130_fd_sc_hd__a21oi_1 _1588_ (.A1(_0145_),
    .A2(_0174_),
    .B1(_0175_),
    .Y(_0071_));
 sky130_fd_sc_hd__a21o_1 _1589_ (.A1(_0735_),
    .A2(_0756_),
    .B1(_0755_),
    .X(_0176_));
 sky130_fd_sc_hd__a21o_1 _1590_ (.A1(_0759_),
    .A2(_0176_),
    .B1(_0758_),
    .X(_0177_));
 sky130_fd_sc_hd__or3_1 _1591_ (.A(_0761_),
    .B(_0782_),
    .C(_0785_),
    .X(_0178_));
 sky130_fd_sc_hd__a21oi_1 _1592_ (.A1(_0762_),
    .A2(_0177_),
    .B1(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__or2_0 _1593_ (.A(_0783_),
    .B(_0782_),
    .X(_0180_));
 sky130_fd_sc_hd__a21oi_1 _1594_ (.A1(_0786_),
    .A2(_0180_),
    .B1(_0785_),
    .Y(_0181_));
 sky130_fd_sc_hd__and2_0 _1595_ (.A(_0789_),
    .B(_0792_),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _1596_ (.A(_0795_),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__a21oi_1 _1597_ (.A1(_0792_),
    .A2(_0788_),
    .B1(_0791_),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_1 _1598_ (.A(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__a21oi_1 _1599_ (.A1(_0795_),
    .A2(_0185_),
    .B1(_0794_),
    .Y(_0186_));
 sky130_fd_sc_hd__o31ai_2 _1600_ (.A1(_0179_),
    .A2(_0181_),
    .A3(_0183_),
    .B1(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__xnor2_1 _1601_ (.A(_0798_),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__nor2_1 _1602_ (.A(_0569_),
    .B(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__a21oi_1 _1603_ (.A1(_0569_),
    .A2(net36),
    .B1(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__nor2_1 _1604_ (.A(_0565_),
    .B(\z[10] ),
    .Y(_0191_));
 sky130_fd_sc_hd__a21oi_1 _1605_ (.A1(_0145_),
    .A2(_0190_),
    .B1(_0191_),
    .Y(_0072_));
 sky130_fd_sc_hd__a21o_1 _1606_ (.A1(_0733_),
    .A2(_0753_),
    .B1(_0752_),
    .X(_0192_));
 sky130_fd_sc_hd__nand2_1 _1607_ (.A(_0756_),
    .B(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__nor2_1 _1608_ (.A(_0755_),
    .B(_0758_),
    .Y(_0194_));
 sky130_fd_sc_hd__o21ai_0 _1609_ (.A1(_0759_),
    .A2(_0758_),
    .B1(_0762_),
    .Y(_0195_));
 sky130_fd_sc_hd__a21oi_1 _1610_ (.A1(_0193_),
    .A2(_0194_),
    .B1(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__o21ba_1 _1611_ (.A1(_0178_),
    .A2(_0196_),
    .B1_N(_0181_),
    .X(_0197_));
 sky130_fd_sc_hd__nand2_1 _1612_ (.A(_0795_),
    .B(_0798_),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2_1 _1613_ (.A(_0798_),
    .B(_0794_),
    .Y(_0199_));
 sky130_fd_sc_hd__o21ai_0 _1614_ (.A1(_0184_),
    .A2(_0198_),
    .B1(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__a41oi_2 _1615_ (.A1(_0795_),
    .A2(_0798_),
    .A3(_0182_),
    .A4(_0197_),
    .B1(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__nor2b_1 _1616_ (.A(_0797_),
    .B_N(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__xnor2_1 _1617_ (.A(_0801_),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__mux2i_1 _1618_ (.A0(net37),
    .A1(_0203_),
    .S(_0173_),
    .Y(_0204_));
 sky130_fd_sc_hd__nor2_1 _1619_ (.A(_0565_),
    .B(\z[11] ),
    .Y(_0205_));
 sky130_fd_sc_hd__a21oi_1 _1620_ (.A1(_0145_),
    .A2(_0204_),
    .B1(_0205_),
    .Y(_0073_));
 sky130_fd_sc_hd__nand3_1 _1621_ (.A(_0798_),
    .B(_0801_),
    .C(_0187_),
    .Y(_0206_));
 sky130_fd_sc_hd__nand2_1 _1622_ (.A(_0801_),
    .B(_0797_),
    .Y(_0207_));
 sky130_fd_sc_hd__and3b_1 _1623_ (.A_N(_0800_),
    .B(_0206_),
    .C(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__xnor2_1 _1624_ (.A(_0804_),
    .B(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__mux2i_1 _1625_ (.A0(net38),
    .A1(_0209_),
    .S(_0173_),
    .Y(_0210_));
 sky130_fd_sc_hd__nor2_1 _1626_ (.A(_0565_),
    .B(\z[12] ),
    .Y(_0211_));
 sky130_fd_sc_hd__a21oi_1 _1627_ (.A1(_0145_),
    .A2(_0210_),
    .B1(_0211_),
    .Y(_0074_));
 sky130_fd_sc_hd__nor3_1 _1628_ (.A(_0797_),
    .B(_0800_),
    .C(_0803_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor3_1 _1629_ (.A(_0801_),
    .B(_0800_),
    .C(_0803_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor2_1 _1630_ (.A(_0804_),
    .B(_0803_),
    .Y(_0214_));
 sky130_fd_sc_hd__a211o_1 _1631_ (.A1(_0201_),
    .A2(_0212_),
    .B1(_0213_),
    .C1(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__xnor2_1 _1632_ (.A(_0807_),
    .B(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__mux2i_1 _1633_ (.A0(net39),
    .A1(_0216_),
    .S(_0173_),
    .Y(_0217_));
 sky130_fd_sc_hd__nor2_1 _1634_ (.A(_0565_),
    .B(\z[13] ),
    .Y(_0218_));
 sky130_fd_sc_hd__a21oi_1 _1635_ (.A1(_0145_),
    .A2(_0217_),
    .B1(_0218_),
    .Y(_0075_));
 sky130_fd_sc_hd__nor3_1 _1636_ (.A(_0800_),
    .B(_0803_),
    .C(_0806_),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_1 _1637_ (.A(_0214_),
    .Y(_0220_));
 sky130_fd_sc_hd__a21oi_1 _1638_ (.A1(_0807_),
    .A2(_0220_),
    .B1(_0806_),
    .Y(_0221_));
 sky130_fd_sc_hd__a31oi_1 _1639_ (.A1(_0206_),
    .A2(_0207_),
    .A3(_0219_),
    .B1(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__xor2_1 _1640_ (.A(_0810_),
    .B(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2i_1 _1641_ (.A0(net40),
    .A1(_0223_),
    .S(_0173_),
    .Y(_0224_));
 sky130_fd_sc_hd__nor2_1 _1642_ (.A(_0565_),
    .B(\z[14] ),
    .Y(_0225_));
 sky130_fd_sc_hd__a21oi_1 _1643_ (.A1(_0561_),
    .A2(_0224_),
    .B1(_0225_),
    .Y(_0076_));
 sky130_fd_sc_hd__nand2_1 _1644_ (.A(_0807_),
    .B(_0810_),
    .Y(_0226_));
 sky130_fd_sc_hd__a21oi_1 _1645_ (.A1(_0810_),
    .A2(_0806_),
    .B1(_0809_),
    .Y(_0227_));
 sky130_fd_sc_hd__o21ai_0 _1646_ (.A1(_0215_),
    .A2(_0226_),
    .B1(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__o21ai_0 _1647_ (.A1(_0765_),
    .A2(_0769_),
    .B1(_0377_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand3_1 _1648_ (.A(_0364_),
    .B(_0527_),
    .C(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__xnor2_1 _1649_ (.A(_0228_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__nand3_1 _1650_ (.A(_0569_),
    .B(net41),
    .C(_0574_),
    .Y(_0232_));
 sky130_fd_sc_hd__o221ai_1 _1651_ (.A1(_0364_),
    .A2(_0112_),
    .B1(_0563_),
    .B2(_0231_),
    .C1(_0232_),
    .Y(_0077_));
 sky130_fd_sc_hd__nor2_1 _1652_ (.A(_0578_),
    .B(net42),
    .Y(_0233_));
 sky130_fd_sc_hd__a21oi_1 _1653_ (.A1(_0578_),
    .A2(_0736_),
    .B1(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__mux2_1 _1654_ (.A0(\z[1] ),
    .A1(_0234_),
    .S(_0570_),
    .X(_0078_));
 sky130_fd_sc_hd__xnor2_1 _1655_ (.A(_0735_),
    .B(_0756_),
    .Y(_0235_));
 sky130_fd_sc_hd__nor2_1 _1656_ (.A(_0562_),
    .B(net43),
    .Y(_0236_));
 sky130_fd_sc_hd__a21oi_1 _1657_ (.A1(_0578_),
    .A2(_0235_),
    .B1(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__mux2_1 _1658_ (.A0(\z[2] ),
    .A1(_0237_),
    .S(_0570_),
    .X(_0079_));
 sky130_fd_sc_hd__a21oi_1 _1659_ (.A1(_0756_),
    .A2(_0192_),
    .B1(_0755_),
    .Y(_0238_));
 sky130_fd_sc_hd__xnor2_1 _1660_ (.A(_0759_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__mux2i_1 _1661_ (.A0(net44),
    .A1(_0239_),
    .S(_0173_),
    .Y(_0240_));
 sky130_fd_sc_hd__nor2_1 _1662_ (.A(_0565_),
    .B(\z[3] ),
    .Y(_0241_));
 sky130_fd_sc_hd__a21oi_1 _1663_ (.A1(_0561_),
    .A2(_0240_),
    .B1(_0241_),
    .Y(_0080_));
 sky130_fd_sc_hd__xor2_1 _1664_ (.A(_0762_),
    .B(_0177_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2i_1 _1665_ (.A0(net45),
    .A1(_0242_),
    .S(_0173_),
    .Y(_0243_));
 sky130_fd_sc_hd__nor2_1 _1666_ (.A(_0565_),
    .B(\z[4] ),
    .Y(_0244_));
 sky130_fd_sc_hd__a21oi_1 _1667_ (.A1(_0561_),
    .A2(_0243_),
    .B1(_0244_),
    .Y(_0081_));
 sky130_fd_sc_hd__nor2_1 _1668_ (.A(_0761_),
    .B(_0196_),
    .Y(_0245_));
 sky130_fd_sc_hd__xnor2_1 _1669_ (.A(_0783_),
    .B(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__mux2i_1 _1670_ (.A0(net46),
    .A1(_0246_),
    .S(_0173_),
    .Y(_0247_));
 sky130_fd_sc_hd__nor2_1 _1671_ (.A(_0574_),
    .B(\z[5] ),
    .Y(_0248_));
 sky130_fd_sc_hd__a21oi_1 _1672_ (.A1(_0561_),
    .A2(_0247_),
    .B1(_0248_),
    .Y(_0082_));
 sky130_fd_sc_hd__a21o_1 _1673_ (.A1(_0762_),
    .A2(_0177_),
    .B1(_0761_),
    .X(_0249_));
 sky130_fd_sc_hd__a21oi_1 _1674_ (.A1(_0783_),
    .A2(_0249_),
    .B1(_0782_),
    .Y(_0250_));
 sky130_fd_sc_hd__xnor2_1 _1675_ (.A(_0786_),
    .B(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__mux2i_1 _1676_ (.A0(net47),
    .A1(_0251_),
    .S(_0173_),
    .Y(_0252_));
 sky130_fd_sc_hd__nor2_1 _1677_ (.A(_0574_),
    .B(\z[6] ),
    .Y(_0253_));
 sky130_fd_sc_hd__a21oi_1 _1678_ (.A1(_0561_),
    .A2(_0252_),
    .B1(_0253_),
    .Y(_0083_));
 sky130_fd_sc_hd__xor2_1 _1679_ (.A(_0789_),
    .B(_0197_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2i_1 _1680_ (.A0(net48),
    .A1(_0254_),
    .S(_0173_),
    .Y(_0255_));
 sky130_fd_sc_hd__nor2_1 _1681_ (.A(_0574_),
    .B(\z[7] ),
    .Y(_0256_));
 sky130_fd_sc_hd__a21oi_1 _1682_ (.A1(_0561_),
    .A2(_0255_),
    .B1(_0256_),
    .Y(_0084_));
 sky130_fd_sc_hd__nor2_1 _1683_ (.A(_0179_),
    .B(_0181_),
    .Y(_0257_));
 sky130_fd_sc_hd__a21oi_1 _1684_ (.A1(_0789_),
    .A2(_0257_),
    .B1(_0788_),
    .Y(_0258_));
 sky130_fd_sc_hd__xnor2_1 _1685_ (.A(_0792_),
    .B(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__mux2i_1 _1686_ (.A0(net49),
    .A1(_0259_),
    .S(_0578_),
    .Y(_0260_));
 sky130_fd_sc_hd__nor2_1 _1687_ (.A(_0574_),
    .B(\z[8] ),
    .Y(_0261_));
 sky130_fd_sc_hd__a21oi_1 _1688_ (.A1(_0561_),
    .A2(_0260_),
    .B1(_0261_),
    .Y(_0085_));
 sky130_fd_sc_hd__a21o_1 _1689_ (.A1(_0182_),
    .A2(_0197_),
    .B1(_0185_),
    .X(_0262_));
 sky130_fd_sc_hd__xor2_1 _1690_ (.A(_0795_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2i_1 _1691_ (.A0(net50),
    .A1(_0263_),
    .S(_0578_),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2_1 _1692_ (.A(_0574_),
    .B(\z[9] ),
    .Y(_0265_));
 sky130_fd_sc_hd__a21oi_1 _1693_ (.A1(_0561_),
    .A2(_0264_),
    .B1(_0265_),
    .Y(_0086_));
 sky130_fd_sc_hd__mux2_1 _1694_ (.A0(net84),
    .A1(\z[0] ),
    .S(_0172_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1695_ (.A0(net85),
    .A1(\z[10] ),
    .S(_0172_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(net86),
    .A1(\z[11] ),
    .S(_0172_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1697_ (.A0(net87),
    .A1(\z[12] ),
    .S(_0172_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _1698_ (.A0(net88),
    .A1(\z[13] ),
    .S(_0172_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1699_ (.A0(net89),
    .A1(\z[14] ),
    .S(_0172_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _1700_ (.A0(net90),
    .A1(_0302_),
    .S(_0172_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1701_ (.A0(net91),
    .A1(\z[1] ),
    .S(_0694_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _1702_ (.A0(net92),
    .A1(\z[2] ),
    .S(_0694_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _1703_ (.A0(net93),
    .A1(\z[3] ),
    .S(_0694_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(net94),
    .A1(\z[4] ),
    .S(_0694_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _1705_ (.A0(net95),
    .A1(\z[5] ),
    .S(_0694_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _1706_ (.A0(net96),
    .A1(\z[6] ),
    .S(_0694_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _1707_ (.A0(net97),
    .A1(\z[7] ),
    .S(_0694_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _1708_ (.A0(net98),
    .A1(\z[8] ),
    .S(_0694_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1709_ (.A0(net99),
    .A1(\z[9] ),
    .S(_0694_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1710_ (.A0(_0695_),
    .A1(net51),
    .S(_0560_),
    .X(_0000_));
 sky130_fd_sc_hd__fa_1 _1711_ (.A(\z[1] ),
    .B(_0733_),
    .CIN(_0734_),
    .COUT(_0735_),
    .SUM(_0736_));
 sky130_fd_sc_hd__fa_1 _1712_ (.A(\y[1] ),
    .B(_0737_),
    .CIN(_0738_),
    .COUT(_0739_),
    .SUM(_0740_));
 sky130_fd_sc_hd__fa_1 _1713_ (.A(_0741_),
    .B(_0742_),
    .CIN(_0743_),
    .COUT(_0744_),
    .SUM(_0745_));
 sky130_fd_sc_hd__ha_1 _1714_ (.A(\z[0] ),
    .B(_0746_),
    .COUT(_0733_),
    .SUM(_0747_));
 sky130_fd_sc_hd__ha_1 _1715_ (.A(_0748_),
    .B(_0749_),
    .COUT(_0750_),
    .SUM(_0751_));
 sky130_fd_sc_hd__ha_1 _1716_ (.A(\z[1] ),
    .B(_0734_),
    .COUT(_0752_),
    .SUM(_0753_));
 sky130_fd_sc_hd__ha_1 _1717_ (.A(\z[2] ),
    .B(_0754_),
    .COUT(_0755_),
    .SUM(_0756_));
 sky130_fd_sc_hd__ha_1 _1718_ (.A(\z[3] ),
    .B(_0757_),
    .COUT(_0758_),
    .SUM(_0759_));
 sky130_fd_sc_hd__ha_1 _1719_ (.A(\z[4] ),
    .B(_0760_),
    .COUT(_0761_),
    .SUM(_0762_));
 sky130_fd_sc_hd__ha_1 _1720_ (.A(_0763_),
    .B(_0764_),
    .COUT(_0765_),
    .SUM(_0766_));
 sky130_fd_sc_hd__ha_1 _1721_ (.A(_0763_),
    .B(_0764_),
    .COUT(_0767_),
    .SUM(_0768_));
 sky130_fd_sc_hd__ha_1 _1722_ (.A(_0763_),
    .B(net103),
    .COUT(_0769_),
    .SUM(_0770_));
 sky130_fd_sc_hd__ha_1 _1723_ (.A(_0763_),
    .B(net103),
    .COUT(_0771_),
    .SUM(_0772_));
 sky130_fd_sc_hd__ha_2 _1724_ (.A(\iteration[0] ),
    .B(_0764_),
    .COUT(_0773_),
    .SUM(_0774_));
 sky130_fd_sc_hd__ha_1 _1725_ (.A(\iteration[0] ),
    .B(_0764_),
    .COUT(_0775_),
    .SUM(_0776_));
 sky130_fd_sc_hd__ha_1 _1726_ (.A(\iteration[0] ),
    .B(net103),
    .COUT(_0777_),
    .SUM(_0778_));
 sky130_fd_sc_hd__ha_1 _1727_ (.A(\iteration[0] ),
    .B(net103),
    .COUT(_0779_),
    .SUM(_0780_));
 sky130_fd_sc_hd__ha_1 _1728_ (.A(\z[5] ),
    .B(_0781_),
    .COUT(_0782_),
    .SUM(_0783_));
 sky130_fd_sc_hd__ha_1 _1729_ (.A(\z[6] ),
    .B(_0784_),
    .COUT(_0785_),
    .SUM(_0786_));
 sky130_fd_sc_hd__ha_1 _1730_ (.A(\z[7] ),
    .B(_0787_),
    .COUT(_0788_),
    .SUM(_0789_));
 sky130_fd_sc_hd__ha_1 _1731_ (.A(\z[8] ),
    .B(_0790_),
    .COUT(_0791_),
    .SUM(_0792_));
 sky130_fd_sc_hd__ha_1 _1732_ (.A(\z[9] ),
    .B(_0793_),
    .COUT(_0794_),
    .SUM(_0795_));
 sky130_fd_sc_hd__ha_1 _1733_ (.A(\z[10] ),
    .B(_0796_),
    .COUT(_0797_),
    .SUM(_0798_));
 sky130_fd_sc_hd__ha_1 _1734_ (.A(\z[11] ),
    .B(_0799_),
    .COUT(_0800_),
    .SUM(_0801_));
 sky130_fd_sc_hd__ha_1 _1735_ (.A(\z[12] ),
    .B(_0802_),
    .COUT(_0803_),
    .SUM(_0804_));
 sky130_fd_sc_hd__ha_1 _1736_ (.A(\z[13] ),
    .B(_0805_),
    .COUT(_0806_),
    .SUM(_0807_));
 sky130_fd_sc_hd__ha_1 _1737_ (.A(\z[14] ),
    .B(_0808_),
    .COUT(_0809_),
    .SUM(_0810_));
 sky130_fd_sc_hd__ha_1 _1738_ (.A(_0811_),
    .B(_0812_),
    .COUT(_0813_),
    .SUM(_0814_));
 sky130_fd_sc_hd__ha_1 _1739_ (.A(_0815_),
    .B(_0816_),
    .COUT(_0817_),
    .SUM(_0818_));
 sky130_fd_sc_hd__ha_1 _1740_ (.A(\y[1] ),
    .B(_0738_),
    .COUT(_0819_),
    .SUM(_0820_));
 sky130_fd_sc_hd__ha_1 _1741_ (.A(\y[2] ),
    .B(_0821_),
    .COUT(_0822_),
    .SUM(_0823_));
 sky130_fd_sc_hd__ha_1 _1742_ (.A(\y[3] ),
    .B(_0824_),
    .COUT(_0825_),
    .SUM(_0826_));
 sky130_fd_sc_hd__ha_1 _1743_ (.A(\y[4] ),
    .B(_0827_),
    .COUT(_0828_),
    .SUM(_0829_));
 sky130_fd_sc_hd__ha_1 _1744_ (.A(\y[5] ),
    .B(_0830_),
    .COUT(_0831_),
    .SUM(_0832_));
 sky130_fd_sc_hd__ha_1 _1745_ (.A(\y[6] ),
    .B(_0833_),
    .COUT(_0834_),
    .SUM(_0835_));
 sky130_fd_sc_hd__ha_1 _1746_ (.A(\y[7] ),
    .B(_0836_),
    .COUT(_0837_),
    .SUM(_0838_));
 sky130_fd_sc_hd__ha_1 _1747_ (.A(\y[8] ),
    .B(_0839_),
    .COUT(_0840_),
    .SUM(_0841_));
 sky130_fd_sc_hd__ha_1 _1748_ (.A(\y[9] ),
    .B(_0842_),
    .COUT(_0843_),
    .SUM(_0844_));
 sky130_fd_sc_hd__ha_1 _1749_ (.A(\y[10] ),
    .B(_0845_),
    .COUT(_0846_),
    .SUM(_0847_));
 sky130_fd_sc_hd__ha_1 _1750_ (.A(\y[11] ),
    .B(_0848_),
    .COUT(_0849_),
    .SUM(_0850_));
 sky130_fd_sc_hd__ha_1 _1751_ (.A(\y[12] ),
    .B(_0851_),
    .COUT(_0852_),
    .SUM(_0853_));
 sky130_fd_sc_hd__ha_1 _1752_ (.A(\y[13] ),
    .B(_0854_),
    .COUT(_0855_),
    .SUM(_0856_));
 sky130_fd_sc_hd__ha_1 _1753_ (.A(\y[14] ),
    .B(_0857_),
    .COUT(_0858_),
    .SUM(_0859_));
 sky130_fd_sc_hd__ha_1 _1754_ (.A(\x[0] ),
    .B(_0860_),
    .COUT(_0861_),
    .SUM(_0862_));
 sky130_fd_sc_hd__ha_1 _1755_ (.A(_0863_),
    .B(_0864_),
    .COUT(_0865_),
    .SUM(_0866_));
 sky130_fd_sc_hd__ha_1 _1756_ (.A(\x[1] ),
    .B(_0867_),
    .COUT(_0868_),
    .SUM(_0869_));
 sky130_fd_sc_hd__ha_1 _1757_ (.A(\x[2] ),
    .B(_0870_),
    .COUT(_0871_),
    .SUM(_0872_));
 sky130_fd_sc_hd__ha_1 _1758_ (.A(\x[3] ),
    .B(_0873_),
    .COUT(_0874_),
    .SUM(_0875_));
 sky130_fd_sc_hd__ha_1 _1759_ (.A(\x[4] ),
    .B(_0876_),
    .COUT(_0877_),
    .SUM(_0878_));
 sky130_fd_sc_hd__ha_1 _1760_ (.A(\x[5] ),
    .B(_0879_),
    .COUT(_0880_),
    .SUM(_0881_));
 sky130_fd_sc_hd__ha_1 _1761_ (.A(\x[6] ),
    .B(_0882_),
    .COUT(_0883_),
    .SUM(_0884_));
 sky130_fd_sc_hd__ha_1 _1762_ (.A(\x[7] ),
    .B(_0885_),
    .COUT(_0886_),
    .SUM(_0887_));
 sky130_fd_sc_hd__ha_1 _1763_ (.A(\x[8] ),
    .B(_0888_),
    .COUT(_0889_),
    .SUM(_0890_));
 sky130_fd_sc_hd__ha_1 _1764_ (.A(_0891_),
    .B(\x[9] ),
    .COUT(_0892_),
    .SUM(_0893_));
 sky130_fd_sc_hd__ha_1 _1765_ (.A(\x[10] ),
    .B(_0894_),
    .COUT(_0895_),
    .SUM(_0896_));
 sky130_fd_sc_hd__ha_1 _1766_ (.A(\x[11] ),
    .B(_0897_),
    .COUT(_0898_),
    .SUM(_0899_));
 sky130_fd_sc_hd__ha_1 _1767_ (.A(_0900_),
    .B(\x[12] ),
    .COUT(_0901_),
    .SUM(_0902_));
 sky130_fd_sc_hd__ha_1 _1768_ (.A(_0903_),
    .B(\x[13] ),
    .COUT(_0904_),
    .SUM(_0905_));
 sky130_fd_sc_hd__ha_1 _1769_ (.A(\x[14] ),
    .B(_0906_),
    .COUT(_0907_),
    .SUM(_0908_));
 sky130_fd_sc_hd__ha_1 _1770_ (.A(_0909_),
    .B(_0910_),
    .COUT(_0911_),
    .SUM(\next_state[1] ));
 sky130_fd_sc_hd__ha_1 _1771_ (.A(_0909_),
    .B(_0910_),
    .COUT(_0912_),
    .SUM(_0913_));
 sky130_fd_sc_hd__ha_1 _1772_ (.A(_0909_),
    .B(\state[1] ),
    .COUT(_0914_),
    .SUM(_0915_));
 sky130_fd_sc_hd__ha_2 _1773_ (.A(\state[0] ),
    .B(\state[1] ),
    .COUT(_0916_),
    .SUM(_0917_));
 sky130_fd_sc_hd__dfrtp_1 \done$_DFFE_PN0P_  (.D(_0000_),
    .Q(net51),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \iteration[0]$_DFFE_PN0P_  (.D(_0001_),
    .Q(\iteration[0] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \iteration[1]$_DFFE_PN0P_  (.D(_0002_),
    .Q(\iteration[1] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \iteration[2]$_DFFE_PN0P_  (.D(_0003_),
    .Q(\iteration[2] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \iteration[3]$_DFFE_PN0P_  (.D(_0004_),
    .Q(\iteration[3] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[0]$_DFFE_PN0P_  (.D(_0005_),
    .Q(\state[0] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[1]$_DFFE_PN0P_  (.D(_0006_),
    .Q(\state[1] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x[0]$_DFFE_PN0P_  (.D(_0007_),
    .Q(\x[0] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[10]$_DFFE_PN0P_  (.D(_0008_),
    .Q(\x[10] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[11]$_DFFE_PN0P_  (.D(_0009_),
    .Q(\x[11] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[12]$_DFFE_PN0P_  (.D(_0010_),
    .Q(\x[12] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[13]$_DFFE_PN0P_  (.D(_0011_),
    .Q(\x[13] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[14]$_DFFE_PN0P_  (.D(_0012_),
    .Q(\x[14] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[15]$_DFFE_PN0P_  (.D(_0013_),
    .Q(\x[15] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \x[1]$_DFFE_PN0P_  (.D(_0014_),
    .Q(\x[1] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \x[2]$_DFFE_PN0P_  (.D(_0015_),
    .Q(\x[2] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[3]$_DFFE_PN0P_  (.D(_0016_),
    .Q(\x[3] ),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \x[4]$_DFFE_PN0P_  (.D(_0017_),
    .Q(\x[4] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \x[5]$_DFFE_PN0P_  (.D(_0018_),
    .Q(\x[5] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \x[6]$_DFFE_PN0P_  (.D(_0019_),
    .Q(\x[6] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[7]$_DFFE_PN0P_  (.D(_0020_),
    .Q(\x[7] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[8]$_DFFE_PN0P_  (.D(_0021_),
    .Q(\x[8] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \x[9]$_DFFE_PN0P_  (.D(_0022_),
    .Q(\x[9] ),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[0]$_DFFE_PN0P_  (.D(_0023_),
    .Q(net52),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[10]$_DFFE_PN0P_  (.D(_0024_),
    .Q(net53),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[11]$_DFFE_PN0P_  (.D(_0025_),
    .Q(net54),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[12]$_DFFE_PN0P_  (.D(_0026_),
    .Q(net55),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[13]$_DFFE_PN0P_  (.D(_0027_),
    .Q(net56),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[14]$_DFFE_PN0P_  (.D(_0028_),
    .Q(net57),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[15]$_DFFE_PN0P_  (.D(_0029_),
    .Q(net58),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[1]$_DFFE_PN0P_  (.D(_0030_),
    .Q(net59),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[2]$_DFFE_PN0P_  (.D(_0031_),
    .Q(net60),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[3]$_DFFE_PN0P_  (.D(_0032_),
    .Q(net61),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[4]$_DFFE_PN0P_  (.D(_0033_),
    .Q(net62),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[5]$_DFFE_PN0P_  (.D(_0034_),
    .Q(net63),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[6]$_DFFE_PN0P_  (.D(_0035_),
    .Q(net64),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[7]$_DFFE_PN0P_  (.D(_0036_),
    .Q(net65),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[8]$_DFFE_PN0P_  (.D(_0037_),
    .Q(net66),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \x_out[9]$_DFFE_PN0P_  (.D(_0038_),
    .Q(net67),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \y[0]$_DFFE_PN0P_  (.D(_0039_),
    .Q(\y[0] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \y[10]$_DFFE_PN0P_  (.D(_0040_),
    .Q(\y[10] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \y[11]$_DFFE_PN0P_  (.D(_0041_),
    .Q(\y[11] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \y[12]$_DFFE_PN0P_  (.D(_0042_),
    .Q(\y[12] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \y[13]$_DFFE_PN0P_  (.D(_0043_),
    .Q(\y[13] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \y[14]$_DFFE_PN0P_  (.D(_0044_),
    .Q(\y[14] ),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y[15]$_DFFE_PN0P_  (.D(_0045_),
    .Q(\y[15] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \y[1]$_DFFE_PN0P_  (.D(_0046_),
    .Q(\y[1] ),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \y[2]$_DFFE_PN0P_  (.D(_0047_),
    .Q(\y[2] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \y[3]$_DFFE_PN0P_  (.D(_0048_),
    .Q(\y[3] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \y[4]$_DFFE_PN0P_  (.D(_0049_),
    .Q(\y[4] ),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \y[5]$_DFFE_PN0P_  (.D(_0050_),
    .Q(\y[5] ),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \y[6]$_DFFE_PN0P_  (.D(_0051_),
    .Q(\y[6] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \y[7]$_DFFE_PN0P_  (.D(_0052_),
    .Q(\y[7] ),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \y[8]$_DFFE_PN0P_  (.D(_0053_),
    .Q(\y[8] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \y[9]$_DFFE_PN0P_  (.D(_0054_),
    .Q(\y[9] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[0]$_DFFE_PN0P_  (.D(_0055_),
    .Q(net68),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[10]$_DFFE_PN0P_  (.D(_0056_),
    .Q(net69),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[11]$_DFFE_PN0P_  (.D(_0057_),
    .Q(net70),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[12]$_DFFE_PN0P_  (.D(_0058_),
    .Q(net71),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[13]$_DFFE_PN0P_  (.D(_0059_),
    .Q(net72),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[14]$_DFFE_PN0P_  (.D(_0060_),
    .Q(net73),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[15]$_DFFE_PN0P_  (.D(_0061_),
    .Q(net74),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[1]$_DFFE_PN0P_  (.D(_0062_),
    .Q(net75),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[2]$_DFFE_PN0P_  (.D(_0063_),
    .Q(net76),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[3]$_DFFE_PN0P_  (.D(_0064_),
    .Q(net77),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[4]$_DFFE_PN0P_  (.D(_0065_),
    .Q(net78),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[5]$_DFFE_PN0P_  (.D(_0066_),
    .Q(net79),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[6]$_DFFE_PN0P_  (.D(_0067_),
    .Q(net80),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[7]$_DFFE_PN0P_  (.D(_0068_),
    .Q(net81),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[8]$_DFFE_PN0P_  (.D(_0069_),
    .Q(net82),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \y_out[9]$_DFFE_PN0P_  (.D(_0070_),
    .Q(net83),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[0]$_DFFE_PN0P_  (.D(_0071_),
    .Q(\z[0] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[10]$_DFFE_PN0P_  (.D(_0072_),
    .Q(\z[10] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[11]$_DFFE_PN0P_  (.D(_0073_),
    .Q(\z[11] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[12]$_DFFE_PN0P_  (.D(_0074_),
    .Q(\z[12] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[13]$_DFFE_PN0P_  (.D(_0075_),
    .Q(\z[13] ),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[14]$_DFFE_PN0P_  (.D(_0076_),
    .Q(\z[14] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[15]$_DFFE_PN0P_  (.D(_0077_),
    .Q(\z[15] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[1]$_DFFE_PN0P_  (.D(_0078_),
    .Q(\z[1] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[2]$_DFFE_PN0P_  (.D(_0079_),
    .Q(\z[2] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[3]$_DFFE_PN0P_  (.D(_0080_),
    .Q(\z[3] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[4]$_DFFE_PN0P_  (.D(_0081_),
    .Q(\z[4] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[5]$_DFFE_PN0P_  (.D(_0082_),
    .Q(\z[5] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[6]$_DFFE_PN0P_  (.D(_0083_),
    .Q(\z[6] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[7]$_DFFE_PN0P_  (.D(_0084_),
    .Q(\z[7] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[8]$_DFFE_PN0P_  (.D(_0085_),
    .Q(\z[8] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z[9]$_DFFE_PN0P_  (.D(_0086_),
    .Q(\z[9] ),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[0]$_DFFE_PN0P_  (.D(_0087_),
    .Q(net84),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[10]$_DFFE_PN0P_  (.D(_0088_),
    .Q(net85),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[11]$_DFFE_PN0P_  (.D(_0089_),
    .Q(net86),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[12]$_DFFE_PN0P_  (.D(_0090_),
    .Q(net87),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[13]$_DFFE_PN0P_  (.D(_0091_),
    .Q(net88),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[14]$_DFFE_PN0P_  (.D(_0092_),
    .Q(net89),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[15]$_DFFE_PN0P_  (.D(_0093_),
    .Q(net90),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[1]$_DFFE_PN0P_  (.D(_0094_),
    .Q(net91),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[2]$_DFFE_PN0P_  (.D(_0095_),
    .Q(net92),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[3]$_DFFE_PN0P_  (.D(_0096_),
    .Q(net93),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[4]$_DFFE_PN0P_  (.D(_0097_),
    .Q(net94),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[5]$_DFFE_PN0P_  (.D(_0098_),
    .Q(net95),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[6]$_DFFE_PN0P_  (.D(_0099_),
    .Q(net96),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[7]$_DFFE_PN0P_  (.D(_0100_),
    .Q(net97),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[8]$_DFFE_PN0P_  (.D(_0101_),
    .Q(net98),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \z_out[9]$_DFFE_PN0P_  (.D(_0102_),
    .Q(net99),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net100),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_210 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(start),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(x_in[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(x_in[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(x_in[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(x_in[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(x_in[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(x_in[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(x_in[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(x_in[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(x_in[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(x_in[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(x_in[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(x_in[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(x_in[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(x_in[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(x_in[8]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(x_in[9]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(y_in[0]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(y_in[10]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(y_in[11]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(y_in[12]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(y_in[13]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(y_in[14]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(y_in[15]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(y_in[1]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(y_in[2]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(y_in[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(y_in[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(y_in[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(y_in[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(y_in[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(y_in[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(y_in[9]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(z_in[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(z_in[10]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(z_in[11]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(z_in[12]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(z_in[13]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(z_in[14]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(z_in[15]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(z_in[1]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(z_in[2]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(z_in[3]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(z_in[4]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(z_in[5]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(z_in[6]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(z_in[7]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(z_in[8]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(z_in[9]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net51),
    .X(done));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net52),
    .X(x_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net53),
    .X(x_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net54),
    .X(x_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net55),
    .X(x_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net56),
    .X(x_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net57),
    .X(x_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net58),
    .X(x_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net59),
    .X(x_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net60),
    .X(x_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net61),
    .X(x_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net62),
    .X(x_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net63),
    .X(x_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net64),
    .X(x_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net65),
    .X(x_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net66),
    .X(x_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net67),
    .X(x_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net68),
    .X(y_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net69),
    .X(y_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net70),
    .X(y_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net71),
    .X(y_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net72),
    .X(y_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net73),
    .X(y_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net74),
    .X(y_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net75),
    .X(y_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net76),
    .X(y_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net77),
    .X(y_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net78),
    .X(y_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net79),
    .X(y_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net80),
    .X(y_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net81),
    .X(y_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net82),
    .X(y_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net83),
    .X(y_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net84),
    .X(z_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net85),
    .X(z_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net86),
    .X(z_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net87),
    .X(z_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net88),
    .X(z_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net89),
    .X(z_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net90),
    .X(z_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net91),
    .X(z_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net92),
    .X(z_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net93),
    .X(z_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net94),
    .X(z_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net95),
    .X(z_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net96),
    .X(z_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net97),
    .X(z_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net98),
    .X(z_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net99),
    .X(z_out[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload5 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(_0303_),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net101),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(\iteration[1] ),
    .X(net103));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer4 (.A(\iteration[1] ),
    .X(net104));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_271 ();
endmodule
