module handshake_synchronizer (dst_clk,
    dst_ready,
    dst_rst_n,
    dst_valid,
    src_clk,
    src_ready,
    src_rst_n,
    src_valid,
    dst_data,
    src_data);
 input dst_clk;
 input dst_ready;
 input dst_rst_n;
 output dst_valid;
 input src_clk;
 output src_ready;
 input src_rst_n;
 input src_valid;
 output [31:0] dst_data;
 input [31:0] src_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire \ack_sync[0] ;
 wire \ack_sync[1] ;
 wire \data_reg[0] ;
 wire \data_reg[10] ;
 wire \data_reg[11] ;
 wire \data_reg[12] ;
 wire \data_reg[13] ;
 wire \data_reg[14] ;
 wire \data_reg[15] ;
 wire \data_reg[16] ;
 wire \data_reg[17] ;
 wire \data_reg[18] ;
 wire \data_reg[19] ;
 wire \data_reg[1] ;
 wire \data_reg[20] ;
 wire \data_reg[21] ;
 wire \data_reg[22] ;
 wire \data_reg[23] ;
 wire \data_reg[24] ;
 wire \data_reg[25] ;
 wire \data_reg[26] ;
 wire \data_reg[27] ;
 wire \data_reg[28] ;
 wire \data_reg[29] ;
 wire \data_reg[2] ;
 wire \data_reg[30] ;
 wire \data_reg[31] ;
 wire \data_reg[3] ;
 wire \data_reg[4] ;
 wire \data_reg[5] ;
 wire \data_reg[6] ;
 wire \data_reg[7] ;
 wire \data_reg[8] ;
 wire \data_reg[9] ;
 wire dst_ack;
 wire dst_req;
 wire \req_sync[0] ;
 wire src_req;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire clknet_0_src_clk;
 wire clknet_2_0__leaf_src_clk;
 wire clknet_2_1__leaf_src_clk;
 wire clknet_2_2__leaf_src_clk;
 wire clknet_2_3__leaf_src_clk;
 wire net72;

 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _079_ (.A1(src_req),
    .A2(\ack_sync[1] ),
    .ZN(net71));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _080_ (.A1(net37),
    .A2(net71),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _081_ (.I(_067_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _082_ (.I0(\data_reg[0] ),
    .I1(net5),
    .S(_068_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _083_ (.I0(\data_reg[10] ),
    .I1(net6),
    .S(_068_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _084_ (.I0(\data_reg[11] ),
    .I1(net7),
    .S(_068_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _085_ (.I0(\data_reg[12] ),
    .I1(net8),
    .S(_068_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _086_ (.I0(\data_reg[13] ),
    .I1(net9),
    .S(_068_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _087_ (.I0(\data_reg[14] ),
    .I1(net10),
    .S(_068_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _088_ (.I0(\data_reg[15] ),
    .I1(net11),
    .S(_068_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _089_ (.I0(\data_reg[16] ),
    .I1(net12),
    .S(_068_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _090_ (.I0(\data_reg[17] ),
    .I1(net13),
    .S(_068_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _091_ (.I0(\data_reg[18] ),
    .I1(net14),
    .S(_068_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _092_ (.I(_067_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _093_ (.I0(\data_reg[19] ),
    .I1(net15),
    .S(_069_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _094_ (.I0(\data_reg[1] ),
    .I1(net16),
    .S(_069_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _095_ (.I0(\data_reg[20] ),
    .I1(net17),
    .S(_069_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _096_ (.I0(\data_reg[21] ),
    .I1(net18),
    .S(_069_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _097_ (.I0(\data_reg[22] ),
    .I1(net19),
    .S(_069_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _098_ (.I0(\data_reg[23] ),
    .I1(net20),
    .S(_069_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _099_ (.I0(\data_reg[24] ),
    .I1(net21),
    .S(_069_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _100_ (.I0(\data_reg[25] ),
    .I1(net22),
    .S(_069_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _101_ (.I0(\data_reg[26] ),
    .I1(net23),
    .S(_069_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _102_ (.I0(\data_reg[27] ),
    .I1(net24),
    .S(_069_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _103_ (.I(_067_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _104_ (.I0(\data_reg[28] ),
    .I1(net25),
    .S(_070_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _105_ (.I0(\data_reg[29] ),
    .I1(net26),
    .S(_070_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _106_ (.I0(\data_reg[2] ),
    .I1(net27),
    .S(_070_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _107_ (.I0(\data_reg[30] ),
    .I1(net28),
    .S(_070_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _108_ (.I0(\data_reg[31] ),
    .I1(net29),
    .S(_070_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _109_ (.I0(\data_reg[3] ),
    .I1(net30),
    .S(_070_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _110_ (.I0(\data_reg[4] ),
    .I1(net31),
    .S(_070_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _111_ (.I0(\data_reg[5] ),
    .I1(net32),
    .S(_070_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _112_ (.I0(\data_reg[6] ),
    .I1(net33),
    .S(_070_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _113_ (.I0(\data_reg[7] ),
    .I1(net34),
    .S(_070_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _114_ (.I0(\data_reg[8] ),
    .I1(net35),
    .S(_067_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _115_ (.I0(\data_reg[9] ),
    .I1(net36),
    .S(_067_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _116_ (.A1(net3),
    .A2(net70),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _117_ (.I0(dst_ack),
    .I1(dst_req),
    .S(_071_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _118_ (.A1(dst_ack),
    .A2(dst_req),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _119_ (.A1(net70),
    .A2(_072_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _120_ (.I(_073_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _121_ (.I0(\data_reg[0] ),
    .I1(net38),
    .S(_074_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _122_ (.I0(\data_reg[10] ),
    .I1(net39),
    .S(_074_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _123_ (.I0(\data_reg[11] ),
    .I1(net40),
    .S(_074_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _124_ (.I0(\data_reg[12] ),
    .I1(net41),
    .S(_074_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _125_ (.I0(\data_reg[13] ),
    .I1(net42),
    .S(_074_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _126_ (.I0(\data_reg[14] ),
    .I1(net43),
    .S(_074_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _127_ (.I0(\data_reg[15] ),
    .I1(net44),
    .S(_074_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _128_ (.I0(\data_reg[16] ),
    .I1(net45),
    .S(_074_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _129_ (.I0(\data_reg[17] ),
    .I1(net46),
    .S(_074_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _130_ (.I0(\data_reg[18] ),
    .I1(net47),
    .S(_074_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _131_ (.I(_073_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _132_ (.I0(\data_reg[19] ),
    .I1(net48),
    .S(_075_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _133_ (.I0(\data_reg[1] ),
    .I1(net49),
    .S(_075_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _134_ (.I0(\data_reg[20] ),
    .I1(net50),
    .S(_075_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _135_ (.I0(\data_reg[21] ),
    .I1(net51),
    .S(_075_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _136_ (.I0(\data_reg[22] ),
    .I1(net52),
    .S(_075_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _137_ (.I0(\data_reg[23] ),
    .I1(net53),
    .S(_075_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _138_ (.I0(\data_reg[24] ),
    .I1(net54),
    .S(_075_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _139_ (.I0(\data_reg[25] ),
    .I1(net55),
    .S(_075_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _140_ (.I0(\data_reg[26] ),
    .I1(net56),
    .S(_075_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _141_ (.I0(\data_reg[27] ),
    .I1(net57),
    .S(_075_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _142_ (.I(_073_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _143_ (.I0(\data_reg[28] ),
    .I1(net58),
    .S(_076_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _144_ (.I0(\data_reg[29] ),
    .I1(net59),
    .S(_076_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _145_ (.I0(\data_reg[2] ),
    .I1(net60),
    .S(_076_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _146_ (.I0(\data_reg[30] ),
    .I1(net61),
    .S(_076_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _147_ (.I0(\data_reg[31] ),
    .I1(net62),
    .S(_076_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _148_ (.I0(\data_reg[3] ),
    .I1(net63),
    .S(_076_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _149_ (.I0(\data_reg[4] ),
    .I1(net64),
    .S(_076_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _150_ (.I0(\data_reg[5] ),
    .I1(net65),
    .S(_076_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _151_ (.I0(\data_reg[6] ),
    .I1(net66),
    .S(_076_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _152_ (.I0(\data_reg[7] ),
    .I1(net67),
    .S(_076_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _153_ (.I0(\data_reg[8] ),
    .I1(net68),
    .S(_073_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _154_ (.I0(\data_reg[9] ),
    .I1(net69),
    .S(_073_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _155_ (.I(net70),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _156_ (.A1(_077_),
    .A2(_072_),
    .B(_071_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _157_ (.I(\ack_sync[1] ),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _158_ (.I0(src_req),
    .I1(_078_),
    .S(net37),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ack_sync[0]$_DFF_PN0_  (.D(dst_ack),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\ack_sync[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ack_sync[1]$_DFF_PN0_  (.D(\ack_sync[0] ),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\ack_sync[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[10]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[11]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[12]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[13]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[14]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[15]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[16]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[17]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\data_reg[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[18]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[19]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[1]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[20]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[21]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[22]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[23]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[24]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[25]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[26]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[27]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\data_reg[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[28]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[29]$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[2]$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[30]$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[31]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[3]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[4]$_DFFE_PN0P_  (.D(_026_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[5]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[6]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[7]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\data_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[8]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[9]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\data_reg[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_ack$_DFFE_PN0P_  (.D(_032_),
    .RN(net4),
    .CLK(net2),
    .Q(dst_ack));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[0]$_DFFE_PN0P_  (.D(_033_),
    .RN(net4),
    .CLK(net2),
    .Q(net38));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[10]$_DFFE_PN0P_  (.D(_034_),
    .RN(net4),
    .CLK(net2),
    .Q(net39));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[11]$_DFFE_PN0P_  (.D(_035_),
    .RN(net4),
    .CLK(net2),
    .Q(net40));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[12]$_DFFE_PN0P_  (.D(_036_),
    .RN(net4),
    .CLK(net2),
    .Q(net41));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[13]$_DFFE_PN0P_  (.D(_037_),
    .RN(net4),
    .CLK(net2),
    .Q(net42));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[14]$_DFFE_PN0P_  (.D(_038_),
    .RN(net4),
    .CLK(net2),
    .Q(net43));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[15]$_DFFE_PN0P_  (.D(_039_),
    .RN(net4),
    .CLK(net2),
    .Q(net44));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[16]$_DFFE_PN0P_  (.D(_040_),
    .RN(net4),
    .CLK(net2),
    .Q(net45));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[17]$_DFFE_PN0P_  (.D(_041_),
    .RN(net4),
    .CLK(net2),
    .Q(net46));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[18]$_DFFE_PN0P_  (.D(_042_),
    .RN(net4),
    .CLK(net2),
    .Q(net47));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[19]$_DFFE_PN0P_  (.D(_043_),
    .RN(net4),
    .CLK(net2),
    .Q(net48));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[1]$_DFFE_PN0P_  (.D(_044_),
    .RN(net4),
    .CLK(net2),
    .Q(net49));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[20]$_DFFE_PN0P_  (.D(_045_),
    .RN(net4),
    .CLK(net2),
    .Q(net50));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[21]$_DFFE_PN0P_  (.D(_046_),
    .RN(net4),
    .CLK(net2),
    .Q(net51));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[22]$_DFFE_PN0P_  (.D(_047_),
    .RN(net4),
    .CLK(net2),
    .Q(net52));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[23]$_DFFE_PN0P_  (.D(_048_),
    .RN(net4),
    .CLK(net2),
    .Q(net53));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[24]$_DFFE_PN0P_  (.D(_049_),
    .RN(net4),
    .CLK(net2),
    .Q(net54));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[25]$_DFFE_PN0P_  (.D(_050_),
    .RN(net4),
    .CLK(net2),
    .Q(net55));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[26]$_DFFE_PN0P_  (.D(_051_),
    .RN(net4),
    .CLK(net2),
    .Q(net56));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[27]$_DFFE_PN0P_  (.D(_052_),
    .RN(net4),
    .CLK(net2),
    .Q(net57));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[28]$_DFFE_PN0P_  (.D(_053_),
    .RN(net4),
    .CLK(net2),
    .Q(net58));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[29]$_DFFE_PN0P_  (.D(_054_),
    .RN(net4),
    .CLK(net2),
    .Q(net59));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[2]$_DFFE_PN0P_  (.D(_055_),
    .RN(net4),
    .CLK(net2),
    .Q(net60));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[30]$_DFFE_PN0P_  (.D(_056_),
    .RN(net4),
    .CLK(net2),
    .Q(net61));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[31]$_DFFE_PN0P_  (.D(_057_),
    .RN(net4),
    .CLK(net2),
    .Q(net62));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[3]$_DFFE_PN0P_  (.D(_058_),
    .RN(net4),
    .CLK(net2),
    .Q(net63));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[4]$_DFFE_PN0P_  (.D(_059_),
    .RN(net4),
    .CLK(net2),
    .Q(net64));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[5]$_DFFE_PN0P_  (.D(_060_),
    .RN(net4),
    .CLK(net2),
    .Q(net65));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[6]$_DFFE_PN0P_  (.D(_061_),
    .RN(net4),
    .CLK(net2),
    .Q(net66));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[7]$_DFFE_PN0P_  (.D(_062_),
    .RN(net4),
    .CLK(net2),
    .Q(net67));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[8]$_DFFE_PN0P_  (.D(_063_),
    .RN(net4),
    .CLK(net2),
    .Q(net68));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data_reg[9]$_DFFE_PN0P_  (.D(_064_),
    .RN(net4),
    .CLK(net2),
    .Q(net69));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_valid_reg$_DFFE_PN0P_  (.D(_065_),
    .RN(net4),
    .CLK(net2),
    .Q(net70));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \req_sync[0]$_DFF_PN0_  (.D(src_req),
    .RN(net4),
    .CLK(net2),
    .Q(\req_sync[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \req_sync[1]$_DFF_PN0_  (.D(\req_sync[0] ),
    .RN(net4),
    .CLK(net2),
    .Q(dst_req));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_req$_DFFE_PN0P_  (.D(_066_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(src_req));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 hold1 (.I(net72),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_67 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_68 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_69 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_70 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_71 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_72 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_73 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_74 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_75 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_76 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_77 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input1 (.I(dst_clk),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(dst_ready),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 input3 (.I(dst_rst_n),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(src_data[0]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(src_data[10]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(src_data[11]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(src_data[12]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(src_data[13]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(src_data[14]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(src_data[15]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(src_data[16]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(src_data[17]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(src_data[18]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(src_data[19]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(src_data[1]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(src_data[20]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(src_data[21]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(src_data[22]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(src_data[23]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(src_data[24]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(src_data[25]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(src_data[26]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(src_data[27]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(src_data[28]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(src_data[29]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(src_data[2]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(src_data[30]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(src_data[31]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(src_data[3]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(src_data[4]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(src_data[5]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(src_data[6]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input33 (.I(src_data[7]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(src_data[8]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(src_data[9]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(src_valid),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output37 (.I(net38),
    .Z(dst_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output38 (.I(net39),
    .Z(dst_data[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net40),
    .Z(dst_data[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output40 (.I(net41),
    .Z(dst_data[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output41 (.I(net42),
    .Z(dst_data[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output42 (.I(net43),
    .Z(dst_data[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output43 (.I(net44),
    .Z(dst_data[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output44 (.I(net45),
    .Z(dst_data[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output45 (.I(net46),
    .Z(dst_data[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output46 (.I(net47),
    .Z(dst_data[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output47 (.I(net48),
    .Z(dst_data[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net49),
    .Z(dst_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net50),
    .Z(dst_data[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net51),
    .Z(dst_data[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output51 (.I(net52),
    .Z(dst_data[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output52 (.I(net53),
    .Z(dst_data[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output53 (.I(net54),
    .Z(dst_data[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output54 (.I(net55),
    .Z(dst_data[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output55 (.I(net56),
    .Z(dst_data[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output56 (.I(net57),
    .Z(dst_data[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output57 (.I(net58),
    .Z(dst_data[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output58 (.I(net59),
    .Z(dst_data[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output59 (.I(net60),
    .Z(dst_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output60 (.I(net61),
    .Z(dst_data[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output61 (.I(net62),
    .Z(dst_data[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net63),
    .Z(dst_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net64),
    .Z(dst_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net65),
    .Z(dst_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net66),
    .Z(dst_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net67),
    .Z(dst_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net68),
    .Z(dst_data[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net69),
    .Z(dst_data[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net70),
    .Z(dst_valid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net71),
    .Z(src_ready));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_src_clk (.I(src_clk),
    .Z(clknet_0_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_0__f_src_clk (.I(clknet_0_src_clk),
    .Z(clknet_2_0__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_1__f_src_clk (.I(clknet_0_src_clk),
    .Z(clknet_2_1__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_2__f_src_clk (.I(clknet_0_src_clk),
    .Z(clknet_2_2__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_3__f_src_clk (.I(clknet_0_src_clk),
    .Z(clknet_2_3__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload0 (.I(clknet_2_0__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload1 (.I(clknet_2_1__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload2 (.I(clknet_2_2__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(src_rst_n),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_285 ();
endmodule
