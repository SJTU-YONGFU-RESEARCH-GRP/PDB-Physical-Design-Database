module configurable_prng (clk,
    enable,
    reseed,
    rst_n,
    valid,
    random,
    seed_in);
 input clk;
 input enable;
 input reseed;
 input rst_n;
 output valid;
 output [15:0] random;
 input [15:0] seed_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 CLKBUF_X3 _093_ (.A(reseed),
    .Z(_038_));
 INV_X2 _094_ (.A(_038_),
    .ZN(_039_));
 BUF_X2 _095_ (.A(rst_n),
    .Z(_040_));
 NAND2_X1 _096_ (.A1(_039_),
    .A2(_040_),
    .ZN(_041_));
 INV_X1 _097_ (.A(net33),
    .ZN(_042_));
 CLKBUF_X3 _098_ (.A(enable),
    .Z(_043_));
 CLKBUF_X3 _099_ (.A(_043_),
    .Z(_044_));
 INV_X1 _100_ (.A(_044_),
    .ZN(_045_));
 AOI21_X1 _101_ (.A(_041_),
    .B1(_042_),
    .B2(_045_),
    .ZN(_016_));
 XOR2_X1 _102_ (.A(net23),
    .B(net18),
    .Z(_046_));
 XNOR2_X1 _103_ (.A(net21),
    .B(net20),
    .ZN(_047_));
 XNOR2_X1 _104_ (.A(_046_),
    .B(_047_),
    .ZN(_048_));
 NOR3_X1 _105_ (.A1(_045_),
    .A2(_041_),
    .A3(_048_),
    .ZN(_049_));
 NOR4_X1 _106_ (.A1(net16),
    .A2(net15),
    .A3(net3),
    .A4(net6),
    .ZN(_050_));
 NOR4_X1 _107_ (.A1(net2),
    .A2(net5),
    .A3(net4),
    .A4(net7),
    .ZN(_051_));
 NOR4_X1 _108_ (.A1(net8),
    .A2(net1),
    .A3(net10),
    .A4(net13),
    .ZN(_052_));
 NOR4_X1 _109_ (.A1(net9),
    .A2(net12),
    .A3(net11),
    .A4(net14),
    .ZN(_053_));
 AND4_X1 _110_ (.A1(_050_),
    .A2(_051_),
    .A3(_052_),
    .A4(_053_),
    .ZN(_054_));
 BUF_X4 _111_ (.A(_054_),
    .Z(_055_));
 NAND2_X1 _112_ (.A1(_038_),
    .A2(_040_),
    .ZN(_056_));
 OAI33_X1 _113_ (.A1(_044_),
    .A2(net17),
    .A3(_041_),
    .B1(_055_),
    .B2(_056_),
    .B3(net1),
    .ZN(_057_));
 NOR2_X1 _114_ (.A1(_049_),
    .A2(_057_),
    .ZN(_000_));
 CLKBUF_X3 _115_ (.A(_040_),
    .Z(_058_));
 MUX2_X1 _116_ (.A(net18),
    .B(net32),
    .S(_044_),
    .Z(_059_));
 NOR2_X1 _117_ (.A1(_038_),
    .A2(_059_),
    .ZN(_060_));
 CLKBUF_X3 _118_ (.A(_039_),
    .Z(_061_));
 NOR3_X1 _119_ (.A1(_061_),
    .A2(net2),
    .A3(_055_),
    .ZN(_062_));
 OAI21_X1 _120_ (.A(_058_),
    .B1(_060_),
    .B2(_062_),
    .ZN(_001_));
 MUX2_X1 _121_ (.A(net19),
    .B(net18),
    .S(_044_),
    .Z(_063_));
 NOR2_X1 _122_ (.A1(_038_),
    .A2(_063_),
    .ZN(_064_));
 NOR3_X1 _123_ (.A1(_061_),
    .A2(net3),
    .A3(_055_),
    .ZN(_065_));
 OAI21_X1 _124_ (.A(_058_),
    .B1(_064_),
    .B2(_065_),
    .ZN(_002_));
 MUX2_X1 _125_ (.A(net20),
    .B(net19),
    .S(_044_),
    .Z(_066_));
 MUX2_X1 _126_ (.A(net4),
    .B(_066_),
    .S(_061_),
    .Z(_067_));
 AND2_X1 _127_ (.A1(_058_),
    .A2(_067_),
    .ZN(_003_));
 MUX2_X1 _128_ (.A(net21),
    .B(net20),
    .S(_044_),
    .Z(_068_));
 NOR2_X1 _129_ (.A1(_038_),
    .A2(_068_),
    .ZN(_069_));
 NOR3_X1 _130_ (.A1(_061_),
    .A2(net5),
    .A3(_055_),
    .ZN(_070_));
 OAI21_X1 _131_ (.A(_058_),
    .B1(_069_),
    .B2(_070_),
    .ZN(_004_));
 MUX2_X1 _132_ (.A(net22),
    .B(net21),
    .S(_043_),
    .Z(_071_));
 MUX2_X1 _133_ (.A(net6),
    .B(_071_),
    .S(_061_),
    .Z(_072_));
 AND2_X1 _134_ (.A1(_058_),
    .A2(_072_),
    .ZN(_005_));
 MUX2_X1 _135_ (.A(net23),
    .B(net22),
    .S(_044_),
    .Z(_073_));
 NOR2_X1 _136_ (.A1(_038_),
    .A2(_073_),
    .ZN(_074_));
 NOR3_X1 _137_ (.A1(_061_),
    .A2(net7),
    .A3(_055_),
    .ZN(_075_));
 OAI21_X1 _138_ (.A(_058_),
    .B1(_074_),
    .B2(_075_),
    .ZN(_006_));
 MUX2_X1 _139_ (.A(net24),
    .B(net17),
    .S(_043_),
    .Z(_017_));
 MUX2_X1 _140_ (.A(net8),
    .B(_017_),
    .S(_061_),
    .Z(_018_));
 AND2_X1 _141_ (.A1(_058_),
    .A2(_018_),
    .ZN(_007_));
 MUX2_X1 _142_ (.A(net25),
    .B(net24),
    .S(_043_),
    .Z(_019_));
 MUX2_X1 _143_ (.A(net9),
    .B(_019_),
    .S(_039_),
    .Z(_020_));
 AND2_X1 _144_ (.A1(_040_),
    .A2(_020_),
    .ZN(_008_));
 MUX2_X1 _145_ (.A(net26),
    .B(net25),
    .S(_043_),
    .Z(_021_));
 MUX2_X1 _146_ (.A(net10),
    .B(_021_),
    .S(_039_),
    .Z(_022_));
 AND2_X1 _147_ (.A1(_040_),
    .A2(_022_),
    .ZN(_009_));
 MUX2_X1 _148_ (.A(net27),
    .B(net26),
    .S(_043_),
    .Z(_023_));
 MUX2_X1 _149_ (.A(net11),
    .B(_023_),
    .S(_039_),
    .Z(_024_));
 AND2_X1 _150_ (.A1(_040_),
    .A2(_024_),
    .ZN(_010_));
 MUX2_X1 _151_ (.A(net28),
    .B(net27),
    .S(_044_),
    .Z(_025_));
 NOR2_X1 _152_ (.A1(_038_),
    .A2(_025_),
    .ZN(_026_));
 NOR3_X1 _153_ (.A1(_061_),
    .A2(net12),
    .A3(_055_),
    .ZN(_027_));
 OAI21_X1 _154_ (.A(_058_),
    .B1(_026_),
    .B2(_027_),
    .ZN(_011_));
 MUX2_X1 _155_ (.A(net29),
    .B(net28),
    .S(_044_),
    .Z(_028_));
 NOR2_X1 _156_ (.A1(_038_),
    .A2(_028_),
    .ZN(_029_));
 NOR3_X1 _157_ (.A1(_061_),
    .A2(net13),
    .A3(_055_),
    .ZN(_030_));
 OAI21_X1 _158_ (.A(_058_),
    .B1(_029_),
    .B2(_030_),
    .ZN(_012_));
 MUX2_X1 _159_ (.A(net30),
    .B(net29),
    .S(_044_),
    .Z(_031_));
 NOR2_X1 _160_ (.A1(_038_),
    .A2(_031_),
    .ZN(_032_));
 NOR3_X1 _161_ (.A1(_061_),
    .A2(net14),
    .A3(_055_),
    .ZN(_033_));
 OAI21_X1 _162_ (.A(_058_),
    .B1(_032_),
    .B2(_033_),
    .ZN(_013_));
 MUX2_X1 _163_ (.A(net31),
    .B(net30),
    .S(_043_),
    .Z(_034_));
 MUX2_X1 _164_ (.A(net15),
    .B(_034_),
    .S(_039_),
    .Z(_035_));
 AND2_X1 _165_ (.A1(_040_),
    .A2(_035_),
    .ZN(_014_));
 MUX2_X1 _166_ (.A(net32),
    .B(net31),
    .S(_043_),
    .Z(_036_));
 MUX2_X1 _167_ (.A(net16),
    .B(_036_),
    .S(_039_),
    .Z(_037_));
 AND2_X1 _168_ (.A1(_040_),
    .A2(_037_),
    .ZN(_015_));
 DFF_X1 \lfsr_reg[0]$_SDFFE_PN1P_  (.D(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net17),
    .QN(_092_));
 DFF_X1 \lfsr_reg[10]$_SDFFE_PN1P_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net18),
    .QN(_091_));
 DFF_X1 \lfsr_reg[11]$_SDFFE_PN1P_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net19),
    .QN(_090_));
 DFF_X1 \lfsr_reg[12]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net20),
    .QN(_089_));
 DFF_X1 \lfsr_reg[13]$_SDFFE_PN1P_  (.D(_004_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net21),
    .QN(_088_));
 DFF_X1 \lfsr_reg[14]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net22),
    .QN(_087_));
 DFF_X1 \lfsr_reg[15]$_SDFFE_PN1P_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net23),
    .QN(_086_));
 DFF_X1 \lfsr_reg[1]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net24),
    .QN(_085_));
 DFF_X1 \lfsr_reg[2]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net25),
    .QN(_084_));
 DFF_X1 \lfsr_reg[3]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net26),
    .QN(_083_));
 DFF_X1 \lfsr_reg[4]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net27),
    .QN(_082_));
 DFF_X1 \lfsr_reg[5]$_SDFFE_PN1P_  (.D(_011_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net28),
    .QN(_081_));
 DFF_X1 \lfsr_reg[6]$_SDFFE_PN1P_  (.D(_012_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net29),
    .QN(_080_));
 DFF_X1 \lfsr_reg[7]$_SDFFE_PN1P_  (.D(_013_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net30),
    .QN(_079_));
 DFF_X1 \lfsr_reg[8]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net31),
    .QN(_078_));
 DFF_X1 \lfsr_reg[9]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net32),
    .QN(_077_));
 DFF_X1 \valid_reg$_SDFFE_PP0P_  (.D(_016_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net33),
    .QN(_076_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_57 ();
 BUF_X1 input1 (.A(seed_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(seed_in[10]),
    .Z(net2));
 BUF_X1 input3 (.A(seed_in[11]),
    .Z(net3));
 BUF_X1 input4 (.A(seed_in[12]),
    .Z(net4));
 BUF_X1 input5 (.A(seed_in[13]),
    .Z(net5));
 BUF_X1 input6 (.A(seed_in[14]),
    .Z(net6));
 BUF_X1 input7 (.A(seed_in[15]),
    .Z(net7));
 BUF_X1 input8 (.A(seed_in[1]),
    .Z(net8));
 BUF_X1 input9 (.A(seed_in[2]),
    .Z(net9));
 BUF_X1 input10 (.A(seed_in[3]),
    .Z(net10));
 BUF_X1 input11 (.A(seed_in[4]),
    .Z(net11));
 BUF_X1 input12 (.A(seed_in[5]),
    .Z(net12));
 BUF_X1 input13 (.A(seed_in[6]),
    .Z(net13));
 BUF_X1 input14 (.A(seed_in[7]),
    .Z(net14));
 BUF_X1 input15 (.A(seed_in[8]),
    .Z(net15));
 BUF_X1 input16 (.A(seed_in[9]),
    .Z(net16));
 BUF_X1 output17 (.A(net17),
    .Z(random[0]));
 BUF_X1 output18 (.A(net18),
    .Z(random[10]));
 BUF_X1 output19 (.A(net19),
    .Z(random[11]));
 BUF_X1 output20 (.A(net20),
    .Z(random[12]));
 BUF_X1 output21 (.A(net21),
    .Z(random[13]));
 BUF_X1 output22 (.A(net22),
    .Z(random[14]));
 BUF_X1 output23 (.A(net23),
    .Z(random[15]));
 BUF_X1 output24 (.A(net24),
    .Z(random[1]));
 BUF_X1 output25 (.A(net25),
    .Z(random[2]));
 BUF_X1 output26 (.A(net26),
    .Z(random[3]));
 BUF_X1 output27 (.A(net27),
    .Z(random[4]));
 BUF_X1 output28 (.A(net28),
    .Z(random[5]));
 BUF_X1 output29 (.A(net29),
    .Z(random[6]));
 BUF_X1 output30 (.A(net30),
    .Z(random[7]));
 BUF_X1 output31 (.A(net31),
    .Z(random[8]));
 BUF_X1 output32 (.A(net32),
    .Z(random[9]));
 BUF_X1 output33 (.A(net33),
    .Z(valid));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X8 FILLER_0_81 ();
 FILLCELL_X2 FILLER_0_89 ();
 FILLCELL_X4 FILLER_0_101 ();
 FILLCELL_X1 FILLER_0_105 ();
 FILLCELL_X2 FILLER_0_121 ();
 FILLCELL_X1 FILLER_0_123 ();
 FILLCELL_X2 FILLER_0_127 ();
 FILLCELL_X1 FILLER_0_129 ();
 FILLCELL_X4 FILLER_0_133 ();
 FILLCELL_X2 FILLER_0_137 ();
 FILLCELL_X1 FILLER_0_139 ();
 FILLCELL_X32 FILLER_0_145 ();
 FILLCELL_X32 FILLER_0_177 ();
 FILLCELL_X8 FILLER_0_209 ();
 FILLCELL_X2 FILLER_0_217 ();
 FILLCELL_X1 FILLER_0_219 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X16 FILLER_1_65 ();
 FILLCELL_X4 FILLER_1_81 ();
 FILLCELL_X2 FILLER_1_85 ();
 FILLCELL_X1 FILLER_1_87 ();
 FILLCELL_X4 FILLER_1_91 ();
 FILLCELL_X2 FILLER_1_95 ();
 FILLCELL_X16 FILLER_1_100 ();
 FILLCELL_X1 FILLER_1_116 ();
 FILLCELL_X32 FILLER_1_134 ();
 FILLCELL_X32 FILLER_1_166 ();
 FILLCELL_X16 FILLER_1_198 ();
 FILLCELL_X4 FILLER_1_214 ();
 FILLCELL_X2 FILLER_1_218 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X16 FILLER_2_65 ();
 FILLCELL_X8 FILLER_2_81 ();
 FILLCELL_X2 FILLER_2_117 ();
 FILLCELL_X2 FILLER_2_123 ();
 FILLCELL_X1 FILLER_2_125 ();
 FILLCELL_X32 FILLER_2_133 ();
 FILLCELL_X32 FILLER_2_165 ();
 FILLCELL_X16 FILLER_2_197 ();
 FILLCELL_X4 FILLER_2_213 ();
 FILLCELL_X2 FILLER_2_217 ();
 FILLCELL_X1 FILLER_2_219 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X8 FILLER_3_97 ();
 FILLCELL_X4 FILLER_3_105 ();
 FILLCELL_X2 FILLER_3_109 ();
 FILLCELL_X4 FILLER_3_118 ();
 FILLCELL_X2 FILLER_3_122 ();
 FILLCELL_X32 FILLER_3_131 ();
 FILLCELL_X32 FILLER_3_163 ();
 FILLCELL_X16 FILLER_3_195 ();
 FILLCELL_X8 FILLER_3_211 ();
 FILLCELL_X1 FILLER_3_219 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X8 FILLER_4_97 ();
 FILLCELL_X4 FILLER_4_105 ();
 FILLCELL_X2 FILLER_4_109 ();
 FILLCELL_X1 FILLER_4_111 ();
 FILLCELL_X32 FILLER_4_117 ();
 FILLCELL_X32 FILLER_4_149 ();
 FILLCELL_X32 FILLER_4_181 ();
 FILLCELL_X4 FILLER_4_213 ();
 FILLCELL_X2 FILLER_4_217 ();
 FILLCELL_X1 FILLER_4_219 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X16 FILLER_5_65 ();
 FILLCELL_X8 FILLER_5_81 ();
 FILLCELL_X1 FILLER_5_89 ();
 FILLCELL_X8 FILLER_5_104 ();
 FILLCELL_X4 FILLER_5_112 ();
 FILLCELL_X2 FILLER_5_116 ();
 FILLCELL_X1 FILLER_5_118 ();
 FILLCELL_X32 FILLER_5_136 ();
 FILLCELL_X32 FILLER_5_168 ();
 FILLCELL_X16 FILLER_5_200 ();
 FILLCELL_X4 FILLER_5_216 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_65 ();
 FILLCELL_X4 FILLER_6_73 ();
 FILLCELL_X1 FILLER_6_77 ();
 FILLCELL_X4 FILLER_6_95 ();
 FILLCELL_X16 FILLER_6_103 ();
 FILLCELL_X4 FILLER_6_130 ();
 FILLCELL_X2 FILLER_6_134 ();
 FILLCELL_X32 FILLER_6_143 ();
 FILLCELL_X32 FILLER_6_175 ();
 FILLCELL_X8 FILLER_6_207 ();
 FILLCELL_X4 FILLER_6_215 ();
 FILLCELL_X1 FILLER_6_219 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X16 FILLER_7_193 ();
 FILLCELL_X8 FILLER_7_209 ();
 FILLCELL_X2 FILLER_7_217 ();
 FILLCELL_X1 FILLER_7_219 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X16 FILLER_8_65 ();
 FILLCELL_X8 FILLER_8_81 ();
 FILLCELL_X2 FILLER_8_89 ();
 FILLCELL_X1 FILLER_8_91 ();
 FILLCELL_X32 FILLER_8_106 ();
 FILLCELL_X32 FILLER_8_138 ();
 FILLCELL_X32 FILLER_8_170 ();
 FILLCELL_X16 FILLER_8_202 ();
 FILLCELL_X2 FILLER_8_218 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X4 FILLER_9_81 ();
 FILLCELL_X2 FILLER_9_85 ();
 FILLCELL_X1 FILLER_9_87 ();
 FILLCELL_X4 FILLER_9_109 ();
 FILLCELL_X8 FILLER_9_121 ();
 FILLCELL_X4 FILLER_9_129 ();
 FILLCELL_X2 FILLER_9_133 ();
 FILLCELL_X1 FILLER_9_135 ();
 FILLCELL_X1 FILLER_9_143 ();
 FILLCELL_X16 FILLER_9_161 ();
 FILLCELL_X4 FILLER_9_177 ();
 FILLCELL_X32 FILLER_9_184 ();
 FILLCELL_X4 FILLER_9_216 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X8 FILLER_10_65 ();
 FILLCELL_X4 FILLER_10_73 ();
 FILLCELL_X2 FILLER_10_77 ();
 FILLCELL_X4 FILLER_10_100 ();
 FILLCELL_X2 FILLER_10_104 ();
 FILLCELL_X2 FILLER_10_110 ();
 FILLCELL_X8 FILLER_10_116 ();
 FILLCELL_X2 FILLER_10_124 ();
 FILLCELL_X4 FILLER_10_131 ();
 FILLCELL_X1 FILLER_10_135 ();
 FILLCELL_X1 FILLER_10_143 ();
 FILLCELL_X32 FILLER_10_148 ();
 FILLCELL_X32 FILLER_10_180 ();
 FILLCELL_X8 FILLER_10_212 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X2 FILLER_11_97 ();
 FILLCELL_X1 FILLER_11_99 ();
 FILLCELL_X2 FILLER_11_104 ();
 FILLCELL_X4 FILLER_11_109 ();
 FILLCELL_X1 FILLER_11_113 ();
 FILLCELL_X4 FILLER_11_119 ();
 FILLCELL_X2 FILLER_11_123 ();
 FILLCELL_X32 FILLER_11_131 ();
 FILLCELL_X16 FILLER_11_163 ();
 FILLCELL_X4 FILLER_11_179 ();
 FILLCELL_X32 FILLER_11_186 ();
 FILLCELL_X2 FILLER_11_218 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_37 ();
 FILLCELL_X4 FILLER_12_69 ();
 FILLCELL_X2 FILLER_12_90 ();
 FILLCELL_X1 FILLER_12_92 ();
 FILLCELL_X16 FILLER_12_103 ();
 FILLCELL_X8 FILLER_12_119 ();
 FILLCELL_X4 FILLER_12_127 ();
 FILLCELL_X1 FILLER_12_131 ();
 FILLCELL_X4 FILLER_12_139 ();
 FILLCELL_X2 FILLER_12_143 ();
 FILLCELL_X1 FILLER_12_145 ();
 FILLCELL_X4 FILLER_12_149 ();
 FILLCELL_X1 FILLER_12_153 ();
 FILLCELL_X4 FILLER_12_171 ();
 FILLCELL_X2 FILLER_12_175 ();
 FILLCELL_X1 FILLER_12_177 ();
 FILLCELL_X32 FILLER_12_181 ();
 FILLCELL_X4 FILLER_12_213 ();
 FILLCELL_X2 FILLER_12_217 ();
 FILLCELL_X1 FILLER_12_219 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X16 FILLER_13_65 ();
 FILLCELL_X4 FILLER_13_81 ();
 FILLCELL_X2 FILLER_13_85 ();
 FILLCELL_X16 FILLER_13_97 ();
 FILLCELL_X4 FILLER_13_113 ();
 FILLCELL_X2 FILLER_13_117 ();
 FILLCELL_X8 FILLER_13_133 ();
 FILLCELL_X2 FILLER_13_141 ();
 FILLCELL_X2 FILLER_13_149 ();
 FILLCELL_X32 FILLER_13_155 ();
 FILLCELL_X4 FILLER_13_187 ();
 FILLCELL_X2 FILLER_13_191 ();
 FILLCELL_X16 FILLER_13_199 ();
 FILLCELL_X4 FILLER_13_215 ();
 FILLCELL_X1 FILLER_13_219 ();
 FILLCELL_X16 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_17 ();
 FILLCELL_X32 FILLER_14_21 ();
 FILLCELL_X32 FILLER_14_53 ();
 FILLCELL_X2 FILLER_14_85 ();
 FILLCELL_X4 FILLER_14_106 ();
 FILLCELL_X2 FILLER_14_110 ();
 FILLCELL_X1 FILLER_14_112 ();
 FILLCELL_X1 FILLER_14_119 ();
 FILLCELL_X16 FILLER_14_127 ();
 FILLCELL_X8 FILLER_14_143 ();
 FILLCELL_X1 FILLER_14_151 ();
 FILLCELL_X2 FILLER_14_154 ();
 FILLCELL_X8 FILLER_14_173 ();
 FILLCELL_X2 FILLER_14_181 ();
 FILLCELL_X32 FILLER_14_186 ();
 FILLCELL_X2 FILLER_14_218 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X4 FILLER_15_17 ();
 FILLCELL_X2 FILLER_15_21 ();
 FILLCELL_X32 FILLER_15_26 ();
 FILLCELL_X16 FILLER_15_58 ();
 FILLCELL_X8 FILLER_15_74 ();
 FILLCELL_X4 FILLER_15_82 ();
 FILLCELL_X2 FILLER_15_86 ();
 FILLCELL_X32 FILLER_15_105 ();
 FILLCELL_X32 FILLER_15_137 ();
 FILLCELL_X32 FILLER_15_169 ();
 FILLCELL_X16 FILLER_15_201 ();
 FILLCELL_X2 FILLER_15_217 ();
 FILLCELL_X1 FILLER_15_219 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X16 FILLER_16_65 ();
 FILLCELL_X2 FILLER_16_81 ();
 FILLCELL_X1 FILLER_16_83 ();
 FILLCELL_X16 FILLER_16_89 ();
 FILLCELL_X2 FILLER_16_105 ();
 FILLCELL_X16 FILLER_16_112 ();
 FILLCELL_X4 FILLER_16_128 ();
 FILLCELL_X2 FILLER_16_132 ();
 FILLCELL_X1 FILLER_16_134 ();
 FILLCELL_X32 FILLER_16_149 ();
 FILLCELL_X4 FILLER_16_181 ();
 FILLCELL_X1 FILLER_16_185 ();
 FILLCELL_X16 FILLER_16_192 ();
 FILLCELL_X8 FILLER_16_208 ();
 FILLCELL_X4 FILLER_16_216 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_9 ();
 FILLCELL_X2 FILLER_17_13 ();
 FILLCELL_X1 FILLER_17_15 ();
 FILLCELL_X32 FILLER_17_19 ();
 FILLCELL_X32 FILLER_17_51 ();
 FILLCELL_X16 FILLER_17_83 ();
 FILLCELL_X8 FILLER_17_99 ();
 FILLCELL_X4 FILLER_17_107 ();
 FILLCELL_X16 FILLER_17_115 ();
 FILLCELL_X1 FILLER_17_131 ();
 FILLCELL_X8 FILLER_17_137 ();
 FILLCELL_X1 FILLER_17_145 ();
 FILLCELL_X4 FILLER_17_150 ();
 FILLCELL_X1 FILLER_17_154 ();
 FILLCELL_X8 FILLER_17_172 ();
 FILLCELL_X32 FILLER_17_183 ();
 FILLCELL_X4 FILLER_17_215 ();
 FILLCELL_X1 FILLER_17_219 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X16 FILLER_18_97 ();
 FILLCELL_X8 FILLER_18_120 ();
 FILLCELL_X4 FILLER_18_128 ();
 FILLCELL_X2 FILLER_18_132 ();
 FILLCELL_X2 FILLER_18_140 ();
 FILLCELL_X32 FILLER_18_148 ();
 FILLCELL_X32 FILLER_18_180 ();
 FILLCELL_X8 FILLER_18_212 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X16 FILLER_19_65 ();
 FILLCELL_X8 FILLER_19_81 ();
 FILLCELL_X4 FILLER_19_89 ();
 FILLCELL_X2 FILLER_19_93 ();
 FILLCELL_X1 FILLER_19_95 ();
 FILLCELL_X2 FILLER_19_103 ();
 FILLCELL_X1 FILLER_19_105 ();
 FILLCELL_X2 FILLER_19_130 ();
 FILLCELL_X32 FILLER_19_145 ();
 FILLCELL_X32 FILLER_19_177 ();
 FILLCELL_X8 FILLER_19_209 ();
 FILLCELL_X2 FILLER_19_217 ();
 FILLCELL_X1 FILLER_19_219 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X16 FILLER_20_100 ();
 FILLCELL_X2 FILLER_20_116 ();
 FILLCELL_X4 FILLER_20_121 ();
 FILLCELL_X4 FILLER_20_132 ();
 FILLCELL_X4 FILLER_20_146 ();
 FILLCELL_X1 FILLER_20_150 ();
 FILLCELL_X32 FILLER_20_168 ();
 FILLCELL_X16 FILLER_20_200 ();
 FILLCELL_X4 FILLER_20_216 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X16 FILLER_21_65 ();
 FILLCELL_X8 FILLER_21_81 ();
 FILLCELL_X4 FILLER_21_89 ();
 FILLCELL_X2 FILLER_21_93 ();
 FILLCELL_X1 FILLER_21_95 ();
 FILLCELL_X8 FILLER_21_100 ();
 FILLCELL_X16 FILLER_21_112 ();
 FILLCELL_X8 FILLER_21_128 ();
 FILLCELL_X4 FILLER_21_136 ();
 FILLCELL_X2 FILLER_21_140 ();
 FILLCELL_X1 FILLER_21_142 ();
 FILLCELL_X32 FILLER_21_147 ();
 FILLCELL_X32 FILLER_21_179 ();
 FILLCELL_X8 FILLER_21_211 ();
 FILLCELL_X1 FILLER_21_219 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X16 FILLER_22_65 ();
 FILLCELL_X8 FILLER_22_81 ();
 FILLCELL_X2 FILLER_22_89 ();
 FILLCELL_X2 FILLER_22_121 ();
 FILLCELL_X32 FILLER_22_138 ();
 FILLCELL_X32 FILLER_22_170 ();
 FILLCELL_X16 FILLER_22_202 ();
 FILLCELL_X2 FILLER_22_218 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X4 FILLER_23_129 ();
 FILLCELL_X2 FILLER_23_133 ();
 FILLCELL_X32 FILLER_23_152 ();
 FILLCELL_X32 FILLER_23_184 ();
 FILLCELL_X4 FILLER_23_216 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X16 FILLER_24_97 ();
 FILLCELL_X1 FILLER_24_113 ();
 FILLCELL_X32 FILLER_24_131 ();
 FILLCELL_X32 FILLER_24_163 ();
 FILLCELL_X16 FILLER_24_195 ();
 FILLCELL_X8 FILLER_24_211 ();
 FILLCELL_X1 FILLER_24_219 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X16 FILLER_25_193 ();
 FILLCELL_X8 FILLER_25_209 ();
 FILLCELL_X2 FILLER_25_217 ();
 FILLCELL_X1 FILLER_25_219 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X16 FILLER_26_193 ();
 FILLCELL_X8 FILLER_26_209 ();
 FILLCELL_X2 FILLER_26_217 ();
 FILLCELL_X1 FILLER_26_219 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X8 FILLER_27_97 ();
 FILLCELL_X4 FILLER_27_105 ();
 FILLCELL_X2 FILLER_27_109 ();
 FILLCELL_X1 FILLER_27_111 ();
 FILLCELL_X16 FILLER_27_115 ();
 FILLCELL_X4 FILLER_27_131 ();
 FILLCELL_X1 FILLER_27_135 ();
 FILLCELL_X32 FILLER_27_139 ();
 FILLCELL_X32 FILLER_27_171 ();
 FILLCELL_X16 FILLER_27_203 ();
 FILLCELL_X1 FILLER_27_219 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X2 FILLER_28_97 ();
 FILLCELL_X1 FILLER_28_99 ();
 FILLCELL_X1 FILLER_28_103 ();
 FILLCELL_X2 FILLER_28_107 ();
 FILLCELL_X4 FILLER_28_115 ();
 FILLCELL_X2 FILLER_28_119 ();
 FILLCELL_X8 FILLER_28_124 ();
 FILLCELL_X2 FILLER_28_132 ();
 FILLCELL_X8 FILLER_28_137 ();
 FILLCELL_X4 FILLER_28_145 ();
 FILLCELL_X2 FILLER_28_149 ();
 FILLCELL_X32 FILLER_28_154 ();
 FILLCELL_X32 FILLER_28_186 ();
 FILLCELL_X2 FILLER_28_218 ();
endmodule
