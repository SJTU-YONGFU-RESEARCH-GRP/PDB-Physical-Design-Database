module configurable_mult (sign_mode,
    a,
    b,
    product);
 input sign_mode;
 input [7:0] a;
 input [7:0] b;
 output [15:0] product;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire _486_;
 wire _487_;
 wire _488_;
 wire _489_;
 wire _490_;
 wire _491_;
 wire _492_;
 wire _493_;
 wire _494_;
 wire _495_;
 wire _496_;
 wire _497_;
 wire _498_;
 wire _499_;
 wire _500_;
 wire _501_;
 wire _502_;
 wire _503_;
 wire _504_;
 wire _505_;
 wire _506_;
 wire _507_;
 wire _508_;
 wire _509_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;

 sky130_fd_sc_hd__buf_2 _510_ (.A(net5),
    .X(_000_));
 sky130_fd_sc_hd__buf_2 _511_ (.A(a[1]),
    .X(_001_));
 sky130_fd_sc_hd__and2_0 _512_ (.A(_000_),
    .B(_001_),
    .X(_387_));
 sky130_fd_sc_hd__buf_2 _513_ (.A(b[1]),
    .X(_002_));
 sky130_fd_sc_hd__and2_0 _514_ (.A(net1),
    .B(_002_),
    .X(_386_));
 sky130_fd_sc_hd__nand2_1 _515_ (.A(net1),
    .B(net6),
    .Y(_111_));
 sky130_fd_sc_hd__buf_2 _516_ (.A(a[3]),
    .X(_003_));
 sky130_fd_sc_hd__nand2_1 _517_ (.A(_000_),
    .B(_003_),
    .Y(_116_));
 sky130_fd_sc_hd__buf_2 _518_ (.A(a[2]),
    .X(_004_));
 sky130_fd_sc_hd__nand2_1 _519_ (.A(_002_),
    .B(_004_),
    .Y(_117_));
 sky130_fd_sc_hd__nand2_1 _520_ (.A(_001_),
    .B(net6),
    .Y(_118_));
 sky130_fd_sc_hd__nand2_1 _521_ (.A(net1),
    .B(net7),
    .Y(_121_));
 sky130_fd_sc_hd__clkbuf_4 _522_ (.A(a[4]),
    .X(_005_));
 sky130_fd_sc_hd__nand2_1 _523_ (.A(_000_),
    .B(_005_),
    .Y(_125_));
 sky130_fd_sc_hd__nand2_1 _524_ (.A(_002_),
    .B(_003_),
    .Y(_124_));
 sky130_fd_sc_hd__nand2_1 _525_ (.A(_004_),
    .B(net6),
    .Y(_126_));
 sky130_fd_sc_hd__and2_0 _526_ (.A(_001_),
    .B(net7),
    .X(_396_));
 sky130_fd_sc_hd__and2_0 _527_ (.A(net1),
    .B(net8),
    .X(_397_));
 sky130_fd_sc_hd__nand2_1 _528_ (.A(_000_),
    .B(net2),
    .Y(_134_));
 sky130_fd_sc_hd__nand2_1 _529_ (.A(_002_),
    .B(_005_),
    .Y(_132_));
 sky130_fd_sc_hd__nand2_1 _530_ (.A(net6),
    .B(_003_),
    .Y(_133_));
 sky130_fd_sc_hd__nand2_1 _531_ (.A(net1),
    .B(net9),
    .Y(_139_));
 sky130_fd_sc_hd__nand2_1 _532_ (.A(_000_),
    .B(net3),
    .Y(_151_));
 sky130_fd_sc_hd__nand2_1 _533_ (.A(_002_),
    .B(net2),
    .Y(_150_));
 sky130_fd_sc_hd__nand2_1 _534_ (.A(net6),
    .B(_005_),
    .Y(_149_));
 sky130_fd_sc_hd__nand2_1 _535_ (.A(_001_),
    .B(net9),
    .Y(_154_));
 sky130_fd_sc_hd__and2_0 _536_ (.A(net1),
    .B(net10),
    .X(_408_));
 sky130_fd_sc_hd__nand2_1 _537_ (.A(_002_),
    .B(net3),
    .Y(_173_));
 sky130_fd_sc_hd__inv_1 _538_ (.A(_173_),
    .Y(_414_));
 sky130_fd_sc_hd__nand2_1 _539_ (.A(net6),
    .B(net2),
    .Y(_174_));
 sky130_fd_sc_hd__nand2_1 _540_ (.A(_004_),
    .B(net9),
    .Y(_177_));
 sky130_fd_sc_hd__buf_2 _541_ (.A(net4),
    .X(_006_));
 sky130_fd_sc_hd__and2_0 _542_ (.A(_002_),
    .B(_006_),
    .X(_425_));
 sky130_fd_sc_hd__and2_0 _543_ (.A(net6),
    .B(net3),
    .X(_426_));
 sky130_fd_sc_hd__and2_0 _544_ (.A(net7),
    .B(net2),
    .X(_209_));
 sky130_fd_sc_hd__and2_0 _545_ (.A(_005_),
    .B(net8),
    .X(_210_));
 sky130_fd_sc_hd__and2_0 _546_ (.A(_003_),
    .B(net9),
    .X(_211_));
 sky130_fd_sc_hd__nand2_1 _547_ (.A(_004_),
    .B(net10),
    .Y(_219_));
 sky130_fd_sc_hd__inv_1 _548_ (.A(_219_),
    .Y(_429_));
 sky130_fd_sc_hd__clkbuf_4 _549_ (.A(net11),
    .X(_007_));
 sky130_fd_sc_hd__nor2b_1 _550_ (.A(_001_),
    .B_N(_007_),
    .Y(_432_));
 sky130_fd_sc_hd__inv_1 _551_ (.A(_239_),
    .Y(_236_));
 sky130_fd_sc_hd__nand2_1 _552_ (.A(net6),
    .B(_006_),
    .Y(_246_));
 sky130_fd_sc_hd__inv_1 _553_ (.A(_246_),
    .Y(_434_));
 sky130_fd_sc_hd__and2_0 _554_ (.A(net7),
    .B(net3),
    .X(_240_));
 sky130_fd_sc_hd__and2_0 _555_ (.A(net8),
    .B(net2),
    .X(_241_));
 sky130_fd_sc_hd__and2_0 _556_ (.A(_005_),
    .B(net9),
    .X(_242_));
 sky130_fd_sc_hd__nand2_1 _557_ (.A(_003_),
    .B(net10),
    .Y(_250_));
 sky130_fd_sc_hd__inv_1 _558_ (.A(_250_),
    .Y(_435_));
 sky130_fd_sc_hd__nor2b_1 _559_ (.A(_004_),
    .B_N(net11),
    .Y(_440_));
 sky130_fd_sc_hd__nand2_1 _560_ (.A(net7),
    .B(_006_),
    .Y(_276_));
 sky130_fd_sc_hd__inv_1 _561_ (.A(_276_),
    .Y(_315_));
 sky130_fd_sc_hd__nand2_1 _562_ (.A(_005_),
    .B(net10),
    .Y(_281_));
 sky130_fd_sc_hd__inv_1 _563_ (.A(_281_),
    .Y(_444_));
 sky130_fd_sc_hd__inv_1 _564_ (.A(_171_),
    .Y(_166_));
 sky130_fd_sc_hd__nand3_1 _565_ (.A(net5),
    .B(_002_),
    .C(net4),
    .Y(_008_));
 sky130_fd_sc_hd__nand2b_1 _566_ (.A_N(_439_),
    .B(_008_),
    .Y(_292_));
 sky130_fd_sc_hd__inv_1 _567_ (.A(_292_),
    .Y(_320_));
 sky130_fd_sc_hd__nor2b_1 _568_ (.A(_003_),
    .B_N(net11),
    .Y(_453_));
 sky130_fd_sc_hd__and2_1 _569_ (.A(net8),
    .B(_006_),
    .X(_316_));
 sky130_fd_sc_hd__and2_0 _570_ (.A(net9),
    .B(net3),
    .X(_317_));
 sky130_fd_sc_hd__nand2_1 _571_ (.A(net2),
    .B(net10),
    .Y(_308_));
 sky130_fd_sc_hd__inv_1 _572_ (.A(_308_),
    .Y(_463_));
 sky130_fd_sc_hd__nor2b_1 _573_ (.A(_005_),
    .B_N(net11),
    .Y(_470_));
 sky130_fd_sc_hd__and2_1 _574_ (.A(net9),
    .B(_006_),
    .X(_346_));
 sky130_fd_sc_hd__and2_0 _575_ (.A(net3),
    .B(net10),
    .X(_337_));
 sky130_fd_sc_hd__and2_0 _576_ (.A(net2),
    .B(_007_),
    .X(_338_));
 sky130_fd_sc_hd__nor2b_1 _577_ (.A(net2),
    .B_N(net11),
    .Y(_479_));
 sky130_fd_sc_hd__and2_1 _578_ (.A(net10),
    .B(_006_),
    .X(_485_));
 sky130_fd_sc_hd__and2_0 _579_ (.A(net3),
    .B(_007_),
    .X(_484_));
 sky130_fd_sc_hd__nor2b_1 _580_ (.A(net3),
    .B_N(net11),
    .Y(_492_));
 sky130_fd_sc_hd__and2_0 _581_ (.A(_006_),
    .B(_007_),
    .X(_497_));
 sky130_fd_sc_hd__nand2_1 _582_ (.A(_004_),
    .B(net7),
    .Y(_137_));
 sky130_fd_sc_hd__nand2_1 _583_ (.A(_000_),
    .B(net4),
    .Y(_172_));
 sky130_fd_sc_hd__nand2_1 _584_ (.A(net1),
    .B(_007_),
    .Y(_184_));
 sky130_fd_sc_hd__nand2_1 _585_ (.A(_003_),
    .B(net8),
    .Y(_178_));
 sky130_fd_sc_hd__nand2_1 _586_ (.A(_001_),
    .B(_007_),
    .Y(_218_));
 sky130_fd_sc_hd__inv_1 _587_ (.A(_427_),
    .Y(_245_));
 sky130_fd_sc_hd__nand2_1 _588_ (.A(net2),
    .B(net9),
    .Y(_275_));
 sky130_fd_sc_hd__nand2_1 _589_ (.A(_005_),
    .B(_007_),
    .Y(_307_));
 sky130_fd_sc_hd__nand2_1 _590_ (.A(_001_),
    .B(_002_),
    .Y(_112_));
 sky130_fd_sc_hd__nand2_1 _591_ (.A(_001_),
    .B(net8),
    .Y(_138_));
 sky130_fd_sc_hd__nand2_1 _592_ (.A(_004_),
    .B(net8),
    .Y(_155_));
 sky130_fd_sc_hd__inv_1 _593_ (.A(_170_),
    .Y(_165_));
 sky130_fd_sc_hd__nand2_1 _594_ (.A(net7),
    .B(_005_),
    .Y(_179_));
 sky130_fd_sc_hd__nand2b_1 _595_ (.A_N(net1),
    .B(net11),
    .Y(_200_));
 sky130_fd_sc_hd__nand2_1 _596_ (.A(_000_),
    .B(_004_),
    .Y(_113_));
 sky130_fd_sc_hd__nand2_1 _597_ (.A(_003_),
    .B(net7),
    .Y(_156_));
 sky130_fd_sc_hd__nand2_1 _598_ (.A(_001_),
    .B(net10),
    .Y(_185_));
 sky130_fd_sc_hd__nand2_1 _599_ (.A(_004_),
    .B(_007_),
    .Y(_252_));
 sky130_fd_sc_hd__nand2_1 _600_ (.A(net8),
    .B(net3),
    .Y(_277_));
 sky130_fd_sc_hd__nand2_1 _601_ (.A(_003_),
    .B(_007_),
    .Y(_282_));
 sky130_fd_sc_hd__inv_1 _602_ (.A(_213_),
    .Y(_215_));
 sky130_fd_sc_hd__inv_1 _603_ (.A(_229_),
    .Y(_233_));
 sky130_fd_sc_hd__inv_1 _604_ (.A(_244_),
    .Y(_247_));
 sky130_fd_sc_hd__inv_1 _605_ (.A(_262_),
    .Y(_268_));
 sky130_fd_sc_hd__inv_1 _606_ (.A(_267_),
    .Y(_270_));
 sky130_fd_sc_hd__inv_1 _607_ (.A(_288_),
    .Y(_289_));
 sky130_fd_sc_hd__inv_1 _608_ (.A(_294_),
    .Y(_300_));
 sky130_fd_sc_hd__inv_1 _609_ (.A(_298_),
    .Y(_301_));
 sky130_fd_sc_hd__inv_1 _610_ (.A(_319_),
    .Y(_321_));
 sky130_fd_sc_hd__inv_1 _611_ (.A(_328_),
    .Y(_330_));
 sky130_fd_sc_hd__inv_1 _612_ (.A(_348_),
    .Y(_349_));
 sky130_fd_sc_hd__inv_1 _613_ (.A(_355_),
    .Y(_356_));
 sky130_fd_sc_hd__inv_1 _614_ (.A(_369_),
    .Y(_370_));
 sky130_fd_sc_hd__inv_1 _615_ (.A(_379_),
    .Y(_380_));
 sky130_fd_sc_hd__inv_1 _616_ (.A(_212_),
    .Y(_251_));
 sky130_fd_sc_hd__inv_1 _617_ (.A(_228_),
    .Y(_269_));
 sky130_fd_sc_hd__inv_1 _618_ (.A(_243_),
    .Y(_280_));
 sky130_fd_sc_hd__inv_1 _619_ (.A(_261_),
    .Y(_299_));
 sky130_fd_sc_hd__inv_1 _620_ (.A(_266_),
    .Y(_304_));
 sky130_fd_sc_hd__inv_1 _621_ (.A(_287_),
    .Y(_311_));
 sky130_fd_sc_hd__inv_1 _622_ (.A(_293_),
    .Y(_329_));
 sky130_fd_sc_hd__inv_1 _623_ (.A(_297_),
    .Y(_333_));
 sky130_fd_sc_hd__inv_1 _624_ (.A(_327_),
    .Y(_359_));
 sky130_fd_sc_hd__inv_1 _625_ (.A(_354_),
    .Y(_373_));
 sky130_fd_sc_hd__inv_1 _626_ (.A(_368_),
    .Y(_383_));
 sky130_fd_sc_hd__inv_1 _627_ (.A(_123_),
    .Y(_393_));
 sky130_fd_sc_hd__inv_1 _628_ (.A(_122_),
    .Y(_399_));
 sky130_fd_sc_hd__inv_1 _629_ (.A(_130_),
    .Y(_145_));
 sky130_fd_sc_hd__inv_1 _630_ (.A(_140_),
    .Y(_407_));
 sky130_fd_sc_hd__inv_1 _631_ (.A(_202_),
    .Y(_421_));
 sky130_fd_sc_hd__inv_1 _632_ (.A(_162_),
    .Y(_190_));
 sky130_fd_sc_hd__xor2_1 _633_ (.A(_000_),
    .B(_002_),
    .X(_009_));
 sky130_fd_sc_hd__and2_0 _634_ (.A(_006_),
    .B(_009_),
    .X(_430_));
 sky130_fd_sc_hd__inv_1 _635_ (.A(_291_),
    .Y(_445_));
 sky130_fd_sc_hd__inv_1 _636_ (.A(_224_),
    .Y(_449_));
 sky130_fd_sc_hd__inv_1 _637_ (.A(_273_),
    .Y(_454_));
 sky130_fd_sc_hd__inv_1 _638_ (.A(_237_),
    .Y(_458_));
 sky130_fd_sc_hd__inv_1 _639_ (.A(_314_),
    .Y(_466_));
 sky130_fd_sc_hd__inv_1 _640_ (.A(_278_),
    .Y(_324_));
 sky130_fd_sc_hd__inv_1 _641_ (.A(_305_),
    .Y(_471_));
 sky130_fd_sc_hd__inv_1 _642_ (.A(_309_),
    .Y(_341_));
 sky130_fd_sc_hd__inv_1 _643_ (.A(_334_),
    .Y(_480_));
 sky130_fd_sc_hd__inv_1 _644_ (.A(_350_),
    .Y(_489_));
 sky130_fd_sc_hd__inv_1 _645_ (.A(_360_),
    .Y(_493_));
 sky130_fd_sc_hd__nor2b_1 _646_ (.A(_006_),
    .B_N(net11),
    .Y(_502_));
 sky130_fd_sc_hd__inv_1 _647_ (.A(_385_),
    .Y(_506_));
 sky130_fd_sc_hd__inv_1 _648_ (.A(_115_),
    .Y(_390_));
 sky130_fd_sc_hd__inv_1 _649_ (.A(_131_),
    .Y(_400_));
 sky130_fd_sc_hd__inv_1 _650_ (.A(_143_),
    .Y(_146_));
 sky130_fd_sc_hd__inv_1 _651_ (.A(_163_),
    .Y(_410_));
 sky130_fd_sc_hd__inv_1 _652_ (.A(_189_),
    .Y(_192_));
 sky130_fd_sc_hd__xnor2_1 _653_ (.A(_007_),
    .B(_172_),
    .Y(_418_));
 sky130_fd_sc_hd__inv_1 _654_ (.A(_157_),
    .Y(_415_));
 sky130_fd_sc_hd__inv_1 _655_ (.A(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__a31o_1 _656_ (.A1(_000_),
    .A2(_006_),
    .A3(net11),
    .B1(_419_),
    .X(_227_));
 sky130_fd_sc_hd__inv_1 _657_ (.A(_225_),
    .Y(_436_));
 sky130_fd_sc_hd__nand2b_1 _658_ (.A_N(_431_),
    .B(_008_),
    .Y(_260_));
 sky130_fd_sc_hd__inv_1 _659_ (.A(_238_),
    .Y(_441_));
 sky130_fd_sc_hd__inv_1 _660_ (.A(_248_),
    .Y(_285_));
 sky130_fd_sc_hd__inv_1 _661_ (.A(_284_),
    .Y(_286_));
 sky130_fd_sc_hd__inv_1 _662_ (.A(_257_),
    .Y(_446_));
 sky130_fd_sc_hd__inv_1 _663_ (.A(_258_),
    .Y(_450_));
 sky130_fd_sc_hd__inv_1 _664_ (.A(_306_),
    .Y(_455_));
 sky130_fd_sc_hd__inv_1 _665_ (.A(_274_),
    .Y(_459_));
 sky130_fd_sc_hd__inv_1 _666_ (.A(_310_),
    .Y(_464_));
 sky130_fd_sc_hd__inv_1 _667_ (.A(_290_),
    .Y(_467_));
 sky130_fd_sc_hd__inv_1 _668_ (.A(_335_),
    .Y(_472_));
 sky130_fd_sc_hd__inv_1 _669_ (.A(_313_),
    .Y(_475_));
 sky130_fd_sc_hd__inv_1 _670_ (.A(_351_),
    .Y(_478_));
 sky130_fd_sc_hd__inv_1 _671_ (.A(_361_),
    .Y(_481_));
 sky130_fd_sc_hd__inv_1 _672_ (.A(_375_),
    .Y(_494_));
 sky130_fd_sc_hd__inv_1 _673_ (.A(_374_),
    .Y(_507_));
 sky130_fd_sc_hd__inv_1 _674_ (.A(_409_),
    .Y(_161_));
 sky130_fd_sc_hd__inv_1 _675_ (.A(_420_),
    .Y(_197_));
 sky130_fd_sc_hd__inv_1 _676_ (.A(_259_),
    .Y(_263_));
 sky130_fd_sc_hd__inv_1 _677_ (.A(_398_),
    .Y(_129_));
 sky130_fd_sc_hd__inv_1 _678_ (.A(_169_),
    .Y(_164_));
 sky130_fd_sc_hd__inv_1 _679_ (.A(_422_),
    .Y(_203_));
 sky130_fd_sc_hd__inv_1 _680_ (.A(_428_),
    .Y(_214_));
 sky130_fd_sc_hd__inv_1 _681_ (.A(_433_),
    .Y(_230_));
 sky130_fd_sc_hd__inv_1 _682_ (.A(_465_),
    .Y(_312_));
 sky130_fd_sc_hd__and2_0 _683_ (.A(_000_),
    .B(net1),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 _684_ (.A(net12),
    .X(_010_));
 sky130_fd_sc_hd__a21oi_2 _685_ (.A1(_171_),
    .A2(_413_),
    .B1(_412_),
    .Y(_011_));
 sky130_fd_sc_hd__nand3_1 _686_ (.A(_443_),
    .B(_461_),
    .C(_424_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_1 _687_ (.A(_461_),
    .B(_442_),
    .Y(_013_));
 sky130_fd_sc_hd__nand3_1 _688_ (.A(_443_),
    .B(_461_),
    .C(_423_),
    .Y(_014_));
 sky130_fd_sc_hd__inv_1 _689_ (.A(_460_),
    .Y(_015_));
 sky130_fd_sc_hd__o2111ai_4 _690_ (.A1(_011_),
    .A2(_012_),
    .B1(_013_),
    .C1(_014_),
    .D1(_015_),
    .Y(_016_));
 sky130_fd_sc_hd__xnor2_1 _691_ (.A(_457_),
    .B(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__nand3_1 _692_ (.A(_438_),
    .B(_452_),
    .C(_417_),
    .Y(_018_));
 sky130_fd_sc_hd__nand2_1 _693_ (.A(_452_),
    .B(_437_),
    .Y(_019_));
 sky130_fd_sc_hd__nand3_1 _694_ (.A(_438_),
    .B(_452_),
    .C(_416_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_1 _695_ (.A(_451_),
    .Y(_021_));
 sky130_fd_sc_hd__o2111ai_2 _696_ (.A1(_011_),
    .A2(_018_),
    .B1(_019_),
    .C1(_020_),
    .D1(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__nand2_1 _697_ (.A(_448_),
    .B(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__or2_0 _698_ (.A(_448_),
    .B(_022_),
    .X(_024_));
 sky130_fd_sc_hd__a21oi_1 _699_ (.A1(_023_),
    .A2(_024_),
    .B1(_010_),
    .Y(_025_));
 sky130_fd_sc_hd__a21oi_1 _700_ (.A1(_010_),
    .A2(_017_),
    .B1(_025_),
    .Y(net14));
 sky130_fd_sc_hd__inv_1 _701_ (.A(net12),
    .Y(_026_));
 sky130_fd_sc_hd__nand2b_1 _702_ (.A_N(_167_),
    .B(_417_),
    .Y(_027_));
 sky130_fd_sc_hd__nor2_1 _703_ (.A(_416_),
    .B(_437_),
    .Y(_028_));
 sky130_fd_sc_hd__o21ai_0 _704_ (.A1(_438_),
    .A2(_437_),
    .B1(_452_),
    .Y(_029_));
 sky130_fd_sc_hd__a21oi_1 _705_ (.A1(_027_),
    .A2(_028_),
    .B1(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__o21ai_0 _706_ (.A1(_451_),
    .A2(_030_),
    .B1(_448_),
    .Y(_031_));
 sky130_fd_sc_hd__nand2b_1 _707_ (.A_N(_447_),
    .B(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_1 _708_ (.A(_469_),
    .B(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__inv_1 _709_ (.A(_456_),
    .Y(_034_));
 sky130_fd_sc_hd__nor2b_1 _710_ (.A(_167_),
    .B_N(_424_),
    .Y(_035_));
 sky130_fd_sc_hd__o211ai_2 _711_ (.A1(_423_),
    .A2(_035_),
    .B1(_443_),
    .C1(_461_),
    .Y(_036_));
 sky130_fd_sc_hd__a21oi_1 _712_ (.A1(_461_),
    .A2(_442_),
    .B1(_460_),
    .Y(_037_));
 sky130_fd_sc_hd__o21ai_0 _713_ (.A1(_457_),
    .A2(_456_),
    .B1(_474_),
    .Y(_038_));
 sky130_fd_sc_hd__a31oi_2 _714_ (.A1(_034_),
    .A2(_036_),
    .A3(_037_),
    .B1(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__nand2_1 _715_ (.A(_036_),
    .B(_037_),
    .Y(_040_));
 sky130_fd_sc_hd__a211oi_1 _716_ (.A1(_457_),
    .A2(_040_),
    .B1(_456_),
    .C1(_474_),
    .Y(_041_));
 sky130_fd_sc_hd__o21ai_0 _717_ (.A1(_039_),
    .A2(_041_),
    .B1(_010_),
    .Y(_042_));
 sky130_fd_sc_hd__a21boi_0 _718_ (.A1(_026_),
    .A2(_033_),
    .B1_N(_042_),
    .Y(net15));
 sky130_fd_sc_hd__a21o_1 _719_ (.A1(_457_),
    .A2(_016_),
    .B1(_456_),
    .X(_043_));
 sky130_fd_sc_hd__a21oi_1 _720_ (.A1(_474_),
    .A2(_043_),
    .B1(_473_),
    .Y(_044_));
 sky130_fd_sc_hd__xor2_1 _721_ (.A(_483_),
    .B(_044_),
    .X(_045_));
 sky130_fd_sc_hd__a21o_1 _722_ (.A1(_448_),
    .A2(_022_),
    .B1(_447_),
    .X(_046_));
 sky130_fd_sc_hd__a21oi_1 _723_ (.A1(_469_),
    .A2(_046_),
    .B1(_468_),
    .Y(_047_));
 sky130_fd_sc_hd__xor2_1 _724_ (.A(_477_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__mux2i_1 _725_ (.A0(_045_),
    .A1(_048_),
    .S(_026_),
    .Y(net16));
 sky130_fd_sc_hd__or2_0 _726_ (.A(_473_),
    .B(_482_),
    .X(_049_));
 sky130_fd_sc_hd__o22ai_1 _727_ (.A1(_483_),
    .A2(_482_),
    .B1(_039_),
    .B2(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__xor2_1 _728_ (.A(_496_),
    .B(_050_),
    .X(_051_));
 sky130_fd_sc_hd__nor2_1 _729_ (.A(_447_),
    .B(_451_),
    .Y(_052_));
 sky130_fd_sc_hd__a21oi_1 _730_ (.A1(_477_),
    .A2(_468_),
    .B1(_476_),
    .Y(_053_));
 sky130_fd_sc_hd__nand2_1 _731_ (.A(_052_),
    .B(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _732_ (.A(_448_),
    .B(_447_),
    .Y(_055_));
 sky130_fd_sc_hd__nand2_1 _733_ (.A(_469_),
    .B(_477_),
    .Y(_056_));
 sky130_fd_sc_hd__o21ai_0 _734_ (.A1(_055_),
    .A2(_056_),
    .B1(_053_),
    .Y(_057_));
 sky130_fd_sc_hd__o21ai_1 _735_ (.A1(_030_),
    .A2(_054_),
    .B1(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__xnor2_1 _736_ (.A(_488_),
    .B(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__nand2_1 _737_ (.A(_026_),
    .B(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__o21ai_0 _738_ (.A1(_026_),
    .A2(_051_),
    .B1(_060_),
    .Y(net17));
 sky130_fd_sc_hd__inv_1 _739_ (.A(_488_),
    .Y(_061_));
 sky130_fd_sc_hd__nor3b_1 _740_ (.A(net12),
    .B(_487_),
    .C_N(_501_),
    .Y(_062_));
 sky130_fd_sc_hd__inv_1 _741_ (.A(_509_),
    .Y(_063_));
 sky130_fd_sc_hd__nor3_1 _742_ (.A(_496_),
    .B(_063_),
    .C(_495_),
    .Y(_064_));
 sky130_fd_sc_hd__a21oi_1 _743_ (.A1(_063_),
    .A2(_495_),
    .B1(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__nor2_1 _744_ (.A(net12),
    .B(_501_),
    .Y(_066_));
 sky130_fd_sc_hd__nand2_1 _745_ (.A(_487_),
    .B(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__o21ai_0 _746_ (.A1(_026_),
    .A2(_065_),
    .B1(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__a21oi_1 _747_ (.A1(_061_),
    .A2(_062_),
    .B1(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__nand2_1 _748_ (.A(_010_),
    .B(_509_),
    .Y(_070_));
 sky130_fd_sc_hd__nor2_1 _749_ (.A(_495_),
    .B(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__nand2_1 _750_ (.A(_010_),
    .B(_496_),
    .Y(_072_));
 sky130_fd_sc_hd__nor2_1 _751_ (.A(_509_),
    .B(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__nand4_1 _752_ (.A(_457_),
    .B(_474_),
    .C(_483_),
    .D(_016_),
    .Y(_074_));
 sky130_fd_sc_hd__a21o_1 _753_ (.A1(_474_),
    .A2(_456_),
    .B1(_473_),
    .X(_075_));
 sky130_fd_sc_hd__a21oi_1 _754_ (.A1(_483_),
    .A2(_075_),
    .B1(_482_),
    .Y(_076_));
 sky130_fd_sc_hd__nand2_1 _755_ (.A(_074_),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__mux2i_1 _756_ (.A0(_071_),
    .A1(_073_),
    .S(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__nor3_1 _757_ (.A(_010_),
    .B(_061_),
    .C(_501_),
    .Y(_079_));
 sky130_fd_sc_hd__a21o_1 _758_ (.A1(_469_),
    .A2(_447_),
    .B1(_468_),
    .X(_080_));
 sky130_fd_sc_hd__a21oi_1 _759_ (.A1(_477_),
    .A2(_080_),
    .B1(_476_),
    .Y(_081_));
 sky130_fd_sc_hd__o21ai_0 _760_ (.A1(_023_),
    .A2(_056_),
    .B1(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__mux2i_1 _761_ (.A0(_062_),
    .A1(_079_),
    .S(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__nand3_1 _762_ (.A(_069_),
    .B(_078_),
    .C(_083_),
    .Y(net18));
 sky130_fd_sc_hd__nand2_1 _763_ (.A(_488_),
    .B(_501_),
    .Y(_084_));
 sky130_fd_sc_hd__a21oi_1 _764_ (.A1(_501_),
    .A2(_487_),
    .B1(_500_),
    .Y(_085_));
 sky130_fd_sc_hd__o21ai_0 _765_ (.A1(_058_),
    .A2(_084_),
    .B1(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__xnor2_1 _766_ (.A(_498_),
    .B(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__o21a_1 _767_ (.A1(_483_),
    .A2(_482_),
    .B1(_496_),
    .X(_088_));
 sky130_fd_sc_hd__o21ai_0 _768_ (.A1(_495_),
    .A2(_088_),
    .B1(_509_),
    .Y(_089_));
 sky130_fd_sc_hd__nand2b_1 _769_ (.A_N(_508_),
    .B(_089_),
    .Y(_090_));
 sky130_fd_sc_hd__o41ai_1 _770_ (.A1(_495_),
    .A2(_508_),
    .A3(_039_),
    .A4(_049_),
    .B1(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__xnor2_1 _771_ (.A(_378_),
    .B(_505_),
    .Y(_092_));
 sky130_fd_sc_hd__xnor2_1 _772_ (.A(_381_),
    .B(_384_),
    .Y(_093_));
 sky130_fd_sc_hd__xnor2_1 _773_ (.A(_092_),
    .B(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__xnor2_1 _774_ (.A(_503_),
    .B(_491_),
    .Y(_095_));
 sky130_fd_sc_hd__xnor2_2 _775_ (.A(_094_),
    .B(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__xnor2_1 _776_ (.A(_091_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__mux2i_1 _777_ (.A0(_087_),
    .A1(_097_),
    .S(_010_),
    .Y(net19));
 sky130_fd_sc_hd__clkbuf_1 _778_ (.A(_389_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 _779_ (.A(_392_),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 _780_ (.A(_395_),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 _781_ (.A(_404_),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 _782_ (.A(_406_),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 _783_ (.A(_168_),
    .X(net25));
 sky130_fd_sc_hd__mux2i_1 _784_ (.A0(_417_),
    .A1(_424_),
    .S(_010_),
    .Y(_098_));
 sky130_fd_sc_hd__xor2_1 _785_ (.A(_167_),
    .B(_098_),
    .X(net26));
 sky130_fd_sc_hd__a21o_1 _786_ (.A1(_171_),
    .A2(_413_),
    .B1(_412_),
    .X(_099_));
 sky130_fd_sc_hd__a21oi_1 _787_ (.A1(_424_),
    .A2(_099_),
    .B1(_423_),
    .Y(_100_));
 sky130_fd_sc_hd__xor2_1 _788_ (.A(_443_),
    .B(_100_),
    .X(_101_));
 sky130_fd_sc_hd__a21oi_1 _789_ (.A1(_417_),
    .A2(_099_),
    .B1(_416_),
    .Y(_102_));
 sky130_fd_sc_hd__xnor2_1 _790_ (.A(_438_),
    .B(_102_),
    .Y(_103_));
 sky130_fd_sc_hd__nor2_1 _791_ (.A(_010_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__a21oi_1 _792_ (.A1(_010_),
    .A2(_101_),
    .B1(_104_),
    .Y(net27));
 sky130_fd_sc_hd__o21ai_0 _793_ (.A1(_423_),
    .A2(_035_),
    .B1(_443_),
    .Y(_105_));
 sky130_fd_sc_hd__nand2b_1 _794_ (.A_N(_442_),
    .B(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__xnor2_1 _795_ (.A(_461_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__nand2b_1 _796_ (.A_N(_416_),
    .B(_027_),
    .Y(_108_));
 sky130_fd_sc_hd__a211oi_1 _797_ (.A1(_438_),
    .A2(_108_),
    .B1(_437_),
    .C1(_452_),
    .Y(_109_));
 sky130_fd_sc_hd__or3_1 _798_ (.A(net12),
    .B(_030_),
    .C(_109_),
    .X(_110_));
 sky130_fd_sc_hd__o21ai_0 _799_ (.A1(_026_),
    .A2(_107_),
    .B1(_110_),
    .Y(net28));
 sky130_fd_sc_hd__fa_1 _800_ (.A(_111_),
    .B(_112_),
    .CIN(_113_),
    .COUT(_114_),
    .SUM(_115_));
 sky130_fd_sc_hd__fa_1 _801_ (.A(_116_),
    .B(_117_),
    .CIN(_118_),
    .COUT(_119_),
    .SUM(_120_));
 sky130_fd_sc_hd__fa_1 _802_ (.A(_121_),
    .B(_114_),
    .CIN(_120_),
    .COUT(_122_),
    .SUM(_123_));
 sky130_fd_sc_hd__fa_1 _803_ (.A(_124_),
    .B(_125_),
    .CIN(_126_),
    .COUT(_127_),
    .SUM(_128_));
 sky130_fd_sc_hd__fa_1 _804_ (.A(_128_),
    .B(_119_),
    .CIN(_129_),
    .COUT(_130_),
    .SUM(_131_));
 sky130_fd_sc_hd__fa_1 _805_ (.A(_132_),
    .B(_133_),
    .CIN(_134_),
    .COUT(_135_),
    .SUM(_136_));
 sky130_fd_sc_hd__fa_1 _806_ (.A(_137_),
    .B(_138_),
    .CIN(_139_),
    .COUT(_140_),
    .SUM(_141_));
 sky130_fd_sc_hd__fa_1 _807_ (.A(_136_),
    .B(_141_),
    .CIN(_127_),
    .COUT(_142_),
    .SUM(_143_));
 sky130_fd_sc_hd__fa_1 _808_ (.A(_144_),
    .B(_145_),
    .CIN(_146_),
    .COUT(_147_),
    .SUM(_148_));
 sky130_fd_sc_hd__fa_2 _809_ (.A(_149_),
    .B(_150_),
    .CIN(_151_),
    .COUT(_152_),
    .SUM(_153_));
 sky130_fd_sc_hd__fa_1 _810_ (.A(_154_),
    .B(_155_),
    .CIN(_156_),
    .COUT(_157_),
    .SUM(_158_));
 sky130_fd_sc_hd__fa_1 _811_ (.A(_153_),
    .B(_158_),
    .CIN(_135_),
    .COUT(_159_),
    .SUM(_160_));
 sky130_fd_sc_hd__fa_1 _812_ (.A(_161_),
    .B(_142_),
    .CIN(_160_),
    .COUT(_162_),
    .SUM(_163_));
 sky130_fd_sc_hd__fa_1 _813_ (.A(_164_),
    .B(_165_),
    .CIN(_166_),
    .COUT(_167_),
    .SUM(_168_));
 sky130_fd_sc_hd__fa_1 _814_ (.A(_172_),
    .B(_173_),
    .CIN(_174_),
    .COUT(_175_),
    .SUM(_176_));
 sky130_fd_sc_hd__fa_1 _815_ (.A(_177_),
    .B(_178_),
    .CIN(_179_),
    .COUT(_180_),
    .SUM(_181_));
 sky130_fd_sc_hd__fa_1 _816_ (.A(_152_),
    .B(_181_),
    .CIN(_176_),
    .COUT(_182_),
    .SUM(_183_));
 sky130_fd_sc_hd__fa_1 _817_ (.A(_184_),
    .B(_185_),
    .CIN(_157_),
    .COUT(_186_),
    .SUM(_187_));
 sky130_fd_sc_hd__fa_1 _818_ (.A(_187_),
    .B(_183_),
    .CIN(_159_),
    .COUT(_188_),
    .SUM(_189_));
 sky130_fd_sc_hd__fa_1 _819_ (.A(_190_),
    .B(_191_),
    .CIN(_192_),
    .COUT(_193_),
    .SUM(_194_));
 sky130_fd_sc_hd__fa_1 _820_ (.A(_178_),
    .B(_179_),
    .CIN(_174_),
    .COUT(_195_),
    .SUM(_196_));
 sky130_fd_sc_hd__fa_1 _821_ (.A(_152_),
    .B(_197_),
    .CIN(_196_),
    .COUT(_198_),
    .SUM(_199_));
 sky130_fd_sc_hd__fa_1 _822_ (.A(_177_),
    .B(_200_),
    .CIN(_185_),
    .COUT(_201_),
    .SUM(_202_));
 sky130_fd_sc_hd__fa_1 _823_ (.A(_203_),
    .B(_159_),
    .CIN(_199_),
    .COUT(_204_),
    .SUM(_205_));
 sky130_fd_sc_hd__fa_1 _824_ (.A(_190_),
    .B(_206_),
    .CIN(_191_),
    .COUT(_207_),
    .SUM(_208_));
 sky130_fd_sc_hd__fa_1 _825_ (.A(_209_),
    .B(_210_),
    .CIN(_211_),
    .COUT(_212_),
    .SUM(_213_));
 sky130_fd_sc_hd__fa_1 _826_ (.A(_175_),
    .B(_214_),
    .CIN(_215_),
    .COUT(_216_),
    .SUM(_217_));
 sky130_fd_sc_hd__fa_1 _827_ (.A(_218_),
    .B(_180_),
    .CIN(_219_),
    .COUT(_220_),
    .SUM(_221_));
 sky130_fd_sc_hd__fa_1 _828_ (.A(_182_),
    .B(_217_),
    .CIN(_221_),
    .COUT(_222_),
    .SUM(_223_));
 sky130_fd_sc_hd__fa_1 _829_ (.A(_186_),
    .B(_223_),
    .CIN(_188_),
    .COUT(_224_),
    .SUM(_225_));
 sky130_fd_sc_hd__fa_1 _830_ (.A(_226_),
    .B(_213_),
    .CIN(_227_),
    .COUT(_228_),
    .SUM(_229_));
 sky130_fd_sc_hd__fa_1 _831_ (.A(_230_),
    .B(_195_),
    .CIN(_201_),
    .COUT(_231_),
    .SUM(_232_));
 sky130_fd_sc_hd__fa_1 _832_ (.A(_198_),
    .B(_233_),
    .CIN(_232_),
    .COUT(_234_),
    .SUM(_235_));
 sky130_fd_sc_hd__fa_1 _833_ (.A(_236_),
    .B(_235_),
    .CIN(_204_),
    .COUT(_237_),
    .SUM(_238_));
 sky130_fd_sc_hd__fa_1 _834_ (.A(_240_),
    .B(_241_),
    .CIN(_242_),
    .COUT(_243_),
    .SUM(_244_));
 sky130_fd_sc_hd__fa_1 _835_ (.A(_245_),
    .B(_246_),
    .CIN(_247_),
    .COUT(_248_),
    .SUM(_249_));
 sky130_fd_sc_hd__fa_1 _836_ (.A(_250_),
    .B(_251_),
    .CIN(_252_),
    .COUT(_253_),
    .SUM(_254_));
 sky130_fd_sc_hd__fa_1 _837_ (.A(_216_),
    .B(_249_),
    .CIN(_254_),
    .COUT(_255_),
    .SUM(_256_));
 sky130_fd_sc_hd__fa_1 _838_ (.A(_222_),
    .B(_256_),
    .CIN(_220_),
    .COUT(_257_),
    .SUM(_258_));
 sky130_fd_sc_hd__fa_1 _839_ (.A(_259_),
    .B(_244_),
    .CIN(_260_),
    .COUT(_261_),
    .SUM(_262_));
 sky130_fd_sc_hd__fa_1 _840_ (.A(_212_),
    .B(_264_),
    .CIN(_265_),
    .COUT(_266_),
    .SUM(_267_));
 sky130_fd_sc_hd__fa_1 _841_ (.A(_268_),
    .B(_269_),
    .CIN(_270_),
    .COUT(_271_),
    .SUM(_272_));
 sky130_fd_sc_hd__fa_1 _842_ (.A(_234_),
    .B(_272_),
    .CIN(_231_),
    .COUT(_273_),
    .SUM(_274_));
 sky130_fd_sc_hd__fa_2 _843_ (.A(_275_),
    .B(_276_),
    .CIN(_277_),
    .COUT(_278_),
    .SUM(_279_));
 sky130_fd_sc_hd__fa_1 _844_ (.A(_280_),
    .B(_281_),
    .CIN(_282_),
    .COUT(_283_),
    .SUM(_284_));
 sky130_fd_sc_hd__fa_1 _845_ (.A(_279_),
    .B(_285_),
    .CIN(_286_),
    .COUT(_287_),
    .SUM(_288_));
 sky130_fd_sc_hd__fa_1 _846_ (.A(_255_),
    .B(_289_),
    .CIN(_253_),
    .COUT(_290_),
    .SUM(_291_));
 sky130_fd_sc_hd__fa_1 _847_ (.A(_279_),
    .B(_259_),
    .CIN(_292_),
    .COUT(_293_),
    .SUM(_294_));
 sky130_fd_sc_hd__fa_1 _848_ (.A(_243_),
    .B(_295_),
    .CIN(_296_),
    .COUT(_297_),
    .SUM(_298_));
 sky130_fd_sc_hd__fa_1 _849_ (.A(_299_),
    .B(_300_),
    .CIN(_301_),
    .COUT(_302_),
    .SUM(_303_));
 sky130_fd_sc_hd__fa_1 _850_ (.A(_303_),
    .B(_271_),
    .CIN(_304_),
    .COUT(_305_),
    .SUM(_306_));
 sky130_fd_sc_hd__fa_1 _851_ (.A(_307_),
    .B(_278_),
    .CIN(_308_),
    .COUT(_309_),
    .SUM(_310_));
 sky130_fd_sc_hd__fa_1 _852_ (.A(_283_),
    .B(_311_),
    .CIN(_312_),
    .COUT(_313_),
    .SUM(_314_));
 sky130_fd_sc_hd__fa_1 _853_ (.A(_315_),
    .B(_316_),
    .CIN(_317_),
    .COUT(_318_),
    .SUM(_319_));
 sky130_fd_sc_hd__fa_1 _854_ (.A(_263_),
    .B(_320_),
    .CIN(_321_),
    .COUT(_322_),
    .SUM(_323_));
 sky130_fd_sc_hd__fa_1 _855_ (.A(_324_),
    .B(_325_),
    .CIN(_326_),
    .COUT(_327_),
    .SUM(_328_));
 sky130_fd_sc_hd__fa_1 _856_ (.A(_323_),
    .B(_329_),
    .CIN(_330_),
    .COUT(_331_),
    .SUM(_332_));
 sky130_fd_sc_hd__fa_1 _857_ (.A(_333_),
    .B(_302_),
    .CIN(_332_),
    .COUT(_334_),
    .SUM(_335_));
 sky130_fd_sc_hd__fa_1 _858_ (.A(_336_),
    .B(_337_),
    .CIN(_338_),
    .COUT(_339_),
    .SUM(_340_));
 sky130_fd_sc_hd__fa_1 _859_ (.A(_341_),
    .B(_342_),
    .CIN(_343_),
    .COUT(_344_),
    .SUM(_345_));
 sky130_fd_sc_hd__fa_2 _860_ (.A(_315_),
    .B(_316_),
    .CIN(_346_),
    .COUT(_347_),
    .SUM(_348_));
 sky130_fd_sc_hd__fa_4 _861_ (.A(_263_),
    .B(_320_),
    .CIN(_349_),
    .COUT(_350_),
    .SUM(_351_));
 sky130_fd_sc_hd__fa_1 _862_ (.A(_352_),
    .B(_353_),
    .CIN(_318_),
    .COUT(_354_),
    .SUM(_355_));
 sky130_fd_sc_hd__fa_1 _863_ (.A(_356_),
    .B(_322_),
    .CIN(_351_),
    .COUT(_357_),
    .SUM(_358_));
 sky130_fd_sc_hd__fa_1 _864_ (.A(_358_),
    .B(_331_),
    .CIN(_359_),
    .COUT(_360_),
    .SUM(_361_));
 sky130_fd_sc_hd__fa_1 _865_ (.A(_362_),
    .B(_363_),
    .CIN(_339_),
    .COUT(_364_),
    .SUM(_365_));
 sky130_fd_sc_hd__fa_1 _866_ (.A(_366_),
    .B(_347_),
    .CIN(_367_),
    .COUT(_368_),
    .SUM(_369_));
 sky130_fd_sc_hd__fa_1 _867_ (.A(_350_),
    .B(_351_),
    .CIN(_370_),
    .COUT(_371_),
    .SUM(_372_));
 sky130_fd_sc_hd__fa_1 _868_ (.A(_357_),
    .B(_373_),
    .CIN(_372_),
    .COUT(_374_),
    .SUM(_375_));
 sky130_fd_sc_hd__fa_1 _869_ (.A(_347_),
    .B(_376_),
    .CIN(_377_),
    .COUT(_378_),
    .SUM(_379_));
 sky130_fd_sc_hd__fa_1 _870_ (.A(_350_),
    .B(_380_),
    .CIN(_351_),
    .COUT(_381_),
    .SUM(_382_));
 sky130_fd_sc_hd__fa_1 _871_ (.A(_383_),
    .B(_382_),
    .CIN(_371_),
    .COUT(_384_),
    .SUM(_385_));
 sky130_fd_sc_hd__ha_1 _872_ (.A(_386_),
    .B(_387_),
    .COUT(_388_),
    .SUM(_389_));
 sky130_fd_sc_hd__ha_1 _873_ (.A(_388_),
    .B(_390_),
    .COUT(_391_),
    .SUM(_392_));
 sky130_fd_sc_hd__ha_1 _874_ (.A(_393_),
    .B(_391_),
    .COUT(_394_),
    .SUM(_395_));
 sky130_fd_sc_hd__ha_1 _875_ (.A(_396_),
    .B(_397_),
    .COUT(_144_),
    .SUM(_398_));
 sky130_fd_sc_hd__ha_1 _876_ (.A(_399_),
    .B(_400_),
    .COUT(_401_),
    .SUM(_402_));
 sky130_fd_sc_hd__ha_1 _877_ (.A(_402_),
    .B(_394_),
    .COUT(_403_),
    .SUM(_404_));
 sky130_fd_sc_hd__ha_1 _878_ (.A(_401_),
    .B(_148_),
    .COUT(_170_),
    .SUM(_405_));
 sky130_fd_sc_hd__ha_1 _879_ (.A(_403_),
    .B(_405_),
    .COUT(_171_),
    .SUM(_406_));
 sky130_fd_sc_hd__ha_1 _880_ (.A(_407_),
    .B(_408_),
    .COUT(_191_),
    .SUM(_409_));
 sky130_fd_sc_hd__ha_1 _881_ (.A(_147_),
    .B(_410_),
    .COUT(_411_),
    .SUM(_169_));
 sky130_fd_sc_hd__ha_1 _882_ (.A(_169_),
    .B(_170_),
    .COUT(_412_),
    .SUM(_413_));
 sky130_fd_sc_hd__ha_1 _883_ (.A(_194_),
    .B(_411_),
    .COUT(_416_),
    .SUM(_417_));
 sky130_fd_sc_hd__ha_1 _884_ (.A(_414_),
    .B(_418_),
    .COUT(_419_),
    .SUM(_420_));
 sky130_fd_sc_hd__ha_1 _885_ (.A(_421_),
    .B(_415_),
    .COUT(_239_),
    .SUM(_422_));
 sky130_fd_sc_hd__ha_1 _886_ (.A(_208_),
    .B(_411_),
    .COUT(_423_),
    .SUM(_424_));
 sky130_fd_sc_hd__ha_1 _887_ (.A(_425_),
    .B(_426_),
    .COUT(_427_),
    .SUM(_428_));
 sky130_fd_sc_hd__ha_1 _888_ (.A(_426_),
    .B(_430_),
    .COUT(_431_),
    .SUM(_226_));
 sky130_fd_sc_hd__ha_1 _889_ (.A(_429_),
    .B(_432_),
    .COUT(_265_),
    .SUM(_433_));
 sky130_fd_sc_hd__ha_1 _890_ (.A(_193_),
    .B(_436_),
    .COUT(_437_),
    .SUM(_438_));
 sky130_fd_sc_hd__ha_1 _891_ (.A(_430_),
    .B(_434_),
    .COUT(_439_),
    .SUM(_259_));
 sky130_fd_sc_hd__ha_1 _892_ (.A(_435_),
    .B(_440_),
    .COUT(_295_),
    .SUM(_264_));
 sky130_fd_sc_hd__ha_1 _893_ (.A(_207_),
    .B(_441_),
    .COUT(_442_),
    .SUM(_443_));
 sky130_fd_sc_hd__ha_1 _894_ (.A(_445_),
    .B(_446_),
    .COUT(_447_),
    .SUM(_448_));
 sky130_fd_sc_hd__ha_1 _895_ (.A(_449_),
    .B(_450_),
    .COUT(_451_),
    .SUM(_452_));
 sky130_fd_sc_hd__ha_1 _896_ (.A(_444_),
    .B(_453_),
    .COUT(_326_),
    .SUM(_296_));
 sky130_fd_sc_hd__ha_1 _897_ (.A(_454_),
    .B(_455_),
    .COUT(_456_),
    .SUM(_457_));
 sky130_fd_sc_hd__ha_1 _898_ (.A(_458_),
    .B(_459_),
    .COUT(_460_),
    .SUM(_461_));
 sky130_fd_sc_hd__ha_1 _899_ (.A(_316_),
    .B(_317_),
    .COUT(_336_),
    .SUM(_462_));
 sky130_fd_sc_hd__ha_1 _900_ (.A(_462_),
    .B(_464_),
    .COUT(_343_),
    .SUM(_465_));
 sky130_fd_sc_hd__ha_1 _901_ (.A(_466_),
    .B(_467_),
    .COUT(_468_),
    .SUM(_469_));
 sky130_fd_sc_hd__ha_1 _902_ (.A(_463_),
    .B(_470_),
    .COUT(_352_),
    .SUM(_325_));
 sky130_fd_sc_hd__ha_1 _903_ (.A(_471_),
    .B(_472_),
    .COUT(_473_),
    .SUM(_474_));
 sky130_fd_sc_hd__ha_1 _904_ (.A(_340_),
    .B(_346_),
    .COUT(_362_),
    .SUM(_342_));
 sky130_fd_sc_hd__ha_1 _905_ (.A(_345_),
    .B(_475_),
    .COUT(_476_),
    .SUM(_477_));
 sky130_fd_sc_hd__ha_1 _906_ (.A(_479_),
    .B(_337_),
    .COUT(_367_),
    .SUM(_353_));
 sky130_fd_sc_hd__ha_1 _907_ (.A(_480_),
    .B(_481_),
    .COUT(_482_),
    .SUM(_483_));
 sky130_fd_sc_hd__ha_1 _908_ (.A(_484_),
    .B(_485_),
    .COUT(_486_),
    .SUM(_363_));
 sky130_fd_sc_hd__ha_1 _909_ (.A(_365_),
    .B(_344_),
    .COUT(_487_),
    .SUM(_488_));
 sky130_fd_sc_hd__ha_1 _910_ (.A(_489_),
    .B(_478_),
    .COUT(_490_),
    .SUM(_491_));
 sky130_fd_sc_hd__ha_1 _911_ (.A(_492_),
    .B(_485_),
    .COUT(_377_),
    .SUM(_366_));
 sky130_fd_sc_hd__ha_1 _912_ (.A(_493_),
    .B(_494_),
    .COUT(_495_),
    .SUM(_496_));
 sky130_fd_sc_hd__ha_1 _913_ (.A(_486_),
    .B(_497_),
    .COUT(_498_),
    .SUM(_499_));
 sky130_fd_sc_hd__ha_1 _914_ (.A(_499_),
    .B(_364_),
    .COUT(_500_),
    .SUM(_501_));
 sky130_fd_sc_hd__ha_1 _915_ (.A(_502_),
    .B(_485_),
    .COUT(_503_),
    .SUM(_376_));
 sky130_fd_sc_hd__ha_1 _916_ (.A(_347_),
    .B(_376_),
    .COUT(_504_),
    .SUM(_505_));
 sky130_fd_sc_hd__ha_1 _917_ (.A(_506_),
    .B(_507_),
    .COUT(_508_),
    .SUM(_509_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_74 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(a[5]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(a[6]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[7]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(b[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(b[2]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(b[3]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(b[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(b[5]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input10 (.A(b[6]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(b[7]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(sign_mode),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net13),
    .X(product[0]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .X(product[10]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(product[11]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(product[12]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(product[13]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(product[14]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(product[15]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(product[1]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(product[2]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(product[3]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(product[4]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(product[5]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(product[6]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(product[7]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(product[8]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(product[9]));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_170 ();
endmodule
