module performance_counter (clear,
    clk,
    enable,
    rst_n,
    all_counts,
    count_value,
    counter_sel,
    event_inc);
 input clear;
 input clk;
 input enable;
 input rst_n;
 output [255:0] all_counts;
 output [31:0] count_value;
 input [7:0] counter_sel;
 input [7:0] event_inc;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire \prev_event_inc[0] ;
 wire \prev_event_inc[1] ;
 wire \prev_event_inc[2] ;
 wire \prev_event_inc[3] ;
 wire \prev_event_inc[4] ;
 wire \prev_event_inc[5] ;
 wire \prev_event_inc[6] ;
 wire \prev_event_inc[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net304;
 wire net305;
 wire net306;
 wire net307;

 gf180mcu_fd_sc_mcu9t5v0__inv_4 _1458_ (.I(net1),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1459_ (.I(_1126_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1460_ (.I(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1461_ (.I(\prev_event_inc[0] ),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1462_ (.A1(net6),
    .A2(net7),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1463_ (.A1(_1129_),
    .A2(_1130_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1464_ (.A1(net16),
    .A2(_1131_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1465_ (.A1(_1128_),
    .A2(_1132_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1466_ (.I(net6),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1467_ (.I(\prev_event_inc[3] ),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1468_ (.A1(net269),
    .A2(net270),
    .A3(_1454_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1469_ (.A1(_1133_),
    .A2(net10),
    .A3(_1134_),
    .A4(_1135_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1470_ (.I(_1136_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1471_ (.A1(net17),
    .A2(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1472_ (.A1(_1128_),
    .A2(_1138_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1473_ (.A1(net267),
    .A2(net268),
    .A3(net269),
    .A4(net270),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _1474_ (.A1(_1133_),
    .A2(net10),
    .A3(_1134_),
    .A4(_1139_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1475_ (.A1(net17),
    .A2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1476_ (.A1(net18),
    .A2(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1477_ (.A1(_1128_),
    .A2(_1142_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1478_ (.I(net1),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1479_ (.A1(net17),
    .A2(net18),
    .A3(_1137_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1480_ (.A1(net19),
    .A2(_1144_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1481_ (.A1(_1143_),
    .A2(_1145_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1482_ (.A1(net17),
    .A2(net18),
    .A3(net19),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1483_ (.A1(_1140_),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1484_ (.A1(net20),
    .A2(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1485_ (.A1(_1128_),
    .A2(_1148_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1486_ (.A1(net20),
    .A2(_1137_),
    .A3(_1146_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1487_ (.A1(net21),
    .A2(_1149_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1488_ (.A1(_1128_),
    .A2(_1150_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1489_ (.A1(net20),
    .A2(net21),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1490_ (.A1(_1140_),
    .A2(_1146_),
    .A3(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1491_ (.A1(net22),
    .A2(_1152_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1492_ (.A1(_1128_),
    .A2(_1153_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1493_ (.A1(net22),
    .A2(_1137_),
    .A3(_1146_),
    .A4(_1151_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1494_ (.A1(net23),
    .A2(_1154_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1495_ (.A1(_1128_),
    .A2(_1155_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1496_ (.A1(net20),
    .A2(net21),
    .A3(net22),
    .A4(net23),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1497_ (.A1(_1140_),
    .A2(_1146_),
    .A3(_1156_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1498_ (.A1(net24),
    .A2(_1157_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1499_ (.A1(_1128_),
    .A2(_1158_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1500_ (.A1(net24),
    .A2(_1137_),
    .A3(_1146_),
    .A4(_1156_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1501_ (.A1(net25),
    .A2(_1159_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1502_ (.A1(_1128_),
    .A2(_1160_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1503_ (.A1(net24),
    .A2(net25),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1504_ (.A1(_1156_),
    .A2(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1505_ (.A1(_1140_),
    .A2(_1146_),
    .A3(_1162_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1506_ (.A1(net26),
    .A2(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1507_ (.A1(_1128_),
    .A2(_1164_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1508_ (.I(_1127_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1509_ (.A1(_1129_),
    .A2(_1444_),
    .A3(net194),
    .A4(_1130_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1510_ (.I(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1511_ (.A1(net205),
    .A2(net216),
    .A3(net227),
    .A4(net238),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1512_ (.A1(net249),
    .A2(net260),
    .A3(_1168_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1513_ (.I(_1169_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1514_ (.A1(net271),
    .A2(_1167_),
    .A3(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1515_ (.A1(net27),
    .A2(_1171_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1516_ (.A1(_1165_),
    .A2(_1172_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1517_ (.A1(net26),
    .A2(_1137_),
    .A3(_1146_),
    .A4(_1162_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1518_ (.A1(net28),
    .A2(_1173_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1519_ (.A1(_1165_),
    .A2(_1174_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1520_ (.A1(net26),
    .A2(net28),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1521_ (.A1(_1146_),
    .A2(_1156_),
    .A3(_1161_),
    .A4(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1522_ (.I(_1176_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1523_ (.A1(_1140_),
    .A2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1524_ (.A1(net29),
    .A2(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1525_ (.A1(_1165_),
    .A2(_1179_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1526_ (.A1(_1146_),
    .A2(_1175_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1527_ (.A1(net29),
    .A2(_1136_),
    .A3(_1162_),
    .A4(_1180_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1528_ (.A1(net30),
    .A2(_1181_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1529_ (.A1(_1165_),
    .A2(_1182_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1530_ (.A1(net29),
    .A2(net30),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1531_ (.A1(_1140_),
    .A2(_1162_),
    .A3(_1180_),
    .A4(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1532_ (.A1(net31),
    .A2(_1184_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1533_ (.A1(_1165_),
    .A2(_1185_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1534_ (.A1(net31),
    .A2(_1136_),
    .A3(_1177_),
    .A4(_1183_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1535_ (.A1(net32),
    .A2(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1536_ (.A1(_1165_),
    .A2(_1187_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1537_ (.A1(net29),
    .A2(net30),
    .A3(net31),
    .A4(net32),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1538_ (.A1(_1140_),
    .A2(_1177_),
    .A3(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1539_ (.A1(net33),
    .A2(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1540_ (.A1(_1165_),
    .A2(_1190_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1541_ (.A1(net33),
    .A2(_1136_),
    .A3(_1177_),
    .A4(_1188_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1542_ (.A1(net34),
    .A2(_1191_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1543_ (.A1(_1165_),
    .A2(_1192_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1544_ (.A1(net33),
    .A2(net34),
    .A3(_1188_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1545_ (.A1(_1140_),
    .A2(_1176_),
    .A3(_1193_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1546_ (.A1(net35),
    .A2(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1547_ (.A1(_1165_),
    .A2(_1195_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1548_ (.A1(net35),
    .A2(_1136_),
    .A3(_1177_),
    .A4(_1193_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1549_ (.A1(net36),
    .A2(_1196_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1550_ (.A1(_1165_),
    .A2(_1197_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1551_ (.I(_1126_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1552_ (.A1(_1198_),
    .A2(net37),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1553_ (.I(net1),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1554_ (.A1(_1200_),
    .A2(net37),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1555_ (.A1(net35),
    .A2(net36),
    .A3(_1194_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1556_ (.I0(_1199_),
    .I1(_1201_),
    .S(_1202_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1557_ (.I(_1127_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1558_ (.A1(net16),
    .A2(net127),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1559_ (.A1(_1129_),
    .A2(net194),
    .A3(_1130_),
    .A4(_1204_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1560_ (.A1(net271),
    .A2(net27),
    .A3(_1169_),
    .A4(_1205_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1561_ (.A1(net38),
    .A2(_1206_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1562_ (.A1(_1203_),
    .A2(_1207_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1563_ (.A1(net35),
    .A2(net36),
    .A3(net37),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1564_ (.A1(_1137_),
    .A2(_1177_),
    .A3(_1193_),
    .A4(_1208_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1565_ (.A1(net39),
    .A2(_1209_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1566_ (.A1(_1203_),
    .A2(_1210_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1567_ (.A1(_1198_),
    .A2(net40),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1568_ (.A1(_1200_),
    .A2(net40),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1569_ (.A1(net35),
    .A2(net36),
    .A3(net37),
    .A4(net39),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1570_ (.A1(_1194_),
    .A2(_1213_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1571_ (.I0(_1211_),
    .I1(_1212_),
    .S(_1214_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1572_ (.A1(net40),
    .A2(_1213_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1573_ (.A1(_1137_),
    .A2(_1177_),
    .A3(_1193_),
    .A4(_1215_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1574_ (.A1(net41),
    .A2(_1216_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1575_ (.A1(_1203_),
    .A2(_1217_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1576_ (.A1(net40),
    .A2(net41),
    .A3(_1213_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1577_ (.A1(_1140_),
    .A2(_1177_),
    .A3(_1193_),
    .A4(_1218_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1578_ (.A1(net42),
    .A2(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1579_ (.A1(_1203_),
    .A2(_1220_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1580_ (.A1(net40),
    .A2(net41),
    .A3(net42),
    .A4(_1213_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1581_ (.A1(_1137_),
    .A2(_1177_),
    .A3(_1193_),
    .A4(_1221_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1582_ (.A1(net43),
    .A2(_1222_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1583_ (.A1(_1203_),
    .A2(_1223_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1584_ (.A1(_1200_),
    .A2(net44),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1585_ (.A1(_1126_),
    .A2(net44),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1586_ (.A1(net43),
    .A2(_1194_),
    .A3(_1221_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1587_ (.I0(_1224_),
    .I1(_1225_),
    .S(_1226_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1588_ (.A1(net40),
    .A2(net41),
    .A3(net42),
    .A4(net43),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1589_ (.A1(net44),
    .A2(_1213_),
    .A3(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1590_ (.A1(_1137_),
    .A2(_1177_),
    .A3(_1193_),
    .A4(_1228_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1591_ (.A1(net45),
    .A2(_1229_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1592_ (.A1(_1203_),
    .A2(_1230_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1593_ (.A1(_1198_),
    .A2(net46),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1594_ (.A1(_1200_),
    .A2(net46),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1595_ (.A1(net45),
    .A2(_1194_),
    .A3(_1228_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1596_ (.I0(_1231_),
    .I1(_1232_),
    .S(_1233_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1597_ (.I(net47),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1598_ (.I(\prev_event_inc[4] ),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1599_ (.A1(net6),
    .A2(net11),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1600_ (.A1(_1235_),
    .A2(_1236_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1601_ (.A1(_1234_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1602_ (.A1(_1203_),
    .A2(_1238_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1603_ (.I0(net48),
    .I1(_1453_),
    .S(_1237_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1604_ (.A1(_1203_),
    .A2(_1239_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _1605_ (.A1(net271),
    .A2(net27),
    .A3(net38),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1606_ (.A1(_1167_),
    .A2(_1170_),
    .A3(_1240_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1607_ (.A1(net49),
    .A2(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1608_ (.A1(_1203_),
    .A2(_1242_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1609_ (.I(net50),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1610_ (.A1(_1452_),
    .A2(_1237_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1611_ (.A1(_1243_),
    .A2(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1612_ (.A1(_1203_),
    .A2(_1245_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1613_ (.I(_1127_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1614_ (.I(net51),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1615_ (.A1(net47),
    .A2(net48),
    .A3(net50),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1616_ (.A1(_1235_),
    .A2(_1236_),
    .A3(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1617_ (.A1(_1247_),
    .A2(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1618_ (.A1(_1246_),
    .A2(_1250_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1619_ (.I(net52),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1620_ (.A1(_1235_),
    .A2(net50),
    .A3(_1452_),
    .A4(_1236_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1621_ (.I(_1252_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1622_ (.A1(net51),
    .A2(_1253_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1623_ (.A1(_1251_),
    .A2(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1624_ (.A1(_1246_),
    .A2(_1255_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1625_ (.I(net53),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1626_ (.A1(net51),
    .A2(net52),
    .A3(_1249_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1627_ (.A1(_1256_),
    .A2(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1628_ (.A1(_1143_),
    .A2(_1258_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1629_ (.I(net54),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1630_ (.A1(net51),
    .A2(net52),
    .A3(net53),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1631_ (.A1(_1253_),
    .A2(_1260_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1632_ (.A1(_1259_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1633_ (.A1(_1246_),
    .A2(_1262_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1634_ (.I(net55),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1635_ (.A1(net51),
    .A2(net52),
    .A3(net53),
    .A4(net54),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1636_ (.A1(_1235_),
    .A2(_1236_),
    .A3(_1248_),
    .A4(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1637_ (.A1(_1263_),
    .A2(_1265_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1638_ (.A1(_1246_),
    .A2(_1266_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1639_ (.I(net56),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1640_ (.A1(net55),
    .A2(_1253_),
    .A3(_1264_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1641_ (.A1(_1267_),
    .A2(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1642_ (.A1(_1246_),
    .A2(_1269_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1643_ (.I(net57),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1644_ (.A1(net55),
    .A2(net56),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1645_ (.A1(_1265_),
    .A2(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1646_ (.A1(_1270_),
    .A2(_1272_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1647_ (.A1(_1246_),
    .A2(_1273_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1648_ (.I(net58),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1649_ (.A1(net57),
    .A2(_1252_),
    .A3(_1264_),
    .A4(_1271_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1650_ (.A1(_1274_),
    .A2(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1651_ (.A1(_1246_),
    .A2(_1276_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1652_ (.I(net59),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1653_ (.A1(net55),
    .A2(net56),
    .A3(net57),
    .A4(net58),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1654_ (.A1(_1265_),
    .A2(_1278_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1655_ (.A1(_1277_),
    .A2(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1656_ (.A1(_1246_),
    .A2(_1280_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1657_ (.A1(_1129_),
    .A2(net194),
    .A3(_1130_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1658_ (.A1(net16),
    .A2(net127),
    .A3(net260),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1659_ (.A1(net249),
    .A2(_1168_),
    .A3(_1240_),
    .A4(_1282_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1660_ (.A1(net49),
    .A2(_1281_),
    .A3(_1283_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1661_ (.A1(net60),
    .A2(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1662_ (.A1(_1246_),
    .A2(_1285_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1663_ (.I(net61),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1664_ (.A1(net59),
    .A2(_1252_),
    .A3(_1264_),
    .A4(_1278_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1665_ (.A1(_1286_),
    .A2(_1287_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1666_ (.A1(_1246_),
    .A2(_1288_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1667_ (.I(_1127_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1668_ (.I(net62),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1669_ (.A1(net59),
    .A2(net61),
    .A3(_1265_),
    .A4(_1278_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1670_ (.A1(_1290_),
    .A2(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1671_ (.A1(_1289_),
    .A2(_1292_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1672_ (.I(net63),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1673_ (.A1(net54),
    .A2(net59),
    .A3(net61),
    .A4(net62),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1674_ (.A1(_1260_),
    .A2(_1278_),
    .A3(_1294_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1675_ (.A1(_1253_),
    .A2(_1295_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1676_ (.A1(_1293_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1677_ (.A1(_1289_),
    .A2(_1297_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1678_ (.I(net64),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1679_ (.A1(net59),
    .A2(net61),
    .A3(net62),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1680_ (.A1(net63),
    .A2(_1265_),
    .A3(_1278_),
    .A4(_1299_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1681_ (.A1(_1298_),
    .A2(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1682_ (.A1(_1289_),
    .A2(_1301_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1683_ (.I(net65),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1684_ (.A1(net63),
    .A2(net64),
    .A3(_1252_),
    .A4(_1295_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1685_ (.A1(_1302_),
    .A2(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1686_ (.A1(_1289_),
    .A2(_1304_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1687_ (.I(net66),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1688_ (.A1(net63),
    .A2(net64),
    .A3(net65),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1689_ (.A1(_1265_),
    .A2(_1278_),
    .A3(_1299_),
    .A4(_1306_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1690_ (.A1(_1305_),
    .A2(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1691_ (.A1(_1289_),
    .A2(_1308_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1692_ (.I(net67),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1693_ (.A1(net63),
    .A2(net64),
    .A3(net65),
    .A4(net66),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1694_ (.A1(_1253_),
    .A2(_1295_),
    .A3(_1310_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1695_ (.A1(_1309_),
    .A2(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1696_ (.A1(_1289_),
    .A2(_1312_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1697_ (.I(net68),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1698_ (.A1(net67),
    .A2(_1310_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1699_ (.A1(_1265_),
    .A2(_1278_),
    .A3(_1299_),
    .A4(_1314_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1700_ (.A1(_1313_),
    .A2(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1701_ (.A1(_1289_),
    .A2(_1316_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1702_ (.I(net69),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _1703_ (.I(_1314_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1704_ (.A1(net68),
    .A2(_1260_),
    .A3(_1278_),
    .A4(_1294_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1705_ (.A1(_1253_),
    .A2(_1318_),
    .A3(_1319_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1706_ (.A1(_1317_),
    .A2(_1320_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1707_ (.A1(_1289_),
    .A2(_1321_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1708_ (.I(net70),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1709_ (.A1(net69),
    .A2(_1249_),
    .A3(_1314_),
    .A4(_1319_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1710_ (.A1(_1322_),
    .A2(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1711_ (.A1(_1289_),
    .A2(_1324_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1712_ (.A1(net49),
    .A2(net60),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1713_ (.A1(_1167_),
    .A2(_1170_),
    .A3(_1240_),
    .A4(_1325_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1714_ (.A1(net71),
    .A2(_1326_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1715_ (.A1(_1289_),
    .A2(_1327_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1716_ (.I(_1127_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1717_ (.I(net72),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1718_ (.A1(net69),
    .A2(net70),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1719_ (.A1(_1253_),
    .A2(_1318_),
    .A3(_1319_),
    .A4(_1330_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1720_ (.A1(_1329_),
    .A2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1721_ (.A1(_1328_),
    .A2(_1332_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1722_ (.I(net73),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1723_ (.A1(net68),
    .A2(net69),
    .A3(net70),
    .A4(net72),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1724_ (.A1(_1260_),
    .A2(_1278_),
    .A3(_1294_),
    .A4(_1334_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1725_ (.A1(_1249_),
    .A2(_1318_),
    .A3(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1726_ (.A1(_1333_),
    .A2(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1727_ (.A1(_1328_),
    .A2(_1337_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1728_ (.I(net74),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1729_ (.A1(net73),
    .A2(_1252_),
    .A3(_1314_),
    .A4(_1335_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1730_ (.A1(_1338_),
    .A2(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1731_ (.A1(_1328_),
    .A2(_1340_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1732_ (.I(net75),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1733_ (.A1(net73),
    .A2(net74),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1734_ (.A1(_1249_),
    .A2(_1318_),
    .A3(_1335_),
    .A4(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1735_ (.A1(_1341_),
    .A2(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1736_ (.A1(_1328_),
    .A2(_1344_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1737_ (.I(net76),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1738_ (.A1(net75),
    .A2(_1342_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1739_ (.A1(_1253_),
    .A2(_1318_),
    .A3(_1335_),
    .A4(_1346_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1740_ (.A1(_1345_),
    .A2(_1347_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1741_ (.A1(_1328_),
    .A2(_1348_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1742_ (.I(net77),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1743_ (.A1(net73),
    .A2(net74),
    .A3(net75),
    .A4(net76),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1744_ (.A1(_1249_),
    .A2(_1318_),
    .A3(_1335_),
    .A4(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1745_ (.A1(_1349_),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1746_ (.A1(_1328_),
    .A2(_1352_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1747_ (.I(net78),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1748_ (.A1(net77),
    .A2(_1350_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1749_ (.A1(_1253_),
    .A2(_1318_),
    .A3(_1335_),
    .A4(_1354_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1750_ (.A1(_1353_),
    .A2(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1751_ (.A1(_1328_),
    .A2(_1356_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1752_ (.I(net79),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1753_ (.A1(net77),
    .A2(net78),
    .A3(_1350_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1754_ (.A1(_1249_),
    .A2(_1318_),
    .A3(_1335_),
    .A4(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1755_ (.A1(_1357_),
    .A2(_1359_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1756_ (.A1(_1328_),
    .A2(_1360_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1757_ (.I(net80),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1758_ (.A1(net77),
    .A2(net78),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1759_ (.A1(net79),
    .A2(_1350_),
    .A3(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1760_ (.A1(_1253_),
    .A2(_1318_),
    .A3(_1335_),
    .A4(_1363_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1761_ (.A1(_1361_),
    .A2(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1762_ (.A1(_1328_),
    .A2(_1365_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1763_ (.I(net81),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1764_ (.A1(net79),
    .A2(net80),
    .A3(_1350_),
    .A4(_1362_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1765_ (.A1(_1249_),
    .A2(_1318_),
    .A3(_1335_),
    .A4(_1367_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1766_ (.A1(_1366_),
    .A2(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1767_ (.A1(_1328_),
    .A2(_1369_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1768_ (.I(_1127_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1769_ (.A1(net71),
    .A2(_1281_),
    .A3(_1283_),
    .A4(_1325_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1770_ (.A1(net82),
    .A2(_1371_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1771_ (.A1(_1370_),
    .A2(_1372_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1772_ (.I(\prev_event_inc[5] ),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1773_ (.A1(net6),
    .A2(net12),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1774_ (.A1(_1373_),
    .A2(_1374_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1775_ (.A1(net83),
    .A2(_1375_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1776_ (.A1(_1370_),
    .A2(_1376_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1777_ (.I0(net84),
    .I1(_1451_),
    .S(_1375_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1778_ (.A1(_1370_),
    .A2(_1377_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1779_ (.A1(_1450_),
    .A2(_1375_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1780_ (.A1(net85),
    .A2(_1378_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1781_ (.A1(_1370_),
    .A2(_1379_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1782_ (.A1(net83),
    .A2(net84),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1783_ (.A1(_1373_),
    .A2(net85),
    .A3(_1374_),
    .A4(_1380_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1784_ (.I(_1381_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1785_ (.A1(net86),
    .A2(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1786_ (.A1(_1370_),
    .A2(_1383_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1787_ (.A1(_1373_),
    .A2(net85),
    .A3(_1450_),
    .A4(_1374_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1788_ (.I(_1384_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1789_ (.A1(net86),
    .A2(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1790_ (.A1(net87),
    .A2(_1386_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1791_ (.A1(_1370_),
    .A2(_1387_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1792_ (.A1(net86),
    .A2(net87),
    .A3(_1382_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1793_ (.A1(net88),
    .A2(_1388_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1794_ (.A1(_1370_),
    .A2(_1389_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1795_ (.A1(net86),
    .A2(net87),
    .A3(net88),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1796_ (.A1(_1385_),
    .A2(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1797_ (.A1(net89),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1798_ (.A1(_1370_),
    .A2(_1392_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1799_ (.A1(net89),
    .A2(_1390_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1800_ (.A1(_1382_),
    .A2(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1801_ (.A1(net90),
    .A2(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1802_ (.A1(_1370_),
    .A2(_1395_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1803_ (.A1(net90),
    .A2(_1385_),
    .A3(_1393_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1804_ (.A1(net91),
    .A2(_1396_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1805_ (.A1(_1370_),
    .A2(_1397_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1806_ (.I(_1127_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1807_ (.A1(net90),
    .A2(net91),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1808_ (.A1(_1382_),
    .A2(_1393_),
    .A3(_1399_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1809_ (.A1(net92),
    .A2(_1400_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1810_ (.A1(_1398_),
    .A2(_1401_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1811_ (.A1(net49),
    .A2(net60),
    .A3(net71),
    .A4(net82),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1812_ (.A1(_1167_),
    .A2(_1170_),
    .A3(_1240_),
    .A4(_1402_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1813_ (.A1(net93),
    .A2(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1814_ (.A1(_1398_),
    .A2(_1404_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1815_ (.A1(net92),
    .A2(_1385_),
    .A3(_1393_),
    .A4(_1399_),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1816_ (.A1(net94),
    .A2(_1405_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1817_ (.A1(_1398_),
    .A2(_1406_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1818_ (.A1(net90),
    .A2(net91),
    .A3(net92),
    .A4(net94),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1819_ (.A1(_1382_),
    .A2(_1393_),
    .A3(_1407_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1820_ (.A1(net95),
    .A2(_1408_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1821_ (.A1(_1398_),
    .A2(_1409_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1822_ (.A1(net95),
    .A2(_1385_),
    .A3(_1393_),
    .A4(_1407_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1823_ (.A1(net96),
    .A2(_1410_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1824_ (.A1(_1398_),
    .A2(_1411_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1825_ (.A1(net95),
    .A2(net96),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1826_ (.A1(_1382_),
    .A2(_1393_),
    .A3(_1407_),
    .A4(_1412_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1827_ (.A1(net97),
    .A2(_1413_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1828_ (.A1(_1398_),
    .A2(_1414_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1829_ (.A1(net95),
    .A2(net96),
    .A3(net97),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1830_ (.A1(net89),
    .A2(_1390_),
    .A3(_1407_),
    .A4(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1831_ (.A1(_1385_),
    .A2(_1416_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1832_ (.A1(net98),
    .A2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1833_ (.A1(_1398_),
    .A2(_1418_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1834_ (.A1(net98),
    .A2(_1415_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1835_ (.A1(_1382_),
    .A2(_1393_),
    .A3(_1407_),
    .A4(_1419_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1836_ (.A1(net99),
    .A2(_1420_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1837_ (.A1(_1398_),
    .A2(_1421_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1838_ (.A1(net98),
    .A2(net99),
    .A3(_1384_),
    .A4(_1416_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1839_ (.A1(net100),
    .A2(_1422_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1840_ (.A1(_1398_),
    .A2(_1423_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1841_ (.A1(net98),
    .A2(net99),
    .A3(net100),
    .A4(_1415_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1842_ (.A1(_1382_),
    .A2(_1393_),
    .A3(_1407_),
    .A4(_1424_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1843_ (.A1(net101),
    .A2(_1425_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1844_ (.A1(_1398_),
    .A2(_1426_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1845_ (.I(_1127_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1846_ (.A1(net98),
    .A2(net99),
    .A3(net100),
    .A4(net101),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1847_ (.A1(_1385_),
    .A2(_1416_),
    .A3(_1428_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1848_ (.A1(net102),
    .A2(_1429_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1849_ (.A1(_1427_),
    .A2(_1430_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1850_ (.A1(net102),
    .A2(_1415_),
    .A3(_1428_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1851_ (.A1(_1382_),
    .A2(_1393_),
    .A3(_1407_),
    .A4(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1852_ (.A1(net103),
    .A2(_1432_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1853_ (.A1(_1427_),
    .A2(_1433_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1854_ (.A1(net93),
    .A2(_1402_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1855_ (.A1(_1281_),
    .A2(_1283_),
    .A3(_1434_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1856_ (.A1(net104),
    .A2(_1435_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1857_ (.A1(_1427_),
    .A2(_1436_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1858_ (.A1(_1373_),
    .A2(net85),
    .A3(_1374_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1859_ (.A1(net102),
    .A2(_1428_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1860_ (.A1(net89),
    .A2(net103),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1861_ (.A1(_1390_),
    .A2(_1407_),
    .A3(_1415_),
    .A4(_1439_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1862_ (.A1(_1450_),
    .A2(_1437_),
    .A3(_1438_),
    .A4(_1440_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1863_ (.A1(net105),
    .A2(_1441_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1864_ (.A1(_1427_),
    .A2(_0264_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1865_ (.I(_1440_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1866_ (.A1(net105),
    .A2(_1380_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1867_ (.A1(_1437_),
    .A2(_1438_),
    .A3(_0265_),
    .A4(_0266_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1868_ (.A1(net106),
    .A2(_0267_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1869_ (.A1(_1427_),
    .A2(_0268_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1870_ (.A1(net105),
    .A2(net106),
    .A3(_1450_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1871_ (.A1(_1437_),
    .A2(_1438_),
    .A3(_0265_),
    .A4(_0269_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1872_ (.A1(net107),
    .A2(_0270_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1873_ (.A1(_1427_),
    .A2(_0271_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1874_ (.A1(net102),
    .A2(net105),
    .A3(net106),
    .A4(net107),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1875_ (.A1(_1428_),
    .A2(_0272_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1876_ (.A1(_1382_),
    .A2(_0265_),
    .A3(_0273_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1877_ (.A1(net108),
    .A2(_0274_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1878_ (.A1(_1427_),
    .A2(_0275_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1879_ (.A1(net108),
    .A2(_1384_),
    .A3(_1440_),
    .A4(_0273_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1880_ (.A1(net109),
    .A2(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1881_ (.A1(_1427_),
    .A2(_0277_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1882_ (.A1(net108),
    .A2(net109),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1883_ (.A1(_1381_),
    .A2(_0265_),
    .A3(_0273_),
    .A4(_0278_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1884_ (.A1(net110),
    .A2(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1885_ (.A1(_1427_),
    .A2(_0280_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1886_ (.A1(net110),
    .A2(_0278_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1887_ (.A1(_1385_),
    .A2(_0265_),
    .A3(_0273_),
    .A4(_0281_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1888_ (.A1(net111),
    .A2(_0282_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1889_ (.A1(_1427_),
    .A2(_0283_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1890_ (.I(_1126_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1891_ (.I(_0284_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1892_ (.A1(net108),
    .A2(net109),
    .A3(net110),
    .A4(net111),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1893_ (.A1(_1381_),
    .A2(_0265_),
    .A3(_0273_),
    .A4(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1894_ (.A1(net112),
    .A2(_0287_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1895_ (.A1(_0285_),
    .A2(_0288_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1896_ (.A1(net112),
    .A2(_0286_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1897_ (.A1(_1385_),
    .A2(_0265_),
    .A3(_0273_),
    .A4(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1898_ (.A1(net113),
    .A2(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1899_ (.A1(_0285_),
    .A2(_0291_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1900_ (.A1(net112),
    .A2(net113),
    .A3(_0286_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1901_ (.A1(_1381_),
    .A2(_0265_),
    .A3(_0273_),
    .A4(_0292_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1902_ (.A1(net114),
    .A2(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1903_ (.A1(_0285_),
    .A2(_0294_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1904_ (.A1(net93),
    .A2(net104),
    .A3(_1402_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1905_ (.A1(_1167_),
    .A2(_1170_),
    .A3(_1240_),
    .A4(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1906_ (.A1(net115),
    .A2(_0296_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1907_ (.A1(_0285_),
    .A2(_0297_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1908_ (.A1(net112),
    .A2(net113),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1909_ (.A1(net114),
    .A2(_0286_),
    .A3(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1910_ (.A1(_1385_),
    .A2(_0265_),
    .A3(_0273_),
    .A4(_0299_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1911_ (.A1(net116),
    .A2(_0300_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1912_ (.A1(_0285_),
    .A2(_0301_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1913_ (.A1(net114),
    .A2(net116),
    .A3(_0286_),
    .A4(_0298_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1914_ (.A1(_1381_),
    .A2(_0265_),
    .A3(_0273_),
    .A4(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1915_ (.A1(net117),
    .A2(_0303_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1916_ (.A1(_0285_),
    .A2(_0304_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1917_ (.I(\prev_event_inc[6] ),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1918_ (.A1(net6),
    .A2(net13),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1919_ (.A1(_0305_),
    .A2(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1920_ (.A1(net118),
    .A2(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1921_ (.A1(_0285_),
    .A2(_0308_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1922_ (.I0(net119),
    .I1(_1449_),
    .S(_0307_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1923_ (.A1(_0285_),
    .A2(_0309_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1924_ (.A1(_1448_),
    .A2(_0307_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1925_ (.A1(net120),
    .A2(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1926_ (.A1(_0285_),
    .A2(_0311_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1927_ (.A1(net118),
    .A2(net119),
    .A3(net120),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1928_ (.A1(_0305_),
    .A2(_0306_),
    .A3(_0312_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1929_ (.A1(net121),
    .A2(_0313_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1930_ (.A1(_0285_),
    .A2(_0314_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1931_ (.I(_0284_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1932_ (.A1(_0305_),
    .A2(net120),
    .A3(_1448_),
    .A4(_0306_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1933_ (.I(_0316_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1934_ (.A1(net121),
    .A2(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1935_ (.A1(net122),
    .A2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1936_ (.A1(_0315_),
    .A2(_0319_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _1937_ (.A1(net121),
    .A2(net122),
    .A3(_0313_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1938_ (.A1(net123),
    .A2(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _1939_ (.A1(_1143_),
    .A2(_0321_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1940_ (.A1(net121),
    .A2(net122),
    .A3(net123),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1941_ (.A1(_0317_),
    .A2(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1942_ (.A1(net124),
    .A2(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1943_ (.A1(_0315_),
    .A2(_0324_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1944_ (.A1(net121),
    .A2(net122),
    .A3(net123),
    .A4(net124),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1945_ (.A1(_0305_),
    .A2(_0306_),
    .A3(_0312_),
    .A4(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1946_ (.A1(net125),
    .A2(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1947_ (.A1(_0315_),
    .A2(_0327_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1948_ (.A1(net115),
    .A2(_1281_),
    .A3(_1283_),
    .A4(_0295_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1949_ (.A1(net126),
    .A2(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1950_ (.A1(_0315_),
    .A2(_0329_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1951_ (.I0(net127),
    .I1(_1445_),
    .S(_1131_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1952_ (.A1(_0315_),
    .A2(_0330_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1953_ (.A1(net125),
    .A2(_0317_),
    .A3(_0325_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1954_ (.A1(net128),
    .A2(_0331_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1955_ (.A1(_0315_),
    .A2(_0332_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1956_ (.A1(net125),
    .A2(net128),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1957_ (.A1(_0326_),
    .A2(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1958_ (.A1(net129),
    .A2(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1959_ (.A1(_0315_),
    .A2(_0335_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1960_ (.A1(net129),
    .A2(_0316_),
    .A3(_0325_),
    .A4(_0333_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1961_ (.A1(net130),
    .A2(_0336_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1962_ (.A1(_0315_),
    .A2(_0337_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1963_ (.A1(net125),
    .A2(net128),
    .A3(net129),
    .A4(net130),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1964_ (.A1(_0326_),
    .A2(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1965_ (.A1(net131),
    .A2(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1966_ (.A1(_0315_),
    .A2(_0340_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1967_ (.A1(net131),
    .A2(_0316_),
    .A3(_0325_),
    .A4(_0338_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1968_ (.A1(net132),
    .A2(_0341_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1969_ (.A1(_0315_),
    .A2(_0342_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1970_ (.I(_0284_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1971_ (.A1(net131),
    .A2(net132),
    .A3(_0326_),
    .A4(_0338_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1972_ (.A1(net133),
    .A2(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1973_ (.A1(_0343_),
    .A2(_0345_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1974_ (.A1(net124),
    .A2(net131),
    .A3(net132),
    .A4(net133),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1975_ (.A1(_0338_),
    .A2(_0346_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1976_ (.A1(_0317_),
    .A2(_0322_),
    .A3(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1977_ (.A1(net134),
    .A2(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1978_ (.A1(_0343_),
    .A2(_0349_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1979_ (.A1(net131),
    .A2(net132),
    .A3(net133),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1980_ (.A1(net134),
    .A2(_0326_),
    .A3(_0338_),
    .A4(_0350_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1981_ (.A1(net135),
    .A2(_0351_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1982_ (.A1(_0343_),
    .A2(_0352_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1983_ (.A1(net134),
    .A2(net135),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1984_ (.A1(_0317_),
    .A2(_0322_),
    .A3(_0347_),
    .A4(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1985_ (.A1(net136),
    .A2(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1986_ (.A1(_0343_),
    .A2(_0355_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1987_ (.A1(net136),
    .A2(_0353_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1988_ (.A1(_0326_),
    .A2(_0338_),
    .A3(_0350_),
    .A4(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1989_ (.A1(net137),
    .A2(_0357_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1990_ (.A1(_0343_),
    .A2(_0358_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1991_ (.A1(net93),
    .A2(net104),
    .A3(net115),
    .A4(net126),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1992_ (.A1(_1402_),
    .A2(_0359_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1993_ (.A1(_1167_),
    .A2(_1170_),
    .A3(_1240_),
    .A4(_0360_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1994_ (.A1(net138),
    .A2(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1995_ (.A1(_0343_),
    .A2(_0362_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1996_ (.A1(net134),
    .A2(net135),
    .A3(net136),
    .A4(net137),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1997_ (.A1(_0317_),
    .A2(_0322_),
    .A3(_0347_),
    .A4(_0363_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1998_ (.A1(net139),
    .A2(_0364_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1999_ (.A1(_0343_),
    .A2(_0365_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2000_ (.A1(net139),
    .A2(_0363_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2001_ (.A1(_0326_),
    .A2(_0338_),
    .A3(_0350_),
    .A4(_0366_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2002_ (.A1(net140),
    .A2(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2003_ (.A1(_0343_),
    .A2(_0368_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 _2004_ (.I(_0366_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2005_ (.A1(net140),
    .A2(_0322_),
    .A3(_0338_),
    .A4(_0346_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2006_ (.A1(_0317_),
    .A2(_0369_),
    .A3(_0370_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2007_ (.A1(net141),
    .A2(_0371_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2008_ (.A1(_0343_),
    .A2(_0372_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2009_ (.A1(net141),
    .A2(_0313_),
    .A3(_0369_),
    .A4(_0370_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2010_ (.A1(net142),
    .A2(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2011_ (.A1(_0343_),
    .A2(_0374_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _2012_ (.I(_0284_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2013_ (.A1(net141),
    .A2(net142),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2014_ (.A1(_0317_),
    .A2(_0369_),
    .A3(_0370_),
    .A4(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2015_ (.A1(net143),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2016_ (.A1(_0375_),
    .A2(_0378_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2017_ (.A1(net140),
    .A2(net141),
    .A3(net142),
    .A4(net143),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2018_ (.A1(_0322_),
    .A2(_0338_),
    .A3(_0346_),
    .A4(_0379_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2019_ (.A1(_0313_),
    .A2(_0369_),
    .A3(_0380_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2020_ (.A1(net144),
    .A2(_0381_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2021_ (.A1(_0375_),
    .A2(_0382_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2022_ (.A1(net144),
    .A2(_0316_),
    .A3(_0366_),
    .A4(_0380_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2023_ (.A1(net145),
    .A2(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2024_ (.A1(_0375_),
    .A2(_0384_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2025_ (.A1(net144),
    .A2(net145),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2026_ (.A1(_0313_),
    .A2(_0369_),
    .A3(_0380_),
    .A4(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2027_ (.A1(net146),
    .A2(_0386_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2028_ (.A1(_0375_),
    .A2(_0387_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2029_ (.A1(net146),
    .A2(_0385_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2030_ (.A1(_0317_),
    .A2(_0369_),
    .A3(_0380_),
    .A4(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2031_ (.A1(net147),
    .A2(_0389_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2032_ (.A1(_0375_),
    .A2(_0390_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2033_ (.A1(net144),
    .A2(net145),
    .A3(net146),
    .A4(net147),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2034_ (.A1(_0313_),
    .A2(_0369_),
    .A3(_0380_),
    .A4(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2035_ (.A1(net148),
    .A2(_0392_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2036_ (.A1(_0375_),
    .A2(_0393_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2037_ (.A1(net138),
    .A2(_1281_),
    .A3(_1283_),
    .A4(_0360_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2038_ (.A1(net149),
    .A2(_0394_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2039_ (.A1(_0375_),
    .A2(_0395_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2040_ (.A1(net148),
    .A2(_0391_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2041_ (.A1(_0317_),
    .A2(_0369_),
    .A3(_0380_),
    .A4(_0396_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2042_ (.A1(net150),
    .A2(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2043_ (.A1(_0375_),
    .A2(_0398_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2044_ (.A1(net148),
    .A2(net150),
    .A3(_0391_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2045_ (.A1(_0313_),
    .A2(_0369_),
    .A3(_0380_),
    .A4(_0399_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2046_ (.A1(net151),
    .A2(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2047_ (.A1(_0375_),
    .A2(_0401_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2048_ (.A1(net148),
    .A2(net150),
    .A3(net151),
    .A4(_0391_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2049_ (.A1(_0316_),
    .A2(_0369_),
    .A3(_0380_),
    .A4(_0402_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2050_ (.A1(net152),
    .A2(_0403_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2051_ (.A1(_0375_),
    .A2(_0404_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2052_ (.A1(_1200_),
    .A2(net153),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2053_ (.A1(_1126_),
    .A2(net153),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2054_ (.A1(net152),
    .A2(_0381_),
    .A3(_0402_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2055_ (.I0(_0405_),
    .I1(_0406_),
    .S(_0407_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _2056_ (.I(_0284_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2057_ (.I(net154),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2058_ (.I(\prev_event_inc[7] ),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2059_ (.A1(_1133_),
    .A2(net14),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2060_ (.A1(_0410_),
    .A2(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2061_ (.A1(_0409_),
    .A2(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2062_ (.A1(_0408_),
    .A2(_0413_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2063_ (.I0(net155),
    .I1(_1447_),
    .S(_0412_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2064_ (.A1(_0408_),
    .A2(_0414_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2065_ (.I(net156),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2066_ (.A1(_0410_),
    .A2(_1446_),
    .A3(_0411_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2067_ (.A1(_0415_),
    .A2(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2068_ (.A1(_0408_),
    .A2(_0417_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2069_ (.I(net157),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2070_ (.A1(net154),
    .A2(net155),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2071_ (.A1(_0410_),
    .A2(_0411_),
    .A3(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2072_ (.A1(net156),
    .A2(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2073_ (.A1(_0418_),
    .A2(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2074_ (.A1(_0408_),
    .A2(_0422_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2075_ (.I(net158),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2076_ (.A1(net156),
    .A2(net157),
    .A3(_0416_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2077_ (.A1(_0423_),
    .A2(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2078_ (.A1(_0408_),
    .A2(_0425_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2079_ (.I(net159),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2080_ (.A1(net156),
    .A2(net157),
    .A3(net158),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2081_ (.A1(_0420_),
    .A2(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2082_ (.A1(_0426_),
    .A2(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2083_ (.A1(_0408_),
    .A2(_0429_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2084_ (.A1(net138),
    .A2(net149),
    .A3(_1402_),
    .A4(_0359_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2085_ (.A1(_1167_),
    .A2(_1170_),
    .A3(_1240_),
    .A4(_0430_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2086_ (.A1(net160),
    .A2(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2087_ (.A1(_0408_),
    .A2(_0432_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2088_ (.I(net161),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2089_ (.A1(_0410_),
    .A2(_1446_),
    .A3(_0411_),
    .A4(_0427_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2090_ (.A1(net159),
    .A2(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2091_ (.A1(_0433_),
    .A2(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2092_ (.A1(_0408_),
    .A2(_0436_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2093_ (.I(net162),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2094_ (.A1(net159),
    .A2(net161),
    .A3(_0420_),
    .A4(_0427_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2095_ (.A1(_0437_),
    .A2(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2096_ (.A1(_0408_),
    .A2(_0439_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2097_ (.I(net163),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2098_ (.A1(net159),
    .A2(net161),
    .A3(net162),
    .A4(_0434_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2099_ (.A1(_0440_),
    .A2(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2100_ (.A1(_0408_),
    .A2(_0442_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _2101_ (.I(_0284_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2102_ (.I(net164),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2103_ (.A1(net159),
    .A2(net161),
    .A3(net162),
    .A4(net163),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2104_ (.A1(_0420_),
    .A2(_0427_),
    .A3(_0445_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2105_ (.A1(_0444_),
    .A2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2106_ (.A1(_0443_),
    .A2(_0447_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2107_ (.I(net165),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2108_ (.A1(net164),
    .A2(_0434_),
    .A3(_0445_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2109_ (.A1(_0448_),
    .A2(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2110_ (.A1(_0443_),
    .A2(_0450_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2111_ (.I(net166),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2112_ (.A1(net164),
    .A2(net165),
    .A3(_0445_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2113_ (.A1(_0420_),
    .A2(_0427_),
    .A3(_0452_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2114_ (.A1(_0451_),
    .A2(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2115_ (.A1(_0443_),
    .A2(_0454_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2116_ (.I(net167),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2117_ (.A1(net166),
    .A2(_0434_),
    .A3(_0452_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2118_ (.A1(_0455_),
    .A2(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2119_ (.A1(_0443_),
    .A2(_0457_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2120_ (.I(net168),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2121_ (.A1(net166),
    .A2(net167),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2122_ (.A1(_0427_),
    .A2(_0459_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2123_ (.A1(_0420_),
    .A2(_0452_),
    .A3(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2124_ (.A1(_0458_),
    .A2(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2125_ (.A1(_0443_),
    .A2(_0462_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2126_ (.I(net169),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2127_ (.A1(net168),
    .A2(_0416_),
    .A3(_0452_),
    .A4(_0460_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2128_ (.A1(_0463_),
    .A2(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2129_ (.A1(_0443_),
    .A2(_0465_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2130_ (.I(net170),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2131_ (.A1(net164),
    .A2(_0427_),
    .A3(_0445_),
    .A4(_0459_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2132_ (.A1(net165),
    .A2(net168),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2133_ (.A1(net169),
    .A2(_0420_),
    .A3(_0467_),
    .A4(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2134_ (.A1(_0466_),
    .A2(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2135_ (.A1(_0443_),
    .A2(_0470_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2136_ (.A1(net160),
    .A2(_1281_),
    .A3(_1283_),
    .A4(_0430_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2137_ (.A1(net171),
    .A2(_0471_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2138_ (.A1(_0443_),
    .A2(_0472_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2139_ (.I(net172),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2140_ (.A1(net165),
    .A2(net168),
    .A3(net169),
    .A4(net170),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2141_ (.A1(_0410_),
    .A2(_1446_),
    .A3(_0411_),
    .A4(_0474_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2142_ (.A1(_0467_),
    .A2(_0475_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2143_ (.A1(_0473_),
    .A2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2144_ (.A1(_0443_),
    .A2(_0477_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2145_ (.I(net173),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2146_ (.A1(_0410_),
    .A2(_0411_),
    .A3(_0419_),
    .A4(_0474_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2147_ (.A1(net172),
    .A2(_0467_),
    .A3(_0479_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2148_ (.A1(_0478_),
    .A2(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2149_ (.A1(_0443_),
    .A2(_0481_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _2150_ (.I(_0284_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2151_ (.I(net174),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2152_ (.A1(net172),
    .A2(net173),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2153_ (.A1(_0467_),
    .A2(_0475_),
    .A3(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2154_ (.A1(_0483_),
    .A2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2155_ (.A1(_0482_),
    .A2(_0486_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2156_ (.I(net175),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2157_ (.A1(net174),
    .A2(_0467_),
    .A3(_0479_),
    .A4(_0484_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2158_ (.A1(_0487_),
    .A2(_0488_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2159_ (.A1(_0482_),
    .A2(_0489_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2160_ (.I(net176),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2161_ (.A1(net172),
    .A2(net173),
    .A3(net174),
    .A4(net175),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2162_ (.A1(_0467_),
    .A2(_0475_),
    .A3(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2163_ (.A1(_0490_),
    .A2(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2164_ (.A1(_0482_),
    .A2(_0493_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2165_ (.I(net177),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2166_ (.A1(net164),
    .A2(net166),
    .A3(net167),
    .A4(net176),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2167_ (.A1(_0427_),
    .A2(_0445_),
    .A3(_0491_),
    .A4(_0495_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _2168_ (.I(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2169_ (.A1(_0479_),
    .A2(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2170_ (.A1(_0494_),
    .A2(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2171_ (.A1(_0482_),
    .A2(_0499_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2172_ (.I(net178),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2173_ (.A1(net177),
    .A2(_0475_),
    .A3(_0497_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2174_ (.A1(_0500_),
    .A2(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2175_ (.A1(_0482_),
    .A2(_0502_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2176_ (.I(net179),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2177_ (.A1(net177),
    .A2(net178),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2178_ (.A1(_0479_),
    .A2(_0497_),
    .A3(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2179_ (.A1(_0503_),
    .A2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2180_ (.A1(_0482_),
    .A2(_0506_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2181_ (.I(net180),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2182_ (.A1(net179),
    .A2(_0475_),
    .A3(_0497_),
    .A4(_0504_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2183_ (.A1(_0507_),
    .A2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2184_ (.A1(_0482_),
    .A2(_0509_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2185_ (.I(net181),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2186_ (.A1(net177),
    .A2(net178),
    .A3(net179),
    .A4(net180),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2187_ (.A1(_0479_),
    .A2(_0497_),
    .A3(_0511_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2188_ (.A1(_0510_),
    .A2(_0512_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2189_ (.A1(_0482_),
    .A2(_0513_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2190_ (.A1(net138),
    .A2(net149),
    .A3(net160),
    .A4(net171),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2191_ (.A1(_1402_),
    .A2(_0359_),
    .A3(_0514_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2192_ (.A1(_1166_),
    .A2(_1170_),
    .A3(_1240_),
    .A4(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2193_ (.A1(net182),
    .A2(_0516_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2194_ (.A1(_0482_),
    .A2(_0517_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2195_ (.I(net183),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2196_ (.A1(net181),
    .A2(_0511_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2197_ (.A1(_0475_),
    .A2(_0497_),
    .A3(_0519_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2198_ (.A1(_0518_),
    .A2(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2199_ (.A1(_0482_),
    .A2(_0521_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2200_ (.I(_0284_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2201_ (.I(net184),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2202_ (.A1(net183),
    .A2(_0479_),
    .A3(_0497_),
    .A4(_0519_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2203_ (.A1(_0523_),
    .A2(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2204_ (.A1(_0522_),
    .A2(_0525_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2205_ (.I(net185),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2206_ (.A1(net181),
    .A2(net183),
    .A3(net184),
    .A4(_0511_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2207_ (.A1(_0475_),
    .A2(_0497_),
    .A3(_0527_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2208_ (.A1(_0526_),
    .A2(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2209_ (.A1(_0522_),
    .A2(_0529_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2210_ (.I(net186),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2211_ (.A1(net185),
    .A2(_0479_),
    .A3(_0497_),
    .A4(_0527_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2212_ (.A1(_0530_),
    .A2(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2213_ (.A1(_0522_),
    .A2(_0532_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2214_ (.I(net187),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2215_ (.A1(net181),
    .A2(net183),
    .A3(net184),
    .A4(net185),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2216_ (.A1(net186),
    .A2(_0511_),
    .A3(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2217_ (.A1(_0475_),
    .A2(_0497_),
    .A3(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2218_ (.A1(_0533_),
    .A2(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2219_ (.A1(_0522_),
    .A2(_0537_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2220_ (.I(net188),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2221_ (.A1(net187),
    .A2(_0479_),
    .A3(_0496_),
    .A4(_0535_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2222_ (.A1(_0538_),
    .A2(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2223_ (.A1(_0522_),
    .A2(_0540_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2224_ (.A1(net182),
    .A2(_1281_),
    .A3(_1283_),
    .A4(_0515_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2225_ (.A1(net189),
    .A2(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2226_ (.A1(_0522_),
    .A2(_0542_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2227_ (.A1(net182),
    .A2(net189),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2228_ (.A1(_1402_),
    .A2(_0359_),
    .A3(_0514_),
    .A4(_0543_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2229_ (.A1(_1166_),
    .A2(_1169_),
    .A3(_1240_),
    .A4(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2230_ (.A1(net190),
    .A2(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2231_ (.A1(_0522_),
    .A2(_0546_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2232_ (.A1(_1281_),
    .A2(_1283_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2233_ (.A1(net190),
    .A2(_0544_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2234_ (.A1(_0547_),
    .A2(_0548_),
    .B(net191),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2235_ (.A1(net191),
    .A2(_0547_),
    .A3(_0548_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2236_ (.A1(_0549_),
    .A2(_0550_),
    .B(_1143_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2237_ (.A1(_1198_),
    .A2(net192),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2238_ (.A1(_1200_),
    .A2(net192),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2239_ (.A1(net190),
    .A2(net191),
    .A3(_0545_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2240_ (.I0(_0551_),
    .I1(_0552_),
    .S(_0553_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _2241_ (.A1(net190),
    .A2(net191),
    .A3(net192),
    .A4(_0544_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2242_ (.A1(_0547_),
    .A2(_0554_),
    .B(net193),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2243_ (.A1(net193),
    .A2(_0547_),
    .A3(_0554_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2244_ (.A1(_0555_),
    .A2(_0556_),
    .B(_1143_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2245_ (.A1(_1444_),
    .A2(_1131_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2246_ (.A1(net194),
    .A2(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2247_ (.A1(_0522_),
    .A2(_0558_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2248_ (.A1(net193),
    .A2(_1167_),
    .A3(_1170_),
    .A4(_1240_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2249_ (.A1(_0554_),
    .A2(_0559_),
    .B(net195),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2250_ (.A1(net195),
    .A2(_0554_),
    .A3(_0559_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2251_ (.A1(_0560_),
    .A2(_0561_),
    .B(_1143_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2252_ (.A1(net193),
    .A2(net195),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2253_ (.A1(_0547_),
    .A2(_0554_),
    .A3(_0562_),
    .B(net196),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _2254_ (.A1(net196),
    .A2(_0547_),
    .A3(_0554_),
    .A4(_0562_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2255_ (.A1(_0563_),
    .A2(_0564_),
    .B(_1143_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2256_ (.I(\prev_event_inc[1] ),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2257_ (.A1(_1133_),
    .A2(net8),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2258_ (.A1(_0565_),
    .A2(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2259_ (.A1(net197),
    .A2(_0567_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2260_ (.A1(_0522_),
    .A2(_0568_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2261_ (.I0(net198),
    .I1(_1443_),
    .S(_0567_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2262_ (.A1(_0522_),
    .A2(_0569_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _2263_ (.I(_0284_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2264_ (.A1(_1442_),
    .A2(_0567_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2265_ (.A1(net199),
    .A2(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2266_ (.A1(_0570_),
    .A2(_0572_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2267_ (.A1(net197),
    .A2(net199),
    .A3(net198),
    .A4(_0567_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2268_ (.A1(net200),
    .A2(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2269_ (.A1(_0570_),
    .A2(_0574_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _2270_ (.I(net201),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2271_ (.A1(net199),
    .A2(net200),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _2272_ (.A1(_0565_),
    .A2(_1442_),
    .A3(_0566_),
    .A4(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2273_ (.A1(_0575_),
    .A2(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2274_ (.A1(_0570_),
    .A2(_0578_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2275_ (.A1(net197),
    .A2(net199),
    .A3(net198),
    .A4(net200),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2276_ (.A1(_0565_),
    .A2(net201),
    .A3(_0566_),
    .A4(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2277_ (.I(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2278_ (.A1(net202),
    .A2(_0581_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2279_ (.A1(_0570_),
    .A2(_0582_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2280_ (.A1(_0575_),
    .A2(net202),
    .A3(_0577_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2281_ (.A1(net203),
    .A2(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2282_ (.A1(_0570_),
    .A2(_0584_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2283_ (.A1(net202),
    .A2(net203),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2284_ (.A1(_0581_),
    .A2(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2285_ (.A1(net204),
    .A2(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2286_ (.A1(_0570_),
    .A2(_0587_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2287_ (.A1(net205),
    .A2(_1205_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2288_ (.A1(_0570_),
    .A2(_0588_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2289_ (.A1(_0575_),
    .A2(net204),
    .A3(_0577_),
    .A4(_0585_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2290_ (.A1(net206),
    .A2(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2291_ (.A1(_0570_),
    .A2(_0590_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2292_ (.A1(net202),
    .A2(net203),
    .A3(net204),
    .A4(net206),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2293_ (.A1(_0581_),
    .A2(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2294_ (.A1(net207),
    .A2(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2295_ (.A1(_0570_),
    .A2(_0593_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2296_ (.A1(_0575_),
    .A2(net207),
    .A3(_0577_),
    .A4(_0591_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2297_ (.A1(net208),
    .A2(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2298_ (.A1(_0570_),
    .A2(_0595_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _2299_ (.I(_0284_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2300_ (.A1(net207),
    .A2(net208),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2301_ (.A1(_0591_),
    .A2(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2302_ (.A1(_0581_),
    .A2(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2303_ (.A1(net209),
    .A2(_0599_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2304_ (.A1(_0596_),
    .A2(_0600_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2305_ (.A1(_0575_),
    .A2(net209),
    .A3(_0577_),
    .A4(_0598_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2306_ (.A1(net210),
    .A2(_0601_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2307_ (.A1(_0596_),
    .A2(_0602_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2308_ (.A1(net209),
    .A2(net210),
    .A3(_0580_),
    .A4(_0598_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2309_ (.A1(net211),
    .A2(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2310_ (.A1(_0596_),
    .A2(_0604_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2311_ (.A1(net209),
    .A2(net210),
    .A3(net211),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2312_ (.A1(_0575_),
    .A2(_0577_),
    .A3(_0598_),
    .A4(_0605_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2313_ (.A1(net212),
    .A2(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2314_ (.A1(_0596_),
    .A2(_0607_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2315_ (.A1(net209),
    .A2(net210),
    .A3(net211),
    .A4(net212),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2316_ (.A1(_0581_),
    .A2(_0598_),
    .A3(_0608_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2317_ (.A1(net213),
    .A2(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2318_ (.A1(_0596_),
    .A2(_0610_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2319_ (.A1(net213),
    .A2(_0608_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2320_ (.A1(_0575_),
    .A2(_0577_),
    .A3(_0598_),
    .A4(_0611_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2321_ (.A1(net214),
    .A2(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2322_ (.A1(_0596_),
    .A2(_0613_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2323_ (.A1(net213),
    .A2(net214),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2324_ (.A1(_0591_),
    .A2(_0597_),
    .A3(_0608_),
    .A4(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2325_ (.I(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2326_ (.A1(_0581_),
    .A2(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2327_ (.A1(net215),
    .A2(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2328_ (.A1(_0596_),
    .A2(_0618_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2329_ (.A1(net205),
    .A2(_1167_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2330_ (.A1(net216),
    .A2(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2331_ (.A1(_0596_),
    .A2(_0620_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2332_ (.A1(_0575_),
    .A2(net215),
    .A3(_0577_),
    .A4(_0615_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2333_ (.A1(net217),
    .A2(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2334_ (.A1(_0596_),
    .A2(_0622_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2335_ (.A1(net215),
    .A2(net217),
    .A3(_0580_),
    .A4(_0615_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2336_ (.A1(net218),
    .A2(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2337_ (.A1(_0596_),
    .A2(_0624_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2338_ (.A1(_1198_),
    .A2(net219),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2339_ (.A1(_1200_),
    .A2(net219),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2340_ (.A1(_0575_),
    .A2(_0577_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2341_ (.A1(net215),
    .A2(net217),
    .A3(net218),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2342_ (.A1(_0627_),
    .A2(_0616_),
    .A3(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2343_ (.I0(_0625_),
    .I1(_0626_),
    .S(_0629_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _2344_ (.I(_1198_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2345_ (.A1(net219),
    .A2(_0628_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2346_ (.A1(_0581_),
    .A2(_0616_),
    .A3(_0631_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2347_ (.A1(net220),
    .A2(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2348_ (.A1(_0630_),
    .A2(_0633_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2349_ (.A1(_1198_),
    .A2(net221),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2350_ (.A1(_1200_),
    .A2(net221),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2351_ (.A1(net201),
    .A2(_0577_),
    .A3(_0631_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2352_ (.A1(net220),
    .A2(_0616_),
    .A3(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2353_ (.I0(_0634_),
    .I1(_0635_),
    .S(_0637_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2354_ (.A1(net220),
    .A2(net221),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2355_ (.A1(_0581_),
    .A2(_0616_),
    .A3(_0631_),
    .A4(_0638_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2356_ (.A1(net222),
    .A2(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2357_ (.A1(_0630_),
    .A2(_0640_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2358_ (.A1(_1126_),
    .A2(net223),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2359_ (.A1(_1200_),
    .A2(net223),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2360_ (.A1(net222),
    .A2(_0616_),
    .A3(_0636_),
    .A4(_0638_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2361_ (.I0(_0641_),
    .I1(_0642_),
    .S(_0643_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2362_ (.A1(net220),
    .A2(net221),
    .A3(net222),
    .A4(net223),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2363_ (.A1(_0581_),
    .A2(_0616_),
    .A3(_0631_),
    .A4(_0644_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2364_ (.A1(net224),
    .A2(_0645_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2365_ (.A1(_0630_),
    .A2(_0646_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2366_ (.A1(_1126_),
    .A2(net225),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2367_ (.A1(net1),
    .A2(net225),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2368_ (.A1(net224),
    .A2(_0616_),
    .A3(_0636_),
    .A4(_0644_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2369_ (.I0(_0647_),
    .I1(_0648_),
    .S(_0649_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2370_ (.A1(net224),
    .A2(net225),
    .A3(_0644_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2371_ (.A1(_0581_),
    .A2(_0615_),
    .A3(_0631_),
    .A4(_0650_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2372_ (.A1(net226),
    .A2(_0651_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2373_ (.A1(_0630_),
    .A2(_0652_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2374_ (.A1(net205),
    .A2(net216),
    .A3(_1205_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2375_ (.A1(net227),
    .A2(_0653_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2376_ (.A1(_0630_),
    .A2(_0654_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2377_ (.A1(_1126_),
    .A2(net228),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2378_ (.A1(net1),
    .A2(net228),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2379_ (.A1(net226),
    .A2(_0616_),
    .A3(_0636_),
    .A4(_0650_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2380_ (.I0(_0655_),
    .I1(_0656_),
    .S(_0657_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2381_ (.A1(net226),
    .A2(net228),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2382_ (.A1(net224),
    .A2(net225),
    .A3(_0644_),
    .A4(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2383_ (.A1(_0580_),
    .A2(_0615_),
    .A3(_0631_),
    .A4(_0659_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2384_ (.A1(net229),
    .A2(_0660_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2385_ (.A1(_0630_),
    .A2(_0661_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2386_ (.A1(_1126_),
    .A2(net230),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2387_ (.A1(net1),
    .A2(net230),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2388_ (.A1(net229),
    .A2(_0659_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2389_ (.A1(_0616_),
    .A2(_0636_),
    .A3(_0664_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2390_ (.I0(_0662_),
    .I1(_0663_),
    .S(_0665_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2391_ (.A1(net224),
    .A2(net225),
    .A3(net226),
    .A4(net228),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2392_ (.A1(net229),
    .A2(net230),
    .A3(_0644_),
    .A4(_0666_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2393_ (.A1(_0580_),
    .A2(_0615_),
    .A3(_0631_),
    .A4(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2394_ (.A1(net231),
    .A2(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2395_ (.A1(_0630_),
    .A2(_0669_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _2396_ (.I(net232),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2397_ (.I(\prev_event_inc[2] ),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2398_ (.A1(net9),
    .A2(_0671_),
    .A3(_1133_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2399_ (.A1(_0670_),
    .A2(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2400_ (.A1(_0630_),
    .A2(_0673_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2401_ (.I0(net233),
    .I1(_1457_),
    .S(_0672_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2402_ (.A1(_0630_),
    .A2(_0674_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2403_ (.I(net234),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2404_ (.A1(_1456_),
    .A2(_0672_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2405_ (.A1(_0675_),
    .A2(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2406_ (.A1(_0630_),
    .A2(_0677_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _2407_ (.I(_1198_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2408_ (.I(net235),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2409_ (.A1(net233),
    .A2(net232),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2410_ (.A1(net9),
    .A2(_0671_),
    .A3(_1133_),
    .A4(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2411_ (.A1(net234),
    .A2(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2412_ (.A1(_0679_),
    .A2(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2413_ (.A1(_0678_),
    .A2(_0683_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2414_ (.I(net236),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2415_ (.A1(net235),
    .A2(net234),
    .A3(_1456_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2416_ (.A1(net9),
    .A2(_0671_),
    .A3(_1133_),
    .A4(_0685_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2417_ (.A1(_0684_),
    .A2(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2418_ (.A1(_0678_),
    .A2(_0687_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2419_ (.I(net237),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2420_ (.A1(net235),
    .A2(net234),
    .A3(net233),
    .A4(net232),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2421_ (.A1(net9),
    .A2(_0671_),
    .A3(_1133_),
    .A4(_0689_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2422_ (.A1(net236),
    .A2(_0690_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2423_ (.A1(_0688_),
    .A2(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2424_ (.A1(_0678_),
    .A2(_0692_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2425_ (.A1(net205),
    .A2(net216),
    .A3(net227),
    .A4(_1166_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2426_ (.A1(net238),
    .A2(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2427_ (.A1(_0678_),
    .A2(_0694_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2428_ (.I(net239),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2429_ (.A1(net237),
    .A2(net236),
    .A3(_0686_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2430_ (.A1(_0695_),
    .A2(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2431_ (.A1(_0678_),
    .A2(_0697_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2432_ (.I(net240),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2433_ (.A1(net239),
    .A2(net237),
    .A3(net236),
    .A4(_0690_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2434_ (.A1(_0698_),
    .A2(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2435_ (.A1(_0678_),
    .A2(_0700_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2436_ (.I(net241),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2437_ (.A1(net240),
    .A2(net239),
    .A3(net237),
    .A4(net236),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2438_ (.A1(_0686_),
    .A2(_0702_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2439_ (.A1(_0701_),
    .A2(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2440_ (.A1(_0678_),
    .A2(_0704_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2441_ (.I(net242),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2442_ (.A1(net241),
    .A2(_0702_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2443_ (.A1(_0690_),
    .A2(_0706_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2444_ (.A1(_0705_),
    .A2(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2445_ (.A1(_0678_),
    .A2(_0708_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2446_ (.I(net243),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2447_ (.A1(net242),
    .A2(_0686_),
    .A3(_0706_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2448_ (.A1(_0709_),
    .A2(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2449_ (.A1(_0678_),
    .A2(_0711_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2450_ (.I(net244),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2451_ (.A1(net243),
    .A2(net242),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2452_ (.A1(_0690_),
    .A2(_0706_),
    .A3(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2453_ (.A1(_0712_),
    .A2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2454_ (.A1(_0678_),
    .A2(_0715_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _2455_ (.I(_1198_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2456_ (.I(net245),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2457_ (.A1(net244),
    .A2(_0686_),
    .A3(_0706_),
    .A4(_0713_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2458_ (.A1(_0717_),
    .A2(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2459_ (.A1(_0716_),
    .A2(_0719_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2460_ (.I(net246),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2461_ (.A1(net245),
    .A2(net244),
    .A3(net243),
    .A4(net242),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2462_ (.A1(_0690_),
    .A2(_0706_),
    .A3(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2463_ (.A1(_0720_),
    .A2(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2464_ (.A1(_0716_),
    .A2(_0723_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2465_ (.I(net247),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2466_ (.A1(net246),
    .A2(_0686_),
    .A3(_0706_),
    .A4(_0721_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2467_ (.A1(_0724_),
    .A2(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2468_ (.A1(_0716_),
    .A2(_0726_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2469_ (.I(net248),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2470_ (.A1(net247),
    .A2(net246),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2471_ (.A1(_0690_),
    .A2(_0706_),
    .A3(_0721_),
    .A4(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2472_ (.A1(_0727_),
    .A2(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2473_ (.A1(_0716_),
    .A2(_0730_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2474_ (.A1(_1168_),
    .A2(_1205_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2475_ (.A1(net249),
    .A2(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2476_ (.A1(_0716_),
    .A2(_0732_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2477_ (.I(net250),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2478_ (.A1(_1133_),
    .A2(_1456_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2479_ (.A1(net248),
    .A2(net235),
    .A3(net234),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2480_ (.A1(net9),
    .A2(_0671_),
    .A3(_0734_),
    .A4(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2481_ (.A1(net241),
    .A2(_0702_),
    .A3(_0721_),
    .A4(_0728_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2482_ (.I(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2483_ (.A1(_0736_),
    .A2(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2484_ (.A1(_0733_),
    .A2(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2485_ (.A1(_0716_),
    .A2(_0740_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2486_ (.I(net251),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2487_ (.A1(net250),
    .A2(net248),
    .A3(_0690_),
    .A4(_0738_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2488_ (.A1(_0741_),
    .A2(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2489_ (.A1(_0716_),
    .A2(_0743_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2490_ (.I(net252),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2491_ (.A1(net251),
    .A2(net250),
    .A3(_0736_),
    .A4(_0737_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2492_ (.A1(_0744_),
    .A2(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2493_ (.A1(_0716_),
    .A2(_0746_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2494_ (.I(net253),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2495_ (.A1(net252),
    .A2(net251),
    .A3(net250),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2496_ (.A1(net248),
    .A2(_0690_),
    .A3(_0738_),
    .A4(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2497_ (.A1(_0747_),
    .A2(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2498_ (.A1(_0716_),
    .A2(_0750_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2499_ (.I(net254),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2500_ (.A1(net253),
    .A2(net252),
    .A3(net251),
    .A4(net250),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2501_ (.A1(_0736_),
    .A2(_0738_),
    .A3(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2502_ (.A1(_0751_),
    .A2(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2503_ (.A1(_0716_),
    .A2(_0754_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2504_ (.I(_1198_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2505_ (.A1(net254),
    .A2(_0752_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _2506_ (.A1(_0681_),
    .A2(_0735_),
    .A3(_0738_),
    .A4(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2507_ (.A1(net255),
    .A2(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2508_ (.A1(_0755_),
    .A2(_0758_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2509_ (.I(net256),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2510_ (.A1(net255),
    .A2(_0736_),
    .A3(_0738_),
    .A4(_0756_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2511_ (.A1(_0759_),
    .A2(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2512_ (.A1(_0755_),
    .A2(_0761_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2513_ (.I(_0757_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2514_ (.A1(net256),
    .A2(net255),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2515_ (.A1(_0762_),
    .A2(_0763_),
    .B(net257),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2516_ (.A1(net257),
    .A2(_0762_),
    .A3(_0763_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2517_ (.A1(_0764_),
    .A2(_0765_),
    .B(_1143_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2518_ (.I(net258),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2519_ (.I(net257),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2520_ (.A1(_0767_),
    .A2(_0763_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2521_ (.A1(_0736_),
    .A2(_0738_),
    .A3(_0756_),
    .A4(_0768_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2522_ (.A1(_0766_),
    .A2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2523_ (.A1(_0755_),
    .A2(_0770_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2524_ (.A1(net258),
    .A2(_0768_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2525_ (.A1(_0762_),
    .A2(_0771_),
    .B(net259),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2526_ (.A1(net259),
    .A2(_0762_),
    .A3(_0771_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2527_ (.A1(_0772_),
    .A2(_0773_),
    .B(_1143_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2528_ (.A1(net249),
    .A2(_1167_),
    .A3(_1168_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2529_ (.A1(net260),
    .A2(_0774_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2530_ (.A1(_0755_),
    .A2(_0775_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2531_ (.I(net261),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2532_ (.A1(net257),
    .A2(net256),
    .A3(net255),
    .A4(net258),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2533_ (.A1(net259),
    .A2(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2534_ (.A1(_0736_),
    .A2(_0738_),
    .A3(_0756_),
    .A4(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2535_ (.A1(_0776_),
    .A2(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2536_ (.A1(_0755_),
    .A2(_0780_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2537_ (.A1(net261),
    .A2(_0778_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2538_ (.A1(_0762_),
    .A2(_0781_),
    .B(net262),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2539_ (.A1(net262),
    .A2(_0762_),
    .A3(_0781_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2540_ (.I(net1),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2541_ (.A1(_0782_),
    .A2(_0783_),
    .B(_0784_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2542_ (.I(net263),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2543_ (.A1(net259),
    .A2(net261),
    .A3(net262),
    .A4(_0777_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2544_ (.A1(_0736_),
    .A2(_0738_),
    .A3(_0756_),
    .A4(_0786_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2545_ (.A1(_0785_),
    .A2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2546_ (.A1(_0755_),
    .A2(_0788_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2547_ (.A1(net263),
    .A2(_0786_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2548_ (.A1(_0762_),
    .A2(_0789_),
    .B(net264),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2549_ (.A1(net264),
    .A2(_0762_),
    .A3(_0789_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2550_ (.A1(_0790_),
    .A2(_0791_),
    .B(_0784_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2551_ (.I(net265),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2552_ (.A1(net261),
    .A2(net262),
    .A3(net263),
    .A4(net264),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2553_ (.A1(net259),
    .A2(_0777_),
    .A3(_0793_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2554_ (.A1(_0736_),
    .A2(_0738_),
    .A3(_0756_),
    .A4(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2555_ (.A1(_0792_),
    .A2(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2556_ (.A1(_0755_),
    .A2(_0796_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2557_ (.A1(net265),
    .A2(_0794_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2558_ (.A1(_0762_),
    .A2(_0797_),
    .B(net266),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _2559_ (.A1(net266),
    .A2(_0762_),
    .A3(_0797_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2560_ (.A1(_0798_),
    .A2(_0799_),
    .B(_0784_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2561_ (.A1(_1133_),
    .A2(net10),
    .A3(_1134_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2562_ (.A1(net267),
    .A2(_0800_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2563_ (.A1(_0755_),
    .A2(_0801_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2564_ (.I0(net268),
    .I1(_1455_),
    .S(_0800_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2565_ (.A1(_0755_),
    .A2(_0802_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2566_ (.A1(_1454_),
    .A2(_0800_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2567_ (.A1(net269),
    .A2(_0803_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2568_ (.A1(_0755_),
    .A2(_0804_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _2569_ (.A1(net267),
    .A2(net268),
    .A3(net269),
    .A4(_0800_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _2570_ (.A1(net270),
    .A2(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2571_ (.A1(_1143_),
    .A2(_0806_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2572_ (.A1(_1170_),
    .A2(_1205_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2573_ (.A1(net271),
    .A2(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2574_ (.A1(_1127_),
    .A2(_0808_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2575_ (.I0(net7),
    .I1(\prev_event_inc[0] ),
    .S(_0784_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2576_ (.I0(net8),
    .I1(\prev_event_inc[1] ),
    .S(_0784_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2577_ (.I0(net9),
    .I1(\prev_event_inc[2] ),
    .S(_0784_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2578_ (.I0(net10),
    .I1(\prev_event_inc[3] ),
    .S(_0784_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2579_ (.I0(net11),
    .I1(\prev_event_inc[4] ),
    .S(_0784_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2580_ (.I0(net12),
    .I1(\prev_event_inc[5] ),
    .S(_0784_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2581_ (.I0(net13),
    .I1(\prev_event_inc[6] ),
    .S(_0784_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2582_ (.I0(net14),
    .I1(\prev_event_inc[7] ),
    .S(_1200_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2583_ (.I(net5),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2584_ (.I(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2585_ (.I(counter_sel[4]),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2586_ (.I(_0811_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2587_ (.I(counter_sel[2]),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2588_ (.I(_0813_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2589_ (.I(net2),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _2590_ (.I(net3),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2591_ (.I(_0816_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2592_ (.A1(net16),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2593_ (.I(net3),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2594_ (.I(_0813_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2595_ (.A1(net197),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2596_ (.I(counter_sel[3]),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2597_ (.I(_0822_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2598_ (.A1(_0670_),
    .A2(_0814_),
    .B1(_0818_),
    .B2(_0821_),
    .C(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2599_ (.A1(net267),
    .A2(_0823_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2600_ (.I(counter_sel[5]),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2601_ (.I(_0826_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2602_ (.A1(_1234_),
    .A2(_0811_),
    .B(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2603_ (.A1(_0812_),
    .A2(_0824_),
    .A3(_0825_),
    .B(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2604_ (.A1(net4),
    .A2(net5),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2605_ (.I(_0830_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2606_ (.A1(net83),
    .A2(_0827_),
    .B(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _2607_ (.I(net4),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2608_ (.I(_0809_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2609_ (.A1(net118),
    .A2(_0833_),
    .A3(_0834_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2610_ (.A1(_0409_),
    .A2(_0810_),
    .B1(_0829_),
    .B2(_0832_),
    .C(_0835_),
    .ZN(net272));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2611_ (.A1(net27),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2612_ (.A1(net208),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2613_ (.A1(_0709_),
    .A2(_0814_),
    .B1(_0836_),
    .B2(_0837_),
    .C(_0823_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _2614_ (.I(_0822_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2615_ (.A1(_0839_),
    .A2(net23),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2616_ (.I(_0811_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2617_ (.A1(_0841_),
    .A2(_1274_),
    .B(_0827_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2618_ (.A1(_0812_),
    .A2(_0838_),
    .A3(_0840_),
    .B(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2619_ (.I(_0826_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2620_ (.A1(_0844_),
    .A2(net94),
    .B(_0831_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2621_ (.I(_0833_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2622_ (.A1(_0846_),
    .A2(net130),
    .A3(_0834_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2623_ (.A1(_0448_),
    .A2(_0810_),
    .B1(_0843_),
    .B2(_0845_),
    .C(_0847_),
    .ZN(net273));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2624_ (.A1(net38),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2625_ (.A1(net209),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2626_ (.A1(_0712_),
    .A2(_0814_),
    .B1(_0848_),
    .B2(_0849_),
    .C(_0823_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2627_ (.A1(_0839_),
    .A2(net24),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2628_ (.A1(_0841_),
    .A2(_1277_),
    .B(_0827_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2629_ (.A1(_0812_),
    .A2(_0850_),
    .A3(_0851_),
    .B(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2630_ (.A1(_0844_),
    .A2(net95),
    .B(_0831_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2631_ (.A1(_0846_),
    .A2(net131),
    .A3(_0834_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2632_ (.A1(_0451_),
    .A2(_0810_),
    .B1(_0853_),
    .B2(_0854_),
    .C(_0855_),
    .ZN(net274));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2633_ (.A1(net49),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2634_ (.A1(net210),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2635_ (.A1(_0717_),
    .A2(_0814_),
    .B1(_0856_),
    .B2(_0857_),
    .C(_0823_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2636_ (.A1(_0839_),
    .A2(net25),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2637_ (.A1(_0841_),
    .A2(_1286_),
    .B(_0827_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2638_ (.A1(_0812_),
    .A2(_0858_),
    .A3(_0859_),
    .B(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2639_ (.A1(_0844_),
    .A2(net96),
    .B(_0831_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2640_ (.A1(_0846_),
    .A2(net132),
    .A3(_0834_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2641_ (.A1(_0455_),
    .A2(_0810_),
    .B1(_0861_),
    .B2(_0862_),
    .C(_0863_),
    .ZN(net275));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2642_ (.A1(net60),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2643_ (.A1(net211),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2644_ (.A1(_0720_),
    .A2(_0814_),
    .B1(_0864_),
    .B2(_0865_),
    .C(_0823_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2645_ (.A1(_0839_),
    .A2(net26),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2646_ (.A1(_0841_),
    .A2(_1290_),
    .B(_0827_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2647_ (.A1(_0812_),
    .A2(_0866_),
    .A3(_0867_),
    .B(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2648_ (.A1(_0844_),
    .A2(net97),
    .B(_0831_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2649_ (.A1(_0846_),
    .A2(net133),
    .A3(_0834_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2650_ (.A1(_0458_),
    .A2(_0810_),
    .B1(_0869_),
    .B2(_0870_),
    .C(_0871_),
    .ZN(net276));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2651_ (.A1(net71),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2652_ (.A1(net212),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2653_ (.A1(_0724_),
    .A2(_0814_),
    .B1(_0872_),
    .B2(_0873_),
    .C(_0823_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2654_ (.A1(_0839_),
    .A2(net28),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2655_ (.A1(_0841_),
    .A2(_1293_),
    .B(_0827_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2656_ (.A1(_0812_),
    .A2(_0874_),
    .A3(_0875_),
    .B(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2657_ (.A1(_0844_),
    .A2(net98),
    .B(_0831_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2658_ (.A1(_0846_),
    .A2(net134),
    .A3(_0834_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2659_ (.A1(_0463_),
    .A2(_0810_),
    .B1(_0877_),
    .B2(_0878_),
    .C(_0879_),
    .ZN(net277));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2660_ (.A1(net82),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2661_ (.A1(net213),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2662_ (.A1(_0727_),
    .A2(_0814_),
    .B1(_0880_),
    .B2(_0881_),
    .C(_0823_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2663_ (.A1(_0839_),
    .A2(net29),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2664_ (.A1(_0841_),
    .A2(_1298_),
    .B(_0827_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2665_ (.A1(_0812_),
    .A2(_0882_),
    .A3(_0883_),
    .B(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2666_ (.A1(_0844_),
    .A2(net99),
    .B(_0831_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2667_ (.A1(_0846_),
    .A2(net135),
    .A3(_0834_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2668_ (.A1(_0466_),
    .A2(_0810_),
    .B1(_0885_),
    .B2(_0886_),
    .C(_0887_),
    .ZN(net278));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2669_ (.A1(net93),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2670_ (.A1(net214),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2671_ (.A1(_0733_),
    .A2(_0814_),
    .B1(_0888_),
    .B2(_0889_),
    .C(_0823_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2672_ (.A1(_0839_),
    .A2(net30),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2673_ (.A1(_0841_),
    .A2(_1302_),
    .B(_0827_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2674_ (.A1(_0812_),
    .A2(_0890_),
    .A3(_0891_),
    .B(_0892_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2675_ (.A1(_0844_),
    .A2(net100),
    .B(_0831_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2676_ (.A1(_0846_),
    .A2(net136),
    .A3(_0834_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2677_ (.A1(_0473_),
    .A2(_0810_),
    .B1(_0893_),
    .B2(_0894_),
    .C(_0895_),
    .ZN(net279));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2678_ (.A1(net104),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2679_ (.I(_0813_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2680_ (.A1(net215),
    .A2(_0819_),
    .B(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2681_ (.I(_0822_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2682_ (.A1(_0741_),
    .A2(_0814_),
    .B1(_0896_),
    .B2(_0898_),
    .C(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2683_ (.A1(_0839_),
    .A2(net31),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2684_ (.I(_0826_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2685_ (.A1(_0841_),
    .A2(_1305_),
    .B(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2686_ (.A1(_0812_),
    .A2(_0900_),
    .A3(_0901_),
    .B(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2687_ (.A1(_0844_),
    .A2(net101),
    .B(_0831_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2688_ (.I(_0809_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2689_ (.A1(_0846_),
    .A2(net137),
    .A3(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2690_ (.A1(_0478_),
    .A2(_0810_),
    .B1(_0904_),
    .B2(_0905_),
    .C(_0907_),
    .ZN(net280));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2691_ (.A1(net115),
    .A2(_0815_),
    .A3(_0817_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2692_ (.A1(net217),
    .A2(_0819_),
    .B(_0897_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2693_ (.A1(_0744_),
    .A2(_0814_),
    .B1(_0908_),
    .B2(_0909_),
    .C(_0899_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2694_ (.A1(_0839_),
    .A2(net32),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2695_ (.I(_0811_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2696_ (.A1(_0912_),
    .A2(_1309_),
    .B(_0902_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2697_ (.A1(_0812_),
    .A2(_0910_),
    .A3(_0911_),
    .B(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2698_ (.A1(_0844_),
    .A2(net102),
    .B(_0831_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2699_ (.A1(_0846_),
    .A2(net139),
    .A3(_0906_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2700_ (.A1(_0483_),
    .A2(_0810_),
    .B1(_0914_),
    .B2(_0915_),
    .C(_0916_),
    .ZN(net281));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2701_ (.I(_0809_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2702_ (.I(_0811_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2703_ (.I(_0813_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2704_ (.I(net2),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2705_ (.I(_0816_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2706_ (.A1(net126),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2707_ (.I(net3),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2708_ (.A1(net218),
    .A2(_0923_),
    .B(_0897_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2709_ (.A1(_0747_),
    .A2(_0919_),
    .B1(_0922_),
    .B2(_0924_),
    .C(_0899_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2710_ (.A1(_0839_),
    .A2(net33),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2711_ (.A1(_0912_),
    .A2(_1313_),
    .B(_0902_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2712_ (.A1(_0918_),
    .A2(_0925_),
    .A3(_0926_),
    .B(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2713_ (.I(_0830_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2714_ (.A1(_0844_),
    .A2(net103),
    .B(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2715_ (.A1(_0846_),
    .A2(net140),
    .A3(_0906_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2716_ (.A1(_0487_),
    .A2(_0917_),
    .B1(_0928_),
    .B2(_0930_),
    .C(_0931_),
    .ZN(net282));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2717_ (.I(net155),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2718_ (.I(net233),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2719_ (.A1(net127),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2720_ (.A1(net198),
    .A2(_0923_),
    .B(_0897_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2721_ (.A1(_0933_),
    .A2(_0919_),
    .B1(_0934_),
    .B2(_0935_),
    .C(_0899_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _2722_ (.I(_0822_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2723_ (.A1(_0937_),
    .A2(net268),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2724_ (.I(net48),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2725_ (.A1(_0912_),
    .A2(_0939_),
    .B(_0902_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _2726_ (.A1(_0918_),
    .A2(_0936_),
    .A3(_0938_),
    .B(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2727_ (.I(_0826_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2728_ (.A1(_0942_),
    .A2(net84),
    .B(_0929_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2729_ (.I(_0833_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2730_ (.A1(_0944_),
    .A2(net119),
    .A3(_0906_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2731_ (.A1(_0932_),
    .A2(_0917_),
    .B1(_0941_),
    .B2(_0943_),
    .C(_0945_),
    .ZN(net283));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2732_ (.A1(net138),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2733_ (.A1(net219),
    .A2(_0923_),
    .B(_0897_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2734_ (.A1(_0751_),
    .A2(_0919_),
    .B1(_0946_),
    .B2(_0947_),
    .C(_0899_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2735_ (.A1(_0937_),
    .A2(net34),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2736_ (.A1(_0912_),
    .A2(_1317_),
    .B(_0902_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2737_ (.A1(_0918_),
    .A2(_0948_),
    .A3(_0949_),
    .B(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2738_ (.A1(_0942_),
    .A2(net105),
    .B(_0929_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2739_ (.A1(_0944_),
    .A2(net141),
    .A3(_0906_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2740_ (.A1(_0490_),
    .A2(_0917_),
    .B1(_0951_),
    .B2(_0952_),
    .C(_0953_),
    .ZN(net284));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2741_ (.I(net255),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2742_ (.A1(net149),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2743_ (.A1(net220),
    .A2(_0923_),
    .B(_0897_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2744_ (.A1(_0954_),
    .A2(_0919_),
    .B1(_0955_),
    .B2(_0956_),
    .C(_0899_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2745_ (.A1(_0937_),
    .A2(net35),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2746_ (.A1(_0912_),
    .A2(_1322_),
    .B(_0902_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2747_ (.A1(_0918_),
    .A2(_0957_),
    .A3(_0958_),
    .B(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2748_ (.A1(_0942_),
    .A2(net106),
    .B(_0929_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2749_ (.A1(_0944_),
    .A2(net142),
    .A3(_0906_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2750_ (.A1(_0494_),
    .A2(_0917_),
    .B1(_0960_),
    .B2(_0961_),
    .C(_0962_),
    .ZN(net285));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2751_ (.A1(net160),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2752_ (.A1(net221),
    .A2(_0923_),
    .B(_0897_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2753_ (.A1(_0759_),
    .A2(_0919_),
    .B1(_0963_),
    .B2(_0964_),
    .C(_0899_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2754_ (.A1(_0937_),
    .A2(net36),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2755_ (.A1(_0912_),
    .A2(_1329_),
    .B(_0902_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2756_ (.A1(_0918_),
    .A2(_0965_),
    .A3(_0966_),
    .B(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2757_ (.A1(_0942_),
    .A2(net107),
    .B(_0929_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2758_ (.A1(_0944_),
    .A2(net143),
    .A3(_0906_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2759_ (.A1(_0500_),
    .A2(_0917_),
    .B1(_0968_),
    .B2(_0969_),
    .C(_0970_),
    .ZN(net286));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2760_ (.A1(net171),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2761_ (.A1(net222),
    .A2(_0923_),
    .B(_0897_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2762_ (.A1(_0767_),
    .A2(_0919_),
    .B1(_0971_),
    .B2(_0972_),
    .C(_0899_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2763_ (.A1(_0937_),
    .A2(net37),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2764_ (.A1(_0912_),
    .A2(_1333_),
    .B(_0902_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2765_ (.A1(_0918_),
    .A2(_0973_),
    .A3(_0974_),
    .B(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2766_ (.A1(_0942_),
    .A2(net108),
    .B(_0929_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2767_ (.A1(_0944_),
    .A2(net144),
    .A3(_0906_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2768_ (.A1(_0503_),
    .A2(_0917_),
    .B1(_0976_),
    .B2(_0977_),
    .C(_0978_),
    .ZN(net287));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2769_ (.A1(net182),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2770_ (.A1(net223),
    .A2(_0923_),
    .B(_0897_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2771_ (.A1(_0766_),
    .A2(_0919_),
    .B1(_0979_),
    .B2(_0980_),
    .C(_0899_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2772_ (.A1(_0937_),
    .A2(net39),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2773_ (.A1(_0912_),
    .A2(_1338_),
    .B(_0902_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2774_ (.A1(_0918_),
    .A2(_0981_),
    .A3(_0982_),
    .B(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2775_ (.A1(_0942_),
    .A2(net109),
    .B(_0929_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2776_ (.A1(_0944_),
    .A2(net145),
    .A3(_0906_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2777_ (.A1(_0507_),
    .A2(_0917_),
    .B1(_0984_),
    .B2(_0985_),
    .C(_0986_),
    .ZN(net288));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2778_ (.I(net259),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2779_ (.A1(net189),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2780_ (.A1(net224),
    .A2(_0923_),
    .B(_0897_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2781_ (.A1(_0987_),
    .A2(_0919_),
    .B1(_0988_),
    .B2(_0989_),
    .C(_0899_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2782_ (.A1(_0937_),
    .A2(net40),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2783_ (.A1(_0912_),
    .A2(_1341_),
    .B(_0902_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2784_ (.A1(_0918_),
    .A2(_0990_),
    .A3(_0991_),
    .B(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2785_ (.A1(_0942_),
    .A2(net110),
    .B(_0929_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2786_ (.A1(_0944_),
    .A2(net146),
    .A3(_0906_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2787_ (.A1(_0510_),
    .A2(_0917_),
    .B1(_0993_),
    .B2(_0994_),
    .C(_0995_),
    .ZN(net289));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2788_ (.A1(net190),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2789_ (.I(_0813_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2790_ (.A1(net225),
    .A2(_0923_),
    .B(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2791_ (.I(_0822_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2792_ (.A1(_0776_),
    .A2(_0919_),
    .B1(_0996_),
    .B2(_0998_),
    .C(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2793_ (.A1(_0937_),
    .A2(net41),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2794_ (.I(_0826_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2795_ (.A1(_0912_),
    .A2(_1345_),
    .B(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2796_ (.A1(_0918_),
    .A2(_1000_),
    .A3(_1001_),
    .B(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2797_ (.A1(_0942_),
    .A2(net111),
    .B(_0929_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2798_ (.I(_0809_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2799_ (.A1(_0944_),
    .A2(net147),
    .A3(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2800_ (.A1(_0518_),
    .A2(_0917_),
    .B1(_1004_),
    .B2(_1005_),
    .C(_1007_),
    .ZN(net290));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2801_ (.I(net262),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2802_ (.A1(net191),
    .A2(_0920_),
    .A3(_0921_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2803_ (.A1(net226),
    .A2(_0923_),
    .B(_0997_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2804_ (.A1(_1008_),
    .A2(_0919_),
    .B1(_1009_),
    .B2(_1010_),
    .C(_0999_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2805_ (.A1(_0937_),
    .A2(net42),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2806_ (.I(_0811_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2807_ (.A1(_1013_),
    .A2(_1349_),
    .B(_1002_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2808_ (.A1(_0918_),
    .A2(_1011_),
    .A3(_1012_),
    .B(_1014_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2809_ (.A1(_0942_),
    .A2(net112),
    .B(_0929_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2810_ (.A1(_0944_),
    .A2(net148),
    .A3(_1006_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2811_ (.A1(_0523_),
    .A2(_0917_),
    .B1(_1015_),
    .B2(_1016_),
    .C(_1017_),
    .ZN(net291));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2812_ (.I(_0809_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2813_ (.I(_0811_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _2814_ (.I(_0813_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2815_ (.I(net2),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2816_ (.I(_0816_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2817_ (.A1(net192),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2818_ (.I(net3),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2819_ (.A1(net228),
    .A2(_1024_),
    .B(_0997_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2820_ (.A1(_0785_),
    .A2(_1020_),
    .B1(_1023_),
    .B2(_1025_),
    .C(_0999_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2821_ (.A1(_0937_),
    .A2(net43),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2822_ (.A1(_1013_),
    .A2(_1353_),
    .B(_1002_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2823_ (.A1(_1019_),
    .A2(_1026_),
    .A3(_1027_),
    .B(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2824_ (.I(_0830_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2825_ (.A1(_0942_),
    .A2(net113),
    .B(_1030_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2826_ (.A1(_0944_),
    .A2(net150),
    .A3(_1006_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2827_ (.A1(_0526_),
    .A2(_1018_),
    .B1(_1029_),
    .B2(_1031_),
    .C(_1032_),
    .ZN(net292));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2828_ (.I(net264),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2829_ (.A1(net193),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2830_ (.A1(net229),
    .A2(_1024_),
    .B(_0997_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2831_ (.A1(_1033_),
    .A2(_1020_),
    .B1(_1034_),
    .B2(_1035_),
    .C(_0999_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _2832_ (.I(_0822_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2833_ (.A1(_1037_),
    .A2(net44),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2834_ (.A1(_1013_),
    .A2(_1357_),
    .B(_1002_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2835_ (.A1(_1019_),
    .A2(_1036_),
    .A3(_1038_),
    .B(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2836_ (.I(_0826_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2837_ (.A1(_1041_),
    .A2(net114),
    .B(_1030_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2838_ (.I(_0833_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2839_ (.A1(_1043_),
    .A2(net151),
    .A3(_1006_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2840_ (.A1(_0530_),
    .A2(_1018_),
    .B1(_1040_),
    .B2(_1042_),
    .C(_1044_),
    .ZN(net293));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2841_ (.A1(net194),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2842_ (.A1(net199),
    .A2(_1024_),
    .B(_0997_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2843_ (.A1(_0675_),
    .A2(_1020_),
    .B1(_1045_),
    .B2(_1046_),
    .C(_0999_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2844_ (.A1(_1037_),
    .A2(net269),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2845_ (.A1(_1013_),
    .A2(_1243_),
    .B(_1002_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2846_ (.A1(_1019_),
    .A2(_1047_),
    .A3(_1048_),
    .B(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2847_ (.A1(_1041_),
    .A2(net85),
    .B(_1030_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2848_ (.A1(_1043_),
    .A2(net120),
    .A3(_1006_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2849_ (.A1(_0415_),
    .A2(_1018_),
    .B1(_1050_),
    .B2(_1051_),
    .C(_1052_),
    .ZN(net294));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2850_ (.A1(net195),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2851_ (.A1(net230),
    .A2(_1024_),
    .B(_0997_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2852_ (.A1(_0792_),
    .A2(_1020_),
    .B1(_1053_),
    .B2(_1054_),
    .C(_0999_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2853_ (.A1(_1037_),
    .A2(net45),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2854_ (.A1(_1013_),
    .A2(_1361_),
    .B(_1002_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2855_ (.A1(_1019_),
    .A2(_1055_),
    .A3(_1056_),
    .B(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2856_ (.A1(_1041_),
    .A2(net116),
    .B(_1030_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2857_ (.A1(_1043_),
    .A2(net152),
    .A3(_1006_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2858_ (.A1(_0533_),
    .A2(_1018_),
    .B1(_1058_),
    .B2(_1059_),
    .C(_1060_),
    .ZN(net295));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2859_ (.I(net266),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2860_ (.A1(net196),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2861_ (.A1(net231),
    .A2(_1024_),
    .B(_0997_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2862_ (.A1(_1061_),
    .A2(_1020_),
    .B1(_1062_),
    .B2(_1063_),
    .C(_0999_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2863_ (.A1(_1037_),
    .A2(net46),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2864_ (.A1(_1013_),
    .A2(_1366_),
    .B(_1002_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2865_ (.A1(_1019_),
    .A2(_1064_),
    .A3(_1065_),
    .B(_1066_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2866_ (.A1(_1041_),
    .A2(net117),
    .B(_1030_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2867_ (.A1(_1043_),
    .A2(net153),
    .A3(_1006_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2868_ (.A1(_0538_),
    .A2(_1018_),
    .B1(_1067_),
    .B2(_1068_),
    .C(_1069_),
    .ZN(net296));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2869_ (.A1(net205),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2870_ (.A1(net200),
    .A2(_1024_),
    .B(_0997_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2871_ (.A1(_0679_),
    .A2(_1020_),
    .B1(_1070_),
    .B2(_1071_),
    .C(_0999_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2872_ (.A1(_1037_),
    .A2(net270),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2873_ (.A1(_1013_),
    .A2(_1247_),
    .B(_1002_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2874_ (.A1(_1019_),
    .A2(_1072_),
    .A3(_1073_),
    .B(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2875_ (.A1(_1041_),
    .A2(net86),
    .B(_1030_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2876_ (.A1(_1043_),
    .A2(net121),
    .A3(_1006_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2877_ (.A1(_0418_),
    .A2(_1018_),
    .B1(_1075_),
    .B2(_1076_),
    .C(_1077_),
    .ZN(net297));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2878_ (.A1(net216),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2879_ (.A1(_0575_),
    .A2(_1024_),
    .B(_0997_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2880_ (.A1(_0684_),
    .A2(_1020_),
    .B1(_1078_),
    .B2(_1079_),
    .C(_0999_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2881_ (.A1(_1037_),
    .A2(net17),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2882_ (.A1(_1013_),
    .A2(_1251_),
    .B(_1002_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2883_ (.A1(_1019_),
    .A2(_1080_),
    .A3(_1081_),
    .B(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2884_ (.A1(_1041_),
    .A2(net87),
    .B(_1030_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2885_ (.A1(_1043_),
    .A2(net122),
    .A3(_1006_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2886_ (.A1(_0423_),
    .A2(_1018_),
    .B1(_1083_),
    .B2(_1084_),
    .C(_1085_),
    .ZN(net298));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2887_ (.A1(net227),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2888_ (.A1(net202),
    .A2(_1024_),
    .B(_0997_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2889_ (.A1(_0688_),
    .A2(_1020_),
    .B1(_1086_),
    .B2(_1087_),
    .C(_0999_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2890_ (.A1(_1037_),
    .A2(net18),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2891_ (.A1(_1013_),
    .A2(_1256_),
    .B(_1002_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2892_ (.A1(_1019_),
    .A2(_1088_),
    .A3(_1089_),
    .B(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2893_ (.A1(_1041_),
    .A2(net88),
    .B(_1030_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _2894_ (.A1(_1043_),
    .A2(net123),
    .A3(_1006_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2895_ (.A1(_0426_),
    .A2(_1018_),
    .B1(_1091_),
    .B2(_1092_),
    .C(_1093_),
    .ZN(net299));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2896_ (.A1(net238),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2897_ (.A1(net203),
    .A2(_1024_),
    .B(_0813_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2898_ (.A1(_0695_),
    .A2(_1020_),
    .B1(_1094_),
    .B2(_1095_),
    .C(_0822_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2899_ (.A1(_1037_),
    .A2(net19),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2900_ (.A1(_1013_),
    .A2(_1259_),
    .B(_0826_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2901_ (.A1(_1019_),
    .A2(_1096_),
    .A3(_1097_),
    .B(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2902_ (.A1(_1041_),
    .A2(net89),
    .B(_1030_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2903_ (.A1(_1043_),
    .A2(net124),
    .A3(_0809_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2904_ (.A1(_0433_),
    .A2(_1018_),
    .B1(_1099_),
    .B2(_1100_),
    .C(_1101_),
    .ZN(net300));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2905_ (.A1(net249),
    .A2(_1021_),
    .A3(_1022_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2906_ (.A1(net204),
    .A2(_1024_),
    .B(_0813_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2907_ (.A1(_0698_),
    .A2(_1020_),
    .B1(_1102_),
    .B2(_1103_),
    .C(_0822_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2908_ (.A1(_1037_),
    .A2(net20),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2909_ (.A1(_0811_),
    .A2(_1263_),
    .B(_0826_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2910_ (.A1(_1019_),
    .A2(_1104_),
    .A3(_1105_),
    .B(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2911_ (.A1(_1041_),
    .A2(net90),
    .B(_1030_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2912_ (.A1(_1043_),
    .A2(net125),
    .A3(_0809_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2913_ (.A1(_0437_),
    .A2(_1018_),
    .B1(_1107_),
    .B2(_1108_),
    .C(_1109_),
    .ZN(net301));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2914_ (.A1(net260),
    .A2(net2),
    .A3(_0816_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2915_ (.A1(net206),
    .A2(net3),
    .B(_0813_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2916_ (.A1(_0701_),
    .A2(_0820_),
    .B1(_1110_),
    .B2(_1111_),
    .C(_0822_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2917_ (.A1(_1037_),
    .A2(net21),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2918_ (.A1(_0811_),
    .A2(_1267_),
    .B(_0826_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2919_ (.A1(_0841_),
    .A2(_1112_),
    .A3(_1113_),
    .B(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2920_ (.A1(_1041_),
    .A2(net91),
    .B(_0830_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2921_ (.A1(_1043_),
    .A2(net128),
    .A3(_0809_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2922_ (.A1(_0440_),
    .A2(_0834_),
    .B1(_1115_),
    .B2(_1116_),
    .C(_1117_),
    .ZN(net302));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _2923_ (.A1(net271),
    .A2(net2),
    .A3(_0816_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2924_ (.A1(net207),
    .A2(net3),
    .B(_0813_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _2925_ (.A1(_0705_),
    .A2(_0820_),
    .B1(_1118_),
    .B2(_1119_),
    .C(_0822_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2926_ (.A1(_0823_),
    .A2(net22),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2927_ (.A1(_0811_),
    .A2(_1270_),
    .B(_0826_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2928_ (.A1(_0841_),
    .A2(_1120_),
    .A3(_1121_),
    .B(_1122_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2929_ (.A1(_0827_),
    .A2(net92),
    .B(_0830_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _2930_ (.A1(_0833_),
    .A2(net129),
    .A3(_0809_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2931_ (.A1(_0444_),
    .A2(_0834_),
    .B1(_1123_),
    .B2(_1124_),
    .C(_1125_),
    .ZN(net303));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2932_ (.A(net197),
    .B(net198),
    .CO(_1442_),
    .S(_1443_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2933_ (.A(net16),
    .B(net127),
    .CO(_1444_),
    .S(_1445_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2934_ (.A(net154),
    .B(net155),
    .CO(_1446_),
    .S(_1447_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2935_ (.A(net118),
    .B(net119),
    .CO(_1448_),
    .S(_1449_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _2936_ (.A(net83),
    .B(net84),
    .CO(_1450_),
    .S(_1451_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2937_ (.A(net47),
    .B(net48),
    .CO(_1452_),
    .S(_1453_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2938_ (.A(net267),
    .B(net268),
    .CO(_1454_),
    .S(_1455_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _2939_ (.A(net232),
    .B(net233),
    .CO(_1456_),
    .S(_1457_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[0]$_DFFE_PN0P_  (.D(_0000_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[100]$_DFFE_PN0P_  (.D(_0001_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[101]$_DFFE_PN0P_  (.D(_0002_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[102]$_DFFE_PN0P_  (.D(_0003_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[103]$_DFFE_PN0P_  (.D(_0004_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[104]$_DFFE_PN0P_  (.D(_0005_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[105]$_DFFE_PN0P_  (.D(_0006_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[106]$_DFFE_PN0P_  (.D(_0007_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[107]$_DFFE_PN0P_  (.D(_0008_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[108]$_DFFE_PN0P_  (.D(_0009_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[109]$_DFFE_PN0P_  (.D(_0010_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[10]$_DFFE_PN0P_  (.D(_0011_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[110]$_DFFE_PN0P_  (.D(_0012_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[111]$_DFFE_PN0P_  (.D(_0013_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[112]$_DFFE_PN0P_  (.D(_0014_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[113]$_DFFE_PN0P_  (.D(_0015_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[114]$_DFFE_PN0P_  (.D(_0016_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[115]$_DFFE_PN0P_  (.D(_0017_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[116]$_DFFE_PN0P_  (.D(_0018_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net34));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[117]$_DFFE_PN0P_  (.D(_0019_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net35));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[118]$_DFFE_PN0P_  (.D(_0020_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net36));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[119]$_DFFE_PN0P_  (.D(_0021_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net37));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[11]$_DFFE_PN0P_  (.D(_0022_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net38));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[120]$_DFFE_PN0P_  (.D(_0023_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net39));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[121]$_DFFE_PN0P_  (.D(_0024_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net40));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[122]$_DFFE_PN0P_  (.D(_0025_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net41));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[123]$_DFFE_PN0P_  (.D(_0026_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net42));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[124]$_DFFE_PN0P_  (.D(_0027_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net43));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[125]$_DFFE_PN0P_  (.D(_0028_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net44));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[126]$_DFFE_PN0P_  (.D(_0029_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net45));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[127]$_DFFE_PN0P_  (.D(_0030_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net46));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[128]$_DFFE_PN0P_  (.D(_0031_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net47));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[129]$_DFFE_PN0P_  (.D(_0032_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net48));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[12]$_DFFE_PN0P_  (.D(_0033_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net49));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[130]$_DFFE_PN0P_  (.D(_0034_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net50));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[131]$_DFFE_PN0P_  (.D(_0035_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net51));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[132]$_DFFE_PN0P_  (.D(_0036_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net52));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[133]$_DFFE_PN0P_  (.D(_0037_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net53));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[134]$_DFFE_PN0P_  (.D(_0038_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net54));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[135]$_DFFE_PN0P_  (.D(_0039_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net55));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[136]$_DFFE_PN0P_  (.D(_0040_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net56));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[137]$_DFFE_PN0P_  (.D(_0041_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net57));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[138]$_DFFE_PN0P_  (.D(_0042_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net58));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[139]$_DFFE_PN0P_  (.D(_0043_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net59));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[13]$_DFFE_PN0P_  (.D(_0044_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net60));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[140]$_DFFE_PN0P_  (.D(_0045_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net61));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[141]$_DFFE_PN0P_  (.D(_0046_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net62));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[142]$_DFFE_PN0P_  (.D(_0047_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net63));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[143]$_DFFE_PN0P_  (.D(_0048_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net64));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[144]$_DFFE_PN0P_  (.D(_0049_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net65));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[145]$_DFFE_PN0P_  (.D(_0050_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net66));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[146]$_DFFE_PN0P_  (.D(_0051_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net67));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[147]$_DFFE_PN0P_  (.D(_0052_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net68));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[148]$_DFFE_PN0P_  (.D(_0053_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net69));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[149]$_DFFE_PN0P_  (.D(_0054_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net70));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[14]$_DFFE_PN0P_  (.D(_0055_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net71));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[150]$_DFFE_PN0P_  (.D(_0056_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net72));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[151]$_DFFE_PN0P_  (.D(_0057_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net73));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[152]$_DFFE_PN0P_  (.D(_0058_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net74));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[153]$_DFFE_PN0P_  (.D(_0059_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net75));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[154]$_DFFE_PN0P_  (.D(_0060_),
    .RN(net15),
    .CLK(clknet_leaf_2_clk),
    .Q(net76));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[155]$_DFFE_PN0P_  (.D(_0061_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net77));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[156]$_DFFE_PN0P_  (.D(_0062_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net78));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[157]$_DFFE_PN0P_  (.D(_0063_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net79));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[158]$_DFFE_PN0P_  (.D(_0064_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net80));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[159]$_DFFE_PN0P_  (.D(_0065_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net81));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[15]$_DFFE_PN0P_  (.D(_0066_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net82));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[160]$_DFFE_PN0P_  (.D(_0067_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net83));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[161]$_DFFE_PN0P_  (.D(_0068_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net84));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[162]$_DFFE_PN0P_  (.D(_0069_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net85));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[163]$_DFFE_PN0P_  (.D(_0070_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net86));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[164]$_DFFE_PN0P_  (.D(_0071_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net87));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[165]$_DFFE_PN0P_  (.D(_0072_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net88));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[166]$_DFFE_PN0P_  (.D(_0073_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net89));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[167]$_DFFE_PN0P_  (.D(_0074_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net90));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[168]$_DFFE_PN0P_  (.D(_0075_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net91));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[169]$_DFFE_PN0P_  (.D(_0076_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net92));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[16]$_DFFE_PN0P_  (.D(_0077_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net93));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[170]$_DFFE_PN0P_  (.D(_0078_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net94));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[171]$_DFFE_PN0P_  (.D(_0079_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net95));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[172]$_DFFE_PN0P_  (.D(_0080_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net96));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[173]$_DFFE_PN0P_  (.D(_0081_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net97));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[174]$_DFFE_PN0P_  (.D(_0082_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net98));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[175]$_DFFE_PN0P_  (.D(_0083_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net99));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[176]$_DFFE_PN0P_  (.D(_0084_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net100));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[177]$_DFFE_PN0P_  (.D(_0085_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net101));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[178]$_DFFE_PN0P_  (.D(_0086_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net102));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[179]$_DFFE_PN0P_  (.D(_0087_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net103));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[17]$_DFFE_PN0P_  (.D(_0088_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net104));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[180]$_DFFE_PN0P_  (.D(_0089_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net105));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[181]$_DFFE_PN0P_  (.D(_0090_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net106));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[182]$_DFFE_PN0P_  (.D(_0091_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net107));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[183]$_DFFE_PN0P_  (.D(_0092_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net108));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[184]$_DFFE_PN0P_  (.D(_0093_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net109));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[185]$_DFFE_PN0P_  (.D(_0094_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net110));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[186]$_DFFE_PN0P_  (.D(_0095_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net111));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[187]$_DFFE_PN0P_  (.D(_0096_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net112));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[188]$_DFFE_PN0P_  (.D(_0097_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(net113));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[189]$_DFFE_PN0P_  (.D(_0098_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net114));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[18]$_DFFE_PN0P_  (.D(_0099_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net115));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[190]$_DFFE_PN0P_  (.D(_0100_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net116));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[191]$_DFFE_PN0P_  (.D(_0101_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net117));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[192]$_DFFE_PN0P_  (.D(_0102_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net118));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[193]$_DFFE_PN0P_  (.D(_0103_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net119));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[194]$_DFFE_PN0P_  (.D(_0104_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net120));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[195]$_DFFE_PN0P_  (.D(_0105_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net121));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[196]$_DFFE_PN0P_  (.D(_0106_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net122));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[197]$_DFFE_PN0P_  (.D(_0107_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net123));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[198]$_DFFE_PN0P_  (.D(_0108_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net124));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[199]$_DFFE_PN0P_  (.D(_0109_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net125));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[19]$_DFFE_PN0P_  (.D(_0110_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net126));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[1]$_DFFE_PN0P_  (.D(_0111_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net127));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[200]$_DFFE_PN0P_  (.D(_0112_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net128));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[201]$_DFFE_PN0P_  (.D(_0113_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net129));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[202]$_DFFE_PN0P_  (.D(_0114_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net130));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[203]$_DFFE_PN0P_  (.D(_0115_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net131));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[204]$_DFFE_PN0P_  (.D(_0116_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net132));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[205]$_DFFE_PN0P_  (.D(_0117_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net133));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[206]$_DFFE_PN0P_  (.D(_0118_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net134));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[207]$_DFFE_PN0P_  (.D(_0119_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net135));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[208]$_DFFE_PN0P_  (.D(_0120_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net136));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[209]$_DFFE_PN0P_  (.D(_0121_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net137));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[20]$_DFFE_PN0P_  (.D(_0122_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net138));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[210]$_DFFE_PN0P_  (.D(_0123_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net139));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[211]$_DFFE_PN0P_  (.D(_0124_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net140));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[212]$_DFFE_PN0P_  (.D(_0125_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net141));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[213]$_DFFE_PN0P_  (.D(_0126_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net142));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[214]$_DFFE_PN0P_  (.D(_0127_),
    .RN(net15),
    .CLK(clknet_leaf_6_clk),
    .Q(net143));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[215]$_DFFE_PN0P_  (.D(_0128_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net144));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[216]$_DFFE_PN0P_  (.D(_0129_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net145));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[217]$_DFFE_PN0P_  (.D(_0130_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net146));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[218]$_DFFE_PN0P_  (.D(_0131_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net147));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[219]$_DFFE_PN0P_  (.D(_0132_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net148));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[21]$_DFFE_PN0P_  (.D(_0133_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net149));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[220]$_DFFE_PN0P_  (.D(_0134_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net150));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[221]$_DFFE_PN0P_  (.D(_0135_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net151));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[222]$_DFFE_PN0P_  (.D(_0136_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net152));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[223]$_DFFE_PN0P_  (.D(_0137_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net153));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[224]$_DFFE_PN0P_  (.D(_0138_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net154));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[225]$_DFFE_PN0P_  (.D(_0139_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net155));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[226]$_DFFE_PN0P_  (.D(_0140_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net156));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[227]$_DFFE_PN0P_  (.D(_0141_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net157));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[228]$_DFFE_PN0P_  (.D(_0142_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net158));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[229]$_DFFE_PN0P_  (.D(_0143_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net159));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[22]$_DFFE_PN0P_  (.D(_0144_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net160));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[230]$_DFFE_PN0P_  (.D(_0145_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net161));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[231]$_DFFE_PN0P_  (.D(_0146_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(net162));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[232]$_DFFE_PN0P_  (.D(_0147_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net163));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[233]$_DFFE_PN0P_  (.D(_0148_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net164));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[234]$_DFFE_PN0P_  (.D(_0149_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net165));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[235]$_DFFE_PN0P_  (.D(_0150_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net166));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[236]$_DFFE_PN0P_  (.D(_0151_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net167));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[237]$_DFFE_PN0P_  (.D(_0152_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net168));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[238]$_DFFE_PN0P_  (.D(_0153_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net169));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[239]$_DFFE_PN0P_  (.D(_0154_),
    .RN(net15),
    .CLK(clknet_leaf_4_clk),
    .Q(net170));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[23]$_DFFE_PN0P_  (.D(_0155_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net171));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[240]$_DFFE_PN0P_  (.D(_0156_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net172));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[241]$_DFFE_PN0P_  (.D(_0157_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net173));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[242]$_DFFE_PN0P_  (.D(_0158_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net174));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[243]$_DFFE_PN0P_  (.D(_0159_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net175));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[244]$_DFFE_PN0P_  (.D(_0160_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net176));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[245]$_DFFE_PN0P_  (.D(_0161_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net177));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[246]$_DFFE_PN0P_  (.D(_0162_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net178));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[247]$_DFFE_PN0P_  (.D(_0163_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net179));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[248]$_DFFE_PN0P_  (.D(_0164_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net180));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[249]$_DFFE_PN0P_  (.D(_0165_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net181));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[24]$_DFFE_PN0P_  (.D(_0166_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(net182));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[250]$_DFFE_PN0P_  (.D(_0167_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net183));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[251]$_DFFE_PN0P_  (.D(_0168_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net184));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[252]$_DFFE_PN0P_  (.D(_0169_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net185));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[253]$_DFFE_PN0P_  (.D(_0170_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net186));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[254]$_DFFE_PN0P_  (.D(_0171_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net187));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[255]$_DFFE_PN0P_  (.D(_0172_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net188));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[25]$_DFFE_PN0P_  (.D(_0173_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net189));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[26]$_DFFE_PN0P_  (.D(_0174_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net190));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[27]$_DFFE_PN0P_  (.D(_0175_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net191));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[28]$_DFFE_PN0P_  (.D(_0176_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net192));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[29]$_DFFE_PN0P_  (.D(_0177_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net193));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[2]$_DFFE_PN0P_  (.D(_0178_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net194));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[30]$_DFFE_PN0P_  (.D(_0179_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net195));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[31]$_DFFE_PN0P_  (.D(_0180_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net196));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[32]$_DFFE_PN0P_  (.D(_0181_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net197));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[33]$_DFFE_PN0P_  (.D(_0182_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net198));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[34]$_DFFE_PN0P_  (.D(_0183_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net199));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[35]$_DFFE_PN0P_  (.D(_0184_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net200));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[36]$_DFFE_PN0P_  (.D(_0185_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net201));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[37]$_DFFE_PN0P_  (.D(_0186_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net202));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[38]$_DFFE_PN0P_  (.D(_0187_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net203));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[39]$_DFFE_PN0P_  (.D(_0188_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net204));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[3]$_DFFE_PN0P_  (.D(_0189_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net205));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[40]$_DFFE_PN0P_  (.D(_0190_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net206));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[41]$_DFFE_PN0P_  (.D(_0191_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net207));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[42]$_DFFE_PN0P_  (.D(_0192_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net208));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[43]$_DFFE_PN0P_  (.D(_0193_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net209));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[44]$_DFFE_PN0P_  (.D(_0194_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net210));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[45]$_DFFE_PN0P_  (.D(_0195_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net211));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[46]$_DFFE_PN0P_  (.D(_0196_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net212));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[47]$_DFFE_PN0P_  (.D(_0197_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net213));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[48]$_DFFE_PN0P_  (.D(_0198_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net214));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[49]$_DFFE_PN0P_  (.D(_0199_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net215));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[4]$_DFFE_PN0P_  (.D(_0200_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net216));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[50]$_DFFE_PN0P_  (.D(_0201_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net217));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[51]$_DFFE_PN0P_  (.D(_0202_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net218));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[52]$_DFFE_PN0P_  (.D(_0203_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net219));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[53]$_DFFE_PN0P_  (.D(_0204_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net220));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[54]$_DFFE_PN0P_  (.D(_0205_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net221));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[55]$_DFFE_PN0P_  (.D(_0206_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net222));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[56]$_DFFE_PN0P_  (.D(_0207_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net223));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[57]$_DFFE_PN0P_  (.D(_0208_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net224));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[58]$_DFFE_PN0P_  (.D(_0209_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net225));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[59]$_DFFE_PN0P_  (.D(_0210_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net226));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[5]$_DFFE_PN0P_  (.D(_0211_),
    .RN(net15),
    .CLK(clknet_leaf_11_clk),
    .Q(net227));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[60]$_DFFE_PN0P_  (.D(_0212_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net228));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[61]$_DFFE_PN0P_  (.D(_0213_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net229));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[62]$_DFFE_PN0P_  (.D(_0214_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net230));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[63]$_DFFE_PN0P_  (.D(_0215_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net231));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[64]$_DFFE_PN0P_  (.D(_0216_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net232));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[65]$_DFFE_PN0P_  (.D(_0217_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net233));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[66]$_DFFE_PN0P_  (.D(_0218_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net234));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[67]$_DFFE_PN0P_  (.D(_0219_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net235));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[68]$_DFFE_PN0P_  (.D(_0220_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net236));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[69]$_DFFE_PN0P_  (.D(_0221_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net237));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[6]$_DFFE_PN0P_  (.D(_0222_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net238));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[70]$_DFFE_PN0P_  (.D(_0223_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net239));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[71]$_DFFE_PN0P_  (.D(_0224_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net240));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[72]$_DFFE_PN0P_  (.D(_0225_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net241));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[73]$_DFFE_PN0P_  (.D(_0226_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net242));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[74]$_DFFE_PN0P_  (.D(_0227_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net243));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[75]$_DFFE_PN0P_  (.D(_0228_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net244));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[76]$_DFFE_PN0P_  (.D(_0229_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net245));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[77]$_DFFE_PN0P_  (.D(_0230_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net246));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[78]$_DFFE_PN0P_  (.D(_0231_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net247));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[79]$_DFFE_PN0P_  (.D(_0232_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net248));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[7]$_DFFE_PN0P_  (.D(_0233_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net249));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[80]$_DFFE_PN0P_  (.D(_0234_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net250));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[81]$_DFFE_PN0P_  (.D(_0235_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net251));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[82]$_DFFE_PN0P_  (.D(_0236_),
    .RN(net15),
    .CLK(clknet_leaf_12_clk),
    .Q(net252));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[83]$_DFFE_PN0P_  (.D(_0237_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net253));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[84]$_DFFE_PN0P_  (.D(_0238_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(net254));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[85]$_DFFE_PN0P_  (.D(_0239_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net255));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[86]$_DFFE_PN0P_  (.D(_0240_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net256));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[87]$_DFFE_PN0P_  (.D(_0241_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net257));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[88]$_DFFE_PN0P_  (.D(_0242_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net258));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[89]$_DFFE_PN0P_  (.D(_0243_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net259));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[8]$_DFFE_PN0P_  (.D(_0244_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net260));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[90]$_DFFE_PN0P_  (.D(_0245_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net261));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[91]$_DFFE_PN0P_  (.D(_0246_),
    .RN(net15),
    .CLK(clknet_leaf_8_clk),
    .Q(net262));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[92]$_DFFE_PN0P_  (.D(_0247_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net263));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[93]$_DFFE_PN0P_  (.D(_0248_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net264));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[94]$_DFFE_PN0P_  (.D(_0249_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net265));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[95]$_DFFE_PN0P_  (.D(_0250_),
    .RN(net15),
    .CLK(clknet_leaf_9_clk),
    .Q(net266));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[96]$_DFFE_PN0P_  (.D(_0251_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net267));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[97]$_DFFE_PN0P_  (.D(_0252_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(net268));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[98]$_DFFE_PN0P_  (.D(_0253_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net269));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[99]$_DFFE_PN0P_  (.D(_0254_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net270));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counters[9]$_DFFE_PN0P_  (.D(_0255_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(net271));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \prev_event_inc[0]$_DFFE_PN0N_  (.D(_0256_),
    .RN(net15),
    .CLK(clknet_leaf_0_clk),
    .Q(\prev_event_inc[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \prev_event_inc[1]$_DFFE_PN0N_  (.D(_0257_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(\prev_event_inc[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \prev_event_inc[2]$_DFFE_PN0N_  (.D(_0258_),
    .RN(net15),
    .CLK(clknet_leaf_10_clk),
    .Q(\prev_event_inc[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \prev_event_inc[3]$_DFFE_PN0N_  (.D(_0259_),
    .RN(net15),
    .CLK(clknet_leaf_1_clk),
    .Q(\prev_event_inc[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \prev_event_inc[4]$_DFFE_PN0N_  (.D(_0260_),
    .RN(net15),
    .CLK(clknet_leaf_3_clk),
    .Q(\prev_event_inc[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \prev_event_inc[5]$_DFFE_PN0N_  (.D(_0261_),
    .RN(net15),
    .CLK(clknet_leaf_5_clk),
    .Q(\prev_event_inc[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \prev_event_inc[6]$_DFFE_PN0N_  (.D(_0262_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(\prev_event_inc[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \prev_event_inc[7]$_DFFE_PN0N_  (.D(_0263_),
    .RN(net15),
    .CLK(clknet_leaf_7_clk),
    .Q(\prev_event_inc[7] ));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_347 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input1 (.I(net307),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input2 (.I(counter_sel[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input3 (.I(counter_sel[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input4 (.I(counter_sel[6]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input5 (.I(counter_sel[7]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input6 (.I(enable),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(event_inc[0]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(event_inc[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input9 (.I(net304),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input10 (.I(net306),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(event_inc[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(event_inc[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(event_inc[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input14 (.I(event_inc[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input15 (.I(net305),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net16),
    .Z(all_counts[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net17),
    .Z(all_counts[100]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net18),
    .Z(all_counts[101]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net19),
    .Z(all_counts[102]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net20),
    .Z(all_counts[103]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net21),
    .Z(all_counts[104]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net22),
    .Z(all_counts[105]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net23),
    .Z(all_counts[106]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net24),
    .Z(all_counts[107]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output25 (.I(net25),
    .Z(all_counts[108]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output26 (.I(net26),
    .Z(all_counts[109]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output27 (.I(net27),
    .Z(all_counts[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output28 (.I(net28),
    .Z(all_counts[110]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output29 (.I(net29),
    .Z(all_counts[111]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output30 (.I(net30),
    .Z(all_counts[112]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output31 (.I(net31),
    .Z(all_counts[113]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output32 (.I(net32),
    .Z(all_counts[114]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output33 (.I(net33),
    .Z(all_counts[115]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output34 (.I(net34),
    .Z(all_counts[116]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output35 (.I(net35),
    .Z(all_counts[117]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output36 (.I(net36),
    .Z(all_counts[118]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output37 (.I(net37),
    .Z(all_counts[119]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output38 (.I(net38),
    .Z(all_counts[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net39),
    .Z(all_counts[120]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output40 (.I(net40),
    .Z(all_counts[121]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output41 (.I(net41),
    .Z(all_counts[122]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output42 (.I(net42),
    .Z(all_counts[123]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output43 (.I(net43),
    .Z(all_counts[124]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output44 (.I(net44),
    .Z(all_counts[125]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output45 (.I(net45),
    .Z(all_counts[126]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output46 (.I(net46),
    .Z(all_counts[127]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output47 (.I(net47),
    .Z(all_counts[128]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net48),
    .Z(all_counts[129]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net49),
    .Z(all_counts[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net50),
    .Z(all_counts[130]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output51 (.I(net51),
    .Z(all_counts[131]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output52 (.I(net52),
    .Z(all_counts[132]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output53 (.I(net53),
    .Z(all_counts[133]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output54 (.I(net54),
    .Z(all_counts[134]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output55 (.I(net55),
    .Z(all_counts[135]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output56 (.I(net56),
    .Z(all_counts[136]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output57 (.I(net57),
    .Z(all_counts[137]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output58 (.I(net58),
    .Z(all_counts[138]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output59 (.I(net59),
    .Z(all_counts[139]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output60 (.I(net60),
    .Z(all_counts[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output61 (.I(net61),
    .Z(all_counts[140]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net62),
    .Z(all_counts[141]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net63),
    .Z(all_counts[142]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net64),
    .Z(all_counts[143]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net65),
    .Z(all_counts[144]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net66),
    .Z(all_counts[145]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net67),
    .Z(all_counts[146]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net68),
    .Z(all_counts[147]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net69),
    .Z(all_counts[148]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net70),
    .Z(all_counts[149]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net71),
    .Z(all_counts[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net72),
    .Z(all_counts[150]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net73),
    .Z(all_counts[151]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net74),
    .Z(all_counts[152]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net75),
    .Z(all_counts[153]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net76),
    .Z(all_counts[154]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net77),
    .Z(all_counts[155]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net78),
    .Z(all_counts[156]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net79),
    .Z(all_counts[157]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net80),
    .Z(all_counts[158]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net81),
    .Z(all_counts[159]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net82),
    .Z(all_counts[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net83),
    .Z(all_counts[160]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output84 (.I(net84),
    .Z(all_counts[161]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output85 (.I(net85),
    .Z(all_counts[162]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output86 (.I(net86),
    .Z(all_counts[163]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output87 (.I(net87),
    .Z(all_counts[164]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output88 (.I(net88),
    .Z(all_counts[165]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net89),
    .Z(all_counts[166]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output90 (.I(net90),
    .Z(all_counts[167]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output91 (.I(net91),
    .Z(all_counts[168]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net92),
    .Z(all_counts[169]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net93),
    .Z(all_counts[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net94),
    .Z(all_counts[170]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net95),
    .Z(all_counts[171]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net96),
    .Z(all_counts[172]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net97),
    .Z(all_counts[173]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net98),
    .Z(all_counts[174]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output99 (.I(net99),
    .Z(all_counts[175]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output100 (.I(net100),
    .Z(all_counts[176]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output101 (.I(net101),
    .Z(all_counts[177]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output102 (.I(net102),
    .Z(all_counts[178]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output103 (.I(net103),
    .Z(all_counts[179]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output104 (.I(net104),
    .Z(all_counts[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output105 (.I(net105),
    .Z(all_counts[180]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output106 (.I(net106),
    .Z(all_counts[181]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output107 (.I(net107),
    .Z(all_counts[182]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output108 (.I(net108),
    .Z(all_counts[183]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output109 (.I(net109),
    .Z(all_counts[184]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output110 (.I(net110),
    .Z(all_counts[185]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output111 (.I(net111),
    .Z(all_counts[186]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output112 (.I(net112),
    .Z(all_counts[187]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output113 (.I(net113),
    .Z(all_counts[188]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output114 (.I(net114),
    .Z(all_counts[189]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output115 (.I(net115),
    .Z(all_counts[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output116 (.I(net116),
    .Z(all_counts[190]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output117 (.I(net117),
    .Z(all_counts[191]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output118 (.I(net118),
    .Z(all_counts[192]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output119 (.I(net119),
    .Z(all_counts[193]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output120 (.I(net120),
    .Z(all_counts[194]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output121 (.I(net121),
    .Z(all_counts[195]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output122 (.I(net122),
    .Z(all_counts[196]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output123 (.I(net123),
    .Z(all_counts[197]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output124 (.I(net124),
    .Z(all_counts[198]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output125 (.I(net125),
    .Z(all_counts[199]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output126 (.I(net126),
    .Z(all_counts[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output127 (.I(net127),
    .Z(all_counts[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output128 (.I(net128),
    .Z(all_counts[200]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output129 (.I(net129),
    .Z(all_counts[201]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output130 (.I(net130),
    .Z(all_counts[202]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output131 (.I(net131),
    .Z(all_counts[203]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output132 (.I(net132),
    .Z(all_counts[204]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output133 (.I(net133),
    .Z(all_counts[205]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output134 (.I(net134),
    .Z(all_counts[206]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output135 (.I(net135),
    .Z(all_counts[207]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output136 (.I(net136),
    .Z(all_counts[208]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output137 (.I(net137),
    .Z(all_counts[209]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output138 (.I(net138),
    .Z(all_counts[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output139 (.I(net139),
    .Z(all_counts[210]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output140 (.I(net140),
    .Z(all_counts[211]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output141 (.I(net141),
    .Z(all_counts[212]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output142 (.I(net142),
    .Z(all_counts[213]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output143 (.I(net143),
    .Z(all_counts[214]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output144 (.I(net144),
    .Z(all_counts[215]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output145 (.I(net145),
    .Z(all_counts[216]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output146 (.I(net146),
    .Z(all_counts[217]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output147 (.I(net147),
    .Z(all_counts[218]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output148 (.I(net148),
    .Z(all_counts[219]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output149 (.I(net149),
    .Z(all_counts[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output150 (.I(net150),
    .Z(all_counts[220]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output151 (.I(net151),
    .Z(all_counts[221]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output152 (.I(net152),
    .Z(all_counts[222]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output153 (.I(net153),
    .Z(all_counts[223]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output154 (.I(net154),
    .Z(all_counts[224]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output155 (.I(net155),
    .Z(all_counts[225]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output156 (.I(net156),
    .Z(all_counts[226]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output157 (.I(net157),
    .Z(all_counts[227]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output158 (.I(net158),
    .Z(all_counts[228]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output159 (.I(net159),
    .Z(all_counts[229]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output160 (.I(net160),
    .Z(all_counts[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output161 (.I(net161),
    .Z(all_counts[230]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output162 (.I(net162),
    .Z(all_counts[231]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output163 (.I(net163),
    .Z(all_counts[232]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output164 (.I(net164),
    .Z(all_counts[233]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output165 (.I(net165),
    .Z(all_counts[234]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output166 (.I(net166),
    .Z(all_counts[235]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output167 (.I(net167),
    .Z(all_counts[236]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output168 (.I(net168),
    .Z(all_counts[237]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output169 (.I(net169),
    .Z(all_counts[238]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output170 (.I(net170),
    .Z(all_counts[239]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output171 (.I(net171),
    .Z(all_counts[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output172 (.I(net172),
    .Z(all_counts[240]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output173 (.I(net173),
    .Z(all_counts[241]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output174 (.I(net174),
    .Z(all_counts[242]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output175 (.I(net175),
    .Z(all_counts[243]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output176 (.I(net176),
    .Z(all_counts[244]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output177 (.I(net177),
    .Z(all_counts[245]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output178 (.I(net178),
    .Z(all_counts[246]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output179 (.I(net179),
    .Z(all_counts[247]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output180 (.I(net180),
    .Z(all_counts[248]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output181 (.I(net181),
    .Z(all_counts[249]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output182 (.I(net182),
    .Z(all_counts[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output183 (.I(net183),
    .Z(all_counts[250]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output184 (.I(net184),
    .Z(all_counts[251]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output185 (.I(net185),
    .Z(all_counts[252]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output186 (.I(net186),
    .Z(all_counts[253]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output187 (.I(net187),
    .Z(all_counts[254]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output188 (.I(net188),
    .Z(all_counts[255]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output189 (.I(net189),
    .Z(all_counts[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output190 (.I(net190),
    .Z(all_counts[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output191 (.I(net191),
    .Z(all_counts[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output192 (.I(net192),
    .Z(all_counts[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output193 (.I(net193),
    .Z(all_counts[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output194 (.I(net194),
    .Z(all_counts[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output195 (.I(net195),
    .Z(all_counts[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output196 (.I(net196),
    .Z(all_counts[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output197 (.I(net197),
    .Z(all_counts[32]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output198 (.I(net198),
    .Z(all_counts[33]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output199 (.I(net199),
    .Z(all_counts[34]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output200 (.I(net200),
    .Z(all_counts[35]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output201 (.I(net201),
    .Z(all_counts[36]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output202 (.I(net202),
    .Z(all_counts[37]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output203 (.I(net203),
    .Z(all_counts[38]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output204 (.I(net204),
    .Z(all_counts[39]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output205 (.I(net205),
    .Z(all_counts[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output206 (.I(net206),
    .Z(all_counts[40]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output207 (.I(net207),
    .Z(all_counts[41]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output208 (.I(net208),
    .Z(all_counts[42]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output209 (.I(net209),
    .Z(all_counts[43]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output210 (.I(net210),
    .Z(all_counts[44]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output211 (.I(net211),
    .Z(all_counts[45]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output212 (.I(net212),
    .Z(all_counts[46]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output213 (.I(net213),
    .Z(all_counts[47]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output214 (.I(net214),
    .Z(all_counts[48]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output215 (.I(net215),
    .Z(all_counts[49]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output216 (.I(net216),
    .Z(all_counts[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output217 (.I(net217),
    .Z(all_counts[50]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output218 (.I(net218),
    .Z(all_counts[51]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output219 (.I(net219),
    .Z(all_counts[52]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output220 (.I(net220),
    .Z(all_counts[53]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output221 (.I(net221),
    .Z(all_counts[54]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output222 (.I(net222),
    .Z(all_counts[55]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output223 (.I(net223),
    .Z(all_counts[56]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output224 (.I(net224),
    .Z(all_counts[57]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output225 (.I(net225),
    .Z(all_counts[58]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output226 (.I(net226),
    .Z(all_counts[59]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output227 (.I(net227),
    .Z(all_counts[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output228 (.I(net228),
    .Z(all_counts[60]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output229 (.I(net229),
    .Z(all_counts[61]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output230 (.I(net230),
    .Z(all_counts[62]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output231 (.I(net231),
    .Z(all_counts[63]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output232 (.I(net232),
    .Z(all_counts[64]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output233 (.I(net233),
    .Z(all_counts[65]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output234 (.I(net234),
    .Z(all_counts[66]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output235 (.I(net235),
    .Z(all_counts[67]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output236 (.I(net236),
    .Z(all_counts[68]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output237 (.I(net237),
    .Z(all_counts[69]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output238 (.I(net238),
    .Z(all_counts[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output239 (.I(net239),
    .Z(all_counts[70]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output240 (.I(net240),
    .Z(all_counts[71]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output241 (.I(net241),
    .Z(all_counts[72]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output242 (.I(net242),
    .Z(all_counts[73]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output243 (.I(net243),
    .Z(all_counts[74]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output244 (.I(net244),
    .Z(all_counts[75]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output245 (.I(net245),
    .Z(all_counts[76]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output246 (.I(net246),
    .Z(all_counts[77]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output247 (.I(net247),
    .Z(all_counts[78]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output248 (.I(net248),
    .Z(all_counts[79]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output249 (.I(net249),
    .Z(all_counts[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output250 (.I(net250),
    .Z(all_counts[80]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output251 (.I(net251),
    .Z(all_counts[81]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output252 (.I(net252),
    .Z(all_counts[82]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output253 (.I(net253),
    .Z(all_counts[83]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output254 (.I(net254),
    .Z(all_counts[84]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output255 (.I(net255),
    .Z(all_counts[85]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output256 (.I(net256),
    .Z(all_counts[86]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output257 (.I(net257),
    .Z(all_counts[87]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output258 (.I(net258),
    .Z(all_counts[88]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output259 (.I(net259),
    .Z(all_counts[89]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output260 (.I(net260),
    .Z(all_counts[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output261 (.I(net261),
    .Z(all_counts[90]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output262 (.I(net262),
    .Z(all_counts[91]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output263 (.I(net263),
    .Z(all_counts[92]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output264 (.I(net264),
    .Z(all_counts[93]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output265 (.I(net265),
    .Z(all_counts[94]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output266 (.I(net266),
    .Z(all_counts[95]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output267 (.I(net267),
    .Z(all_counts[96]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output268 (.I(net268),
    .Z(all_counts[97]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output269 (.I(net269),
    .Z(all_counts[98]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output270 (.I(net270),
    .Z(all_counts[99]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output271 (.I(net271),
    .Z(all_counts[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output272 (.I(net272),
    .Z(count_value[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output273 (.I(net273),
    .Z(count_value[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output274 (.I(net274),
    .Z(count_value[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output275 (.I(net275),
    .Z(count_value[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output276 (.I(net276),
    .Z(count_value[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output277 (.I(net277),
    .Z(count_value[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output278 (.I(net278),
    .Z(count_value[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output279 (.I(net279),
    .Z(count_value[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output280 (.I(net280),
    .Z(count_value[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output281 (.I(net281),
    .Z(count_value[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output282 (.I(net282),
    .Z(count_value[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output283 (.I(net283),
    .Z(count_value[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output284 (.I(net284),
    .Z(count_value[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output285 (.I(net285),
    .Z(count_value[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output286 (.I(net286),
    .Z(count_value[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output287 (.I(net287),
    .Z(count_value[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output288 (.I(net288),
    .Z(count_value[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output289 (.I(net289),
    .Z(count_value[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output290 (.I(net290),
    .Z(count_value[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output291 (.I(net291),
    .Z(count_value[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output292 (.I(net292),
    .Z(count_value[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output293 (.I(net293),
    .Z(count_value[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output294 (.I(net294),
    .Z(count_value[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output295 (.I(net295),
    .Z(count_value[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output296 (.I(net296),
    .Z(count_value[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output297 (.I(net297),
    .Z(count_value[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output298 (.I(net298),
    .Z(count_value[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output299 (.I(net299),
    .Z(count_value[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output300 (.I(net300),
    .Z(count_value[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output301 (.I(net301),
    .Z(count_value[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output302 (.I(net302),
    .Z(count_value[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output303 (.I(net303),
    .Z(count_value[9]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_1_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_1_0__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload0 (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload1 (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload2 (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload3 (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload4 (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload5 (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload6 (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload7 (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload8 (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload9 (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload10 (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload11 (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold1 (.I(event_inc[2]),
    .Z(net304));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net305));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold3 (.I(event_inc[3]),
    .Z(net306));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold4 (.I(clear),
    .Z(net307));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(net16));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(net43));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_3 (.I(net155));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_4 (.I(net172));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_5 (.I(net281));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_6 (.I(net282));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_7 (.I(net285));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_8 (.I(net297));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_9 (.I(net279));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_777 ();
endmodule
