module pipelined_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    rd_en,
    rst_n,
    wr_en,
    data_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input rd_en;
 input rst_n;
 input wr_en;
 output [4:0] data_count;
 output [31:0] rd_data;
 input [31:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire clknet_0_clk;
 wire \pipeline_count[0] ;
 wire \pipeline_count[1] ;
 wire \pipeline_count[2] ;
 wire \pipeline_count[3] ;
 wire \pipeline_count[4] ;
 wire rd_en_pipe;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_en_pipe[0] ;
 wire \wr_en_pipe[1] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _166_ (.A(_125_),
    .ZN(_130_));
 INV_X1 _167_ (.A(_137_),
    .ZN(_164_));
 BUF_X2 _168_ (.A(_162_),
    .Z(_105_));
 XNOR2_X2 _169_ (.A(_105_),
    .B(_124_),
    .ZN(_106_));
 INV_X1 _170_ (.A(_106_),
    .ZN(_143_));
 BUF_X4 _171_ (.A(_159_),
    .Z(_107_));
 INV_X1 _172_ (.A(_107_),
    .ZN(_108_));
 INV_X1 _173_ (.A(_136_),
    .ZN(_123_));
 NAND3_X2 _174_ (.A1(_105_),
    .A2(_123_),
    .A3(_135_),
    .ZN(_109_));
 AOI21_X4 _175_ (.A(_161_),
    .B1(_163_),
    .B2(_105_),
    .ZN(_110_));
 AOI21_X4 _176_ (.A(_108_),
    .B1(_109_),
    .B2(_110_),
    .ZN(_111_));
 AND3_X1 _177_ (.A1(_105_),
    .A2(_123_),
    .A3(_135_),
    .ZN(_023_));
 INV_X1 _178_ (.A(_110_),
    .ZN(_024_));
 NOR3_X4 _179_ (.A1(_107_),
    .A2(_023_),
    .A3(_024_),
    .ZN(_025_));
 NOR2_X2 _180_ (.A1(_111_),
    .A2(_025_),
    .ZN(_146_));
 OR4_X1 _181_ (.A1(\pipeline_count[1] ),
    .A2(\pipeline_count[3] ),
    .A3(\pipeline_count[2] ),
    .A4(\pipeline_count[4] ),
    .ZN(_026_));
 AND2_X1 _182_ (.A1(_107_),
    .A2(_105_),
    .ZN(_027_));
 AOI221_X2 _183_ (.A(_158_),
    .B1(_161_),
    .B2(_107_),
    .C1(_027_),
    .C2(_124_),
    .ZN(_028_));
 XNOR2_X2 _184_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .ZN(_029_));
 XOR2_X2 _185_ (.A(_028_),
    .B(_029_),
    .Z(_030_));
 NOR3_X1 _186_ (.A1(_125_),
    .A2(_164_),
    .A3(\pipeline_count[0] ),
    .ZN(_031_));
 NAND3_X1 _187_ (.A1(_106_),
    .A2(_030_),
    .A3(_031_),
    .ZN(_032_));
 NOR3_X1 _188_ (.A1(_146_),
    .A2(_026_),
    .A3(_032_),
    .ZN(net11));
 NAND2_X2 _189_ (.A1(_125_),
    .A2(_143_),
    .ZN(_033_));
 OR3_X2 _190_ (.A1(_111_),
    .A2(_025_),
    .A3(_033_),
    .ZN(_034_));
 NAND2_X1 _191_ (.A1(_030_),
    .A2(_034_),
    .ZN(net12));
 INV_X1 _192_ (.A(_134_),
    .ZN(_131_));
 INV_X1 _193_ (.A(_133_),
    .ZN(net7));
 INV_X2 _194_ (.A(_139_),
    .ZN(_126_));
 BUF_X2 _195_ (.A(net2),
    .Z(_035_));
 BUF_X2 _196_ (.A(_140_),
    .Z(_036_));
 MUX2_X1 _197_ (.A(_002_),
    .B(\pipeline_count[0] ),
    .S(_036_),
    .Z(_037_));
 AND2_X1 _198_ (.A1(_035_),
    .A2(_037_),
    .ZN(_005_));
 INV_X1 _199_ (.A(net2),
    .ZN(_038_));
 CLKBUF_X3 _200_ (.A(_038_),
    .Z(_039_));
 NOR2_X1 _201_ (.A1(_128_),
    .A2(_036_),
    .ZN(_040_));
 AOI21_X1 _202_ (.A(_040_),
    .B1(_036_),
    .B2(\pipeline_count[1] ),
    .ZN(_041_));
 NOR2_X1 _203_ (.A1(_039_),
    .A2(_041_),
    .ZN(_006_));
 XOR2_X1 _204_ (.A(_127_),
    .B(_154_),
    .Z(_042_));
 MUX2_X1 _205_ (.A(_042_),
    .B(\pipeline_count[2] ),
    .S(_036_),
    .Z(_043_));
 AND2_X1 _206_ (.A1(_035_),
    .A2(_043_),
    .ZN(_007_));
 AOI21_X1 _207_ (.A(_151_),
    .B1(_152_),
    .B2(\pipeline_count[0] ),
    .ZN(_044_));
 INV_X1 _208_ (.A(_044_),
    .ZN(_045_));
 AOI21_X1 _209_ (.A(_153_),
    .B1(_045_),
    .B2(_154_),
    .ZN(_046_));
 XNOR2_X1 _210_ (.A(_156_),
    .B(_046_),
    .ZN(_047_));
 MUX2_X1 _211_ (.A(_047_),
    .B(\pipeline_count[3] ),
    .S(_036_),
    .Z(_048_));
 AND2_X1 _212_ (.A1(_035_),
    .A2(_048_),
    .ZN(_008_));
 INV_X1 _213_ (.A(_155_),
    .ZN(_049_));
 AOI21_X1 _214_ (.A(_153_),
    .B1(_154_),
    .B2(_127_),
    .ZN(_050_));
 INV_X1 _215_ (.A(_156_),
    .ZN(_051_));
 OAI21_X1 _216_ (.A(_049_),
    .B1(_050_),
    .B2(_051_),
    .ZN(_052_));
 XNOR2_X1 _217_ (.A(_126_),
    .B(_052_),
    .ZN(_053_));
 NOR2_X1 _218_ (.A1(_036_),
    .A2(_053_),
    .ZN(_054_));
 XNOR2_X1 _219_ (.A(\pipeline_count[4] ),
    .B(_054_),
    .ZN(_055_));
 NOR2_X1 _220_ (.A1(_039_),
    .A2(_055_),
    .ZN(_009_));
 INV_X1 _221_ (.A(net1),
    .ZN(_056_));
 XNOR2_X1 _222_ (.A(_028_),
    .B(_029_),
    .ZN(_057_));
 NOR2_X1 _223_ (.A1(_143_),
    .A2(_026_),
    .ZN(_058_));
 NAND2_X1 _224_ (.A1(_031_),
    .A2(_058_),
    .ZN(_059_));
 OAI21_X1 _225_ (.A(_107_),
    .B1(_023_),
    .B2(_024_),
    .ZN(_060_));
 NAND3_X1 _226_ (.A1(_108_),
    .A2(_109_),
    .A3(_110_),
    .ZN(_061_));
 AOI211_X4 _227_ (.A(_057_),
    .B(_059_),
    .C1(_060_),
    .C2(_061_),
    .ZN(_062_));
 NOR3_X1 _228_ (.A1(_056_),
    .A2(_039_),
    .A3(_062_),
    .ZN(_010_));
 AND2_X1 _229_ (.A1(\rd_ptr[0] ),
    .A2(_035_),
    .ZN(_063_));
 AND2_X1 _230_ (.A1(_000_),
    .A2(_035_),
    .ZN(_064_));
 NOR2_X1 _231_ (.A1(_056_),
    .A2(_062_),
    .ZN(_065_));
 MUX2_X1 _232_ (.A(_063_),
    .B(_064_),
    .S(_065_),
    .Z(_011_));
 AND2_X1 _233_ (.A1(\rd_ptr[1] ),
    .A2(_035_),
    .ZN(_066_));
 AND2_X1 _234_ (.A1(_001_),
    .A2(_035_),
    .ZN(_067_));
 MUX2_X1 _235_ (.A(_066_),
    .B(_067_),
    .S(_065_),
    .Z(_012_));
 NAND2_X1 _236_ (.A1(net1),
    .A2(_150_),
    .ZN(_068_));
 OAI21_X1 _237_ (.A(\rd_ptr[2] ),
    .B1(_062_),
    .B2(_068_),
    .ZN(_069_));
 OR3_X1 _238_ (.A1(\rd_ptr[2] ),
    .A2(_062_),
    .A3(_068_),
    .ZN(_070_));
 AOI21_X1 _239_ (.A(_039_),
    .B1(_069_),
    .B2(_070_),
    .ZN(_013_));
 AND2_X1 _240_ (.A1(\rd_ptr[3] ),
    .A2(_035_),
    .ZN(_071_));
 NOR2_X1 _241_ (.A1(\rd_ptr[3] ),
    .A2(_039_),
    .ZN(_072_));
 NAND3_X1 _242_ (.A1(\rd_ptr[2] ),
    .A2(\rd_ptr[1] ),
    .A3(\rd_ptr[0] ),
    .ZN(_073_));
 NOR3_X1 _243_ (.A1(_056_),
    .A2(_062_),
    .A3(_073_),
    .ZN(_074_));
 MUX2_X1 _244_ (.A(_071_),
    .B(_072_),
    .S(_074_),
    .Z(_014_));
 NAND4_X1 _245_ (.A1(net1),
    .A2(_150_),
    .A3(\rd_ptr[2] ),
    .A4(\rd_ptr[3] ),
    .ZN(_075_));
 OAI21_X1 _246_ (.A(\rd_ptr[4] ),
    .B1(_062_),
    .B2(_075_),
    .ZN(_076_));
 OR3_X1 _247_ (.A1(\rd_ptr[4] ),
    .A2(_062_),
    .A3(_075_),
    .ZN(_077_));
 AOI21_X1 _248_ (.A(_039_),
    .B1(_076_),
    .B2(_077_),
    .ZN(_015_));
 NOR3_X4 _249_ (.A1(_111_),
    .A2(_025_),
    .A3(_033_),
    .ZN(_078_));
 NAND2_X2 _250_ (.A1(net3),
    .A2(_030_),
    .ZN(_079_));
 NOR3_X1 _251_ (.A1(_039_),
    .A2(_078_),
    .A3(_079_),
    .ZN(_016_));
 AND2_X1 _252_ (.A1(_035_),
    .A2(\wr_en_pipe[0] ),
    .ZN(_017_));
 AND2_X1 _253_ (.A1(net3),
    .A2(_030_),
    .ZN(_080_));
 NAND3_X1 _254_ (.A1(_003_),
    .A2(_034_),
    .A3(_080_),
    .ZN(_081_));
 OAI21_X1 _255_ (.A(\wr_ptr[0] ),
    .B1(_078_),
    .B2(_079_),
    .ZN(_082_));
 AOI21_X1 _256_ (.A(_039_),
    .B1(_081_),
    .B2(_082_),
    .ZN(_018_));
 NAND3_X1 _257_ (.A1(_004_),
    .A2(_034_),
    .A3(_080_),
    .ZN(_083_));
 OAI21_X1 _258_ (.A(\wr_ptr[1] ),
    .B1(_078_),
    .B2(_079_),
    .ZN(_084_));
 AOI21_X1 _259_ (.A(_039_),
    .B1(_083_),
    .B2(_084_),
    .ZN(_019_));
 NOR2_X1 _260_ (.A1(\wr_ptr[2] ),
    .A2(_038_),
    .ZN(_085_));
 AND2_X1 _261_ (.A1(\wr_ptr[2] ),
    .A2(_035_),
    .ZN(_086_));
 NAND3_X1 _262_ (.A1(_149_),
    .A2(_034_),
    .A3(_080_),
    .ZN(_087_));
 MUX2_X1 _263_ (.A(_085_),
    .B(_086_),
    .S(_087_),
    .Z(_020_));
 AND2_X1 _264_ (.A1(\wr_ptr[3] ),
    .A2(net2),
    .ZN(_088_));
 NOR2_X1 _265_ (.A1(\wr_ptr[3] ),
    .A2(_039_),
    .ZN(_089_));
 NAND3_X1 _266_ (.A1(\wr_ptr[2] ),
    .A2(\wr_ptr[1] ),
    .A3(\wr_ptr[0] ),
    .ZN(_090_));
 NOR3_X1 _267_ (.A1(_078_),
    .A2(_079_),
    .A3(_090_),
    .ZN(_091_));
 MUX2_X1 _268_ (.A(_088_),
    .B(_089_),
    .S(_091_),
    .Z(_021_));
 AND2_X1 _269_ (.A1(\wr_ptr[4] ),
    .A2(net2),
    .ZN(_092_));
 NOR2_X1 _270_ (.A1(\wr_ptr[4] ),
    .A2(_038_),
    .ZN(_093_));
 NAND3_X1 _271_ (.A1(_149_),
    .A2(\wr_ptr[2] ),
    .A3(\wr_ptr[3] ),
    .ZN(_094_));
 NOR3_X1 _272_ (.A1(_078_),
    .A2(_079_),
    .A3(_094_),
    .ZN(_095_));
 MUX2_X1 _273_ (.A(_092_),
    .B(_093_),
    .S(_095_),
    .Z(_022_));
 AOI21_X1 _274_ (.A(_106_),
    .B1(_137_),
    .B2(_130_),
    .ZN(_096_));
 NOR4_X1 _275_ (.A1(_146_),
    .A2(_026_),
    .A3(_057_),
    .A4(_096_),
    .ZN(net4));
 NAND2_X1 _276_ (.A1(_143_),
    .A2(_146_),
    .ZN(_097_));
 NAND2_X1 _277_ (.A1(_030_),
    .A2(_097_),
    .ZN(net5));
 XNOR2_X1 _278_ (.A(_145_),
    .B(_132_),
    .ZN(net8));
 INV_X1 _279_ (.A(_144_),
    .ZN(_098_));
 AOI21_X1 _280_ (.A(_141_),
    .B1(_134_),
    .B2(_142_),
    .ZN(_099_));
 INV_X1 _281_ (.A(_145_),
    .ZN(_100_));
 OAI21_X1 _282_ (.A(_098_),
    .B1(_099_),
    .B2(_100_),
    .ZN(_101_));
 XOR2_X1 _283_ (.A(_148_),
    .B(_101_),
    .Z(net9));
 OAI21_X1 _284_ (.A(_098_),
    .B1(_132_),
    .B2(_100_),
    .ZN(_102_));
 AOI21_X1 _285_ (.A(_147_),
    .B1(_102_),
    .B2(_148_),
    .ZN(_103_));
 XNOR2_X1 _286_ (.A(\pipeline_count[4] ),
    .B(_103_),
    .ZN(_104_));
 XNOR2_X1 _287_ (.A(_030_),
    .B(_104_),
    .ZN(net10));
 FA_X1 _288_ (.A(_122_),
    .B(\wr_ptr[1] ),
    .CI(_123_),
    .CO(_124_),
    .S(_125_));
 FA_X1 _289_ (.A(\pipeline_count[0] ),
    .B(\pipeline_count[1] ),
    .CI(_126_),
    .CO(_127_),
    .S(_128_));
 FA_X1 _290_ (.A(_129_),
    .B(_130_),
    .CI(_131_),
    .CO(_132_),
    .S(_133_));
 HA_X1 _291_ (.A(\rd_ptr[0] ),
    .B(_003_),
    .CO(_136_),
    .S(_137_));
 HA_X1 _292_ (.A(_138_),
    .B(\wr_en_pipe[1] ),
    .CO(_139_),
    .S(_140_));
 HA_X1 _293_ (.A(\pipeline_count[1] ),
    .B(_125_),
    .CO(_141_),
    .S(_142_));
 HA_X1 _294_ (.A(\pipeline_count[2] ),
    .B(_143_),
    .CO(_144_),
    .S(_145_));
 HA_X1 _295_ (.A(\pipeline_count[3] ),
    .B(_146_),
    .CO(_147_),
    .S(_148_));
 HA_X1 _296_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .CO(_149_),
    .S(_004_));
 HA_X1 _297_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .CO(_150_),
    .S(_001_));
 HA_X1 _298_ (.A(\pipeline_count[1] ),
    .B(_126_),
    .CO(_151_),
    .S(_152_));
 HA_X1 _299_ (.A(\pipeline_count[2] ),
    .B(_126_),
    .CO(_153_),
    .S(_154_));
 HA_X1 _300_ (.A(\pipeline_count[3] ),
    .B(_126_),
    .CO(_155_),
    .S(_156_));
 HA_X1 _301_ (.A(_157_),
    .B(\wr_ptr[3] ),
    .CO(_158_),
    .S(_159_));
 HA_X1 _302_ (.A(_160_),
    .B(\wr_ptr[2] ),
    .CO(_161_),
    .S(_162_));
 HA_X1 _303_ (.A(_122_),
    .B(\wr_ptr[1] ),
    .CO(_163_),
    .S(_135_));
 HA_X1 _304_ (.A(\pipeline_count[0] ),
    .B(_164_),
    .CO(_134_),
    .S(net6));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X1 _306_ (.A(net13),
    .Z(rd_data[0]));
 BUF_X1 _307_ (.A(net14),
    .Z(rd_data[1]));
 BUF_X1 _308_ (.A(net15),
    .Z(rd_data[2]));
 BUF_X1 _309_ (.A(net16),
    .Z(rd_data[3]));
 BUF_X1 _310_ (.A(net17),
    .Z(rd_data[4]));
 BUF_X1 _311_ (.A(net18),
    .Z(rd_data[5]));
 BUF_X1 _312_ (.A(net19),
    .Z(rd_data[6]));
 BUF_X1 _313_ (.A(net20),
    .Z(rd_data[7]));
 BUF_X1 _314_ (.A(net21),
    .Z(rd_data[8]));
 BUF_X1 _315_ (.A(net22),
    .Z(rd_data[9]));
 BUF_X1 _316_ (.A(net23),
    .Z(rd_data[10]));
 BUF_X1 _317_ (.A(net24),
    .Z(rd_data[11]));
 BUF_X1 _318_ (.A(net25),
    .Z(rd_data[12]));
 BUF_X1 _319_ (.A(net26),
    .Z(rd_data[13]));
 BUF_X1 _320_ (.A(net27),
    .Z(rd_data[14]));
 BUF_X1 _321_ (.A(net28),
    .Z(rd_data[15]));
 BUF_X1 _322_ (.A(net29),
    .Z(rd_data[16]));
 BUF_X1 _323_ (.A(net30),
    .Z(rd_data[17]));
 BUF_X1 _324_ (.A(net31),
    .Z(rd_data[18]));
 BUF_X1 _325_ (.A(net32),
    .Z(rd_data[19]));
 BUF_X1 _326_ (.A(net33),
    .Z(rd_data[20]));
 BUF_X1 _327_ (.A(net34),
    .Z(rd_data[21]));
 BUF_X1 _328_ (.A(net35),
    .Z(rd_data[22]));
 BUF_X1 _329_ (.A(net36),
    .Z(rd_data[23]));
 BUF_X1 _330_ (.A(net37),
    .Z(rd_data[24]));
 BUF_X1 _331_ (.A(net38),
    .Z(rd_data[25]));
 BUF_X1 _332_ (.A(net39),
    .Z(rd_data[26]));
 BUF_X1 _333_ (.A(net40),
    .Z(rd_data[27]));
 BUF_X1 _334_ (.A(net41),
    .Z(rd_data[28]));
 BUF_X1 _335_ (.A(net42),
    .Z(rd_data[29]));
 BUF_X1 _336_ (.A(net43),
    .Z(rd_data[30]));
 BUF_X1 _337_ (.A(net44),
    .Z(rd_data[31]));
 DFF_X2 \pipeline_count[0]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\pipeline_count[0] ),
    .QN(_002_));
 DFF_X2 \pipeline_count[1]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\pipeline_count[1] ),
    .QN(_129_));
 DFF_X2 \pipeline_count[2]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\pipeline_count[2] ),
    .QN(_121_));
 DFF_X2 \pipeline_count[3]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\pipeline_count[3] ),
    .QN(_120_));
 DFF_X1 \pipeline_count[4]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\pipeline_count[4] ),
    .QN(_119_));
 DFF_X1 \rd_en_pipe$_SDFF_PN0_  (.D(_010_),
    .CK(clknet_1_1__leaf_clk),
    .Q(rd_en_pipe),
    .QN(_138_));
 DFF_X2 \rd_ptr[0]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\rd_ptr[0] ),
    .QN(_000_));
 DFF_X1 \rd_ptr[1]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\rd_ptr[1] ),
    .QN(_122_));
 DFF_X1 \rd_ptr[2]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\rd_ptr[2] ),
    .QN(_160_));
 DFF_X1 \rd_ptr[3]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\rd_ptr[3] ),
    .QN(_157_));
 DFF_X1 \rd_ptr[4]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\rd_ptr[4] ),
    .QN(_118_));
 DFF_X1 \wr_en_pipe[0]$_SDFF_PN0_  (.D(_016_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\wr_en_pipe[0] ),
    .QN(_117_));
 DFF_X1 \wr_en_pipe[1]$_SDFF_PN0_  (.D(_017_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\wr_en_pipe[1] ),
    .QN(_116_));
 DFF_X1 \wr_ptr[0]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\wr_ptr[0] ),
    .QN(_003_));
 DFF_X2 \wr_ptr[1]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\wr_ptr[1] ),
    .QN(_115_));
 DFF_X2 \wr_ptr[2]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\wr_ptr[2] ),
    .QN(_114_));
 DFF_X2 \wr_ptr[3]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\wr_ptr[3] ),
    .QN(_113_));
 DFF_X1 \wr_ptr[4]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\wr_ptr[4] ),
    .QN(_112_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_75 ();
 BUF_X1 input1 (.A(rd_en),
    .Z(net1));
 BUF_X1 input2 (.A(rst_n),
    .Z(net2));
 BUF_X1 input3 (.A(wr_en),
    .Z(net3));
 BUF_X1 output4 (.A(net4),
    .Z(almost_empty));
 BUF_X1 output5 (.A(net5),
    .Z(almost_full));
 BUF_X1 output6 (.A(net6),
    .Z(data_count[0]));
 BUF_X1 output7 (.A(net7),
    .Z(data_count[1]));
 BUF_X1 output8 (.A(net8),
    .Z(data_count[2]));
 BUF_X1 output9 (.A(net9),
    .Z(data_count[3]));
 BUF_X1 output10 (.A(net10),
    .Z(data_count[4]));
 BUF_X1 output11 (.A(net11),
    .Z(empty));
 BUF_X1 output12 (.A(net12),
    .Z(full));
 LOGIC0_X1 _306__13 (.Z(net13));
 LOGIC0_X1 _307__14 (.Z(net14));
 LOGIC0_X1 _308__15 (.Z(net15));
 LOGIC0_X1 _309__16 (.Z(net16));
 LOGIC0_X1 _310__17 (.Z(net17));
 LOGIC0_X1 _311__18 (.Z(net18));
 LOGIC0_X1 _312__19 (.Z(net19));
 LOGIC0_X1 _313__20 (.Z(net20));
 LOGIC0_X1 _314__21 (.Z(net21));
 LOGIC0_X1 _315__22 (.Z(net22));
 LOGIC0_X1 _316__23 (.Z(net23));
 LOGIC0_X1 _317__24 (.Z(net24));
 LOGIC0_X1 _318__25 (.Z(net25));
 LOGIC0_X1 _319__26 (.Z(net26));
 LOGIC0_X1 _320__27 (.Z(net27));
 LOGIC0_X1 _321__28 (.Z(net28));
 LOGIC0_X1 _322__29 (.Z(net29));
 LOGIC0_X1 _323__30 (.Z(net30));
 LOGIC0_X1 _324__31 (.Z(net31));
 LOGIC0_X1 _325__32 (.Z(net32));
 LOGIC0_X1 _326__33 (.Z(net33));
 LOGIC0_X1 _327__34 (.Z(net34));
 LOGIC0_X1 _328__35 (.Z(net35));
 LOGIC0_X1 _329__36 (.Z(net36));
 LOGIC0_X1 _330__37 (.Z(net37));
 LOGIC0_X1 _331__38 (.Z(net38));
 LOGIC0_X1 _332__39 (.Z(net39));
 LOGIC0_X1 _333__40 (.Z(net40));
 LOGIC0_X1 _334__41 (.Z(net41));
 LOGIC0_X1 _335__42 (.Z(net42));
 LOGIC0_X1 _336__43 (.Z(net43));
 LOGIC0_X1 _337__44 (.Z(net44));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 INV_X1 clkload0 (.A(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_97 ();
 FILLCELL_X2 FILLER_0_101 ();
 FILLCELL_X1 FILLER_0_103 ();
 FILLCELL_X32 FILLER_0_107 ();
 FILLCELL_X8 FILLER_0_139 ();
 FILLCELL_X4 FILLER_0_147 ();
 FILLCELL_X32 FILLER_0_154 ();
 FILLCELL_X32 FILLER_0_186 ();
 FILLCELL_X32 FILLER_0_218 ();
 FILLCELL_X32 FILLER_0_250 ();
 FILLCELL_X2 FILLER_0_282 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X16 FILLER_1_129 ();
 FILLCELL_X4 FILLER_1_145 ();
 FILLCELL_X32 FILLER_1_152 ();
 FILLCELL_X32 FILLER_1_184 ();
 FILLCELL_X32 FILLER_1_216 ();
 FILLCELL_X32 FILLER_1_248 ();
 FILLCELL_X4 FILLER_1_280 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X16 FILLER_2_257 ();
 FILLCELL_X8 FILLER_2_273 ();
 FILLCELL_X2 FILLER_2_281 ();
 FILLCELL_X1 FILLER_2_283 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X16 FILLER_3_257 ();
 FILLCELL_X8 FILLER_3_273 ();
 FILLCELL_X2 FILLER_3_281 ();
 FILLCELL_X1 FILLER_3_283 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X16 FILLER_4_257 ();
 FILLCELL_X8 FILLER_4_273 ();
 FILLCELL_X2 FILLER_4_281 ();
 FILLCELL_X1 FILLER_4_283 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X16 FILLER_5_257 ();
 FILLCELL_X8 FILLER_5_273 ();
 FILLCELL_X2 FILLER_5_281 ();
 FILLCELL_X1 FILLER_5_283 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X16 FILLER_6_257 ();
 FILLCELL_X8 FILLER_6_273 ();
 FILLCELL_X2 FILLER_6_281 ();
 FILLCELL_X1 FILLER_6_283 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X16 FILLER_7_257 ();
 FILLCELL_X8 FILLER_7_273 ();
 FILLCELL_X2 FILLER_7_281 ();
 FILLCELL_X1 FILLER_7_283 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X16 FILLER_8_257 ();
 FILLCELL_X8 FILLER_8_273 ();
 FILLCELL_X2 FILLER_8_281 ();
 FILLCELL_X1 FILLER_8_283 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X16 FILLER_9_257 ();
 FILLCELL_X8 FILLER_9_273 ();
 FILLCELL_X2 FILLER_9_281 ();
 FILLCELL_X1 FILLER_9_283 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X16 FILLER_10_257 ();
 FILLCELL_X8 FILLER_10_273 ();
 FILLCELL_X2 FILLER_10_281 ();
 FILLCELL_X1 FILLER_10_283 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X16 FILLER_11_257 ();
 FILLCELL_X4 FILLER_11_273 ();
 FILLCELL_X1 FILLER_11_277 ();
 FILLCELL_X1 FILLER_11_283 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X8 FILLER_12_257 ();
 FILLCELL_X4 FILLER_12_265 ();
 FILLCELL_X2 FILLER_12_269 ();
 FILLCELL_X1 FILLER_12_271 ();
 FILLCELL_X2 FILLER_12_277 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X8 FILLER_13_257 ();
 FILLCELL_X4 FILLER_13_265 ();
 FILLCELL_X1 FILLER_13_276 ();
 FILLCELL_X1 FILLER_13_280 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X2 FILLER_14_97 ();
 FILLCELL_X8 FILLER_14_103 ();
 FILLCELL_X4 FILLER_14_111 ();
 FILLCELL_X2 FILLER_14_115 ();
 FILLCELL_X8 FILLER_14_136 ();
 FILLCELL_X4 FILLER_14_144 ();
 FILLCELL_X1 FILLER_14_148 ();
 FILLCELL_X32 FILLER_14_152 ();
 FILLCELL_X32 FILLER_14_184 ();
 FILLCELL_X32 FILLER_14_216 ();
 FILLCELL_X16 FILLER_14_248 ();
 FILLCELL_X4 FILLER_14_264 ();
 FILLCELL_X1 FILLER_14_268 ();
 FILLCELL_X2 FILLER_14_271 ();
 FILLCELL_X1 FILLER_14_273 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X16 FILLER_15_65 ();
 FILLCELL_X8 FILLER_15_81 ();
 FILLCELL_X4 FILLER_15_89 ();
 FILLCELL_X1 FILLER_15_93 ();
 FILLCELL_X4 FILLER_15_101 ();
 FILLCELL_X2 FILLER_15_105 ();
 FILLCELL_X1 FILLER_15_107 ();
 FILLCELL_X1 FILLER_15_111 ();
 FILLCELL_X1 FILLER_15_119 ();
 FILLCELL_X16 FILLER_15_124 ();
 FILLCELL_X4 FILLER_15_140 ();
 FILLCELL_X2 FILLER_15_144 ();
 FILLCELL_X32 FILLER_15_155 ();
 FILLCELL_X32 FILLER_15_187 ();
 FILLCELL_X32 FILLER_15_219 ();
 FILLCELL_X16 FILLER_15_251 ();
 FILLCELL_X2 FILLER_15_267 ();
 FILLCELL_X1 FILLER_15_276 ();
 FILLCELL_X1 FILLER_15_280 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X1 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_37 ();
 FILLCELL_X8 FILLER_16_69 ();
 FILLCELL_X2 FILLER_16_77 ();
 FILLCELL_X8 FILLER_16_114 ();
 FILLCELL_X4 FILLER_16_122 ();
 FILLCELL_X1 FILLER_16_126 ();
 FILLCELL_X1 FILLER_16_131 ();
 FILLCELL_X1 FILLER_16_136 ();
 FILLCELL_X1 FILLER_16_147 ();
 FILLCELL_X1 FILLER_16_152 ();
 FILLCELL_X1 FILLER_16_157 ();
 FILLCELL_X1 FILLER_16_162 ();
 FILLCELL_X1 FILLER_16_167 ();
 FILLCELL_X32 FILLER_16_187 ();
 FILLCELL_X32 FILLER_16_219 ();
 FILLCELL_X16 FILLER_16_251 ();
 FILLCELL_X4 FILLER_16_267 ();
 FILLCELL_X1 FILLER_16_271 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X8 FILLER_17_97 ();
 FILLCELL_X2 FILLER_17_105 ();
 FILLCELL_X8 FILLER_17_114 ();
 FILLCELL_X4 FILLER_17_122 ();
 FILLCELL_X2 FILLER_17_126 ();
 FILLCELL_X1 FILLER_17_128 ();
 FILLCELL_X32 FILLER_17_137 ();
 FILLCELL_X32 FILLER_17_169 ();
 FILLCELL_X32 FILLER_17_201 ();
 FILLCELL_X32 FILLER_17_233 ();
 FILLCELL_X4 FILLER_17_265 ();
 FILLCELL_X1 FILLER_17_279 ();
 FILLCELL_X1 FILLER_17_283 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X4 FILLER_18_97 ();
 FILLCELL_X4 FILLER_18_120 ();
 FILLCELL_X4 FILLER_18_153 ();
 FILLCELL_X1 FILLER_18_157 ();
 FILLCELL_X1 FILLER_18_162 ();
 FILLCELL_X32 FILLER_18_184 ();
 FILLCELL_X32 FILLER_18_216 ();
 FILLCELL_X16 FILLER_18_248 ();
 FILLCELL_X4 FILLER_18_264 ();
 FILLCELL_X1 FILLER_18_268 ();
 FILLCELL_X2 FILLER_18_271 ();
 FILLCELL_X1 FILLER_18_273 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X8 FILLER_19_65 ();
 FILLCELL_X2 FILLER_19_73 ();
 FILLCELL_X1 FILLER_19_75 ();
 FILLCELL_X1 FILLER_19_85 ();
 FILLCELL_X16 FILLER_19_90 ();
 FILLCELL_X4 FILLER_19_106 ();
 FILLCELL_X32 FILLER_19_113 ();
 FILLCELL_X32 FILLER_19_145 ();
 FILLCELL_X2 FILLER_19_177 ();
 FILLCELL_X1 FILLER_19_179 ();
 FILLCELL_X32 FILLER_19_197 ();
 FILLCELL_X32 FILLER_19_229 ();
 FILLCELL_X8 FILLER_19_261 ();
 FILLCELL_X1 FILLER_19_274 ();
 FILLCELL_X1 FILLER_19_280 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X8 FILLER_20_65 ();
 FILLCELL_X1 FILLER_20_73 ();
 FILLCELL_X1 FILLER_20_91 ();
 FILLCELL_X16 FILLER_20_102 ();
 FILLCELL_X8 FILLER_20_118 ();
 FILLCELL_X32 FILLER_20_131 ();
 FILLCELL_X32 FILLER_20_163 ();
 FILLCELL_X32 FILLER_20_195 ();
 FILLCELL_X32 FILLER_20_227 ();
 FILLCELL_X8 FILLER_20_259 ();
 FILLCELL_X4 FILLER_20_267 ();
 FILLCELL_X1 FILLER_20_273 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X16 FILLER_21_65 ();
 FILLCELL_X4 FILLER_21_81 ();
 FILLCELL_X4 FILLER_21_102 ();
 FILLCELL_X2 FILLER_21_106 ();
 FILLCELL_X1 FILLER_21_108 ();
 FILLCELL_X4 FILLER_21_119 ();
 FILLCELL_X1 FILLER_21_123 ();
 FILLCELL_X32 FILLER_21_133 ();
 FILLCELL_X32 FILLER_21_165 ();
 FILLCELL_X32 FILLER_21_197 ();
 FILLCELL_X32 FILLER_21_229 ();
 FILLCELL_X8 FILLER_21_261 ();
 FILLCELL_X1 FILLER_21_276 ();
 FILLCELL_X1 FILLER_21_283 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X1 FILLER_22_65 ();
 FILLCELL_X1 FILLER_22_69 ();
 FILLCELL_X2 FILLER_22_83 ();
 FILLCELL_X16 FILLER_22_88 ();
 FILLCELL_X8 FILLER_22_104 ();
 FILLCELL_X2 FILLER_22_112 ();
 FILLCELL_X1 FILLER_22_114 ();
 FILLCELL_X2 FILLER_22_122 ();
 FILLCELL_X32 FILLER_22_150 ();
 FILLCELL_X8 FILLER_22_182 ();
 FILLCELL_X4 FILLER_22_190 ();
 FILLCELL_X32 FILLER_22_204 ();
 FILLCELL_X32 FILLER_22_236 ();
 FILLCELL_X4 FILLER_22_268 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X1 FILLER_23_65 ();
 FILLCELL_X1 FILLER_23_71 ();
 FILLCELL_X2 FILLER_23_76 ();
 FILLCELL_X1 FILLER_23_80 ();
 FILLCELL_X8 FILLER_23_88 ();
 FILLCELL_X2 FILLER_23_96 ();
 FILLCELL_X1 FILLER_23_98 ();
 FILLCELL_X4 FILLER_23_103 ();
 FILLCELL_X2 FILLER_23_136 ();
 FILLCELL_X1 FILLER_23_138 ();
 FILLCELL_X8 FILLER_23_157 ();
 FILLCELL_X2 FILLER_23_165 ();
 FILLCELL_X1 FILLER_23_167 ();
 FILLCELL_X4 FILLER_23_189 ();
 FILLCELL_X2 FILLER_23_193 ();
 FILLCELL_X1 FILLER_23_195 ();
 FILLCELL_X32 FILLER_23_200 ();
 FILLCELL_X32 FILLER_23_232 ();
 FILLCELL_X2 FILLER_23_264 ();
 FILLCELL_X1 FILLER_23_266 ();
 FILLCELL_X1 FILLER_23_279 ();
 FILLCELL_X1 FILLER_23_283 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X2 FILLER_24_65 ();
 FILLCELL_X1 FILLER_24_84 ();
 FILLCELL_X32 FILLER_24_89 ();
 FILLCELL_X4 FILLER_24_121 ();
 FILLCELL_X2 FILLER_24_125 ();
 FILLCELL_X1 FILLER_24_127 ();
 FILLCELL_X1 FILLER_24_141 ();
 FILLCELL_X1 FILLER_24_144 ();
 FILLCELL_X32 FILLER_24_151 ();
 FILLCELL_X1 FILLER_24_183 ();
 FILLCELL_X32 FILLER_24_206 ();
 FILLCELL_X32 FILLER_24_238 ();
 FILLCELL_X8 FILLER_24_270 ();
 FILLCELL_X1 FILLER_24_278 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X8 FILLER_25_65 ();
 FILLCELL_X4 FILLER_25_73 ();
 FILLCELL_X1 FILLER_25_77 ();
 FILLCELL_X32 FILLER_25_85 ();
 FILLCELL_X4 FILLER_25_117 ();
 FILLCELL_X2 FILLER_25_121 ();
 FILLCELL_X32 FILLER_25_157 ();
 FILLCELL_X4 FILLER_25_189 ();
 FILLCELL_X2 FILLER_25_193 ();
 FILLCELL_X1 FILLER_25_195 ();
 FILLCELL_X32 FILLER_25_203 ();
 FILLCELL_X32 FILLER_25_235 ();
 FILLCELL_X16 FILLER_25_267 ();
 FILLCELL_X1 FILLER_25_283 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X8 FILLER_26_65 ();
 FILLCELL_X4 FILLER_26_73 ();
 FILLCELL_X2 FILLER_26_77 ();
 FILLCELL_X1 FILLER_26_79 ();
 FILLCELL_X32 FILLER_26_90 ();
 FILLCELL_X4 FILLER_26_122 ();
 FILLCELL_X2 FILLER_26_126 ();
 FILLCELL_X32 FILLER_26_150 ();
 FILLCELL_X32 FILLER_26_182 ();
 FILLCELL_X32 FILLER_26_214 ();
 FILLCELL_X4 FILLER_26_249 ();
 FILLCELL_X1 FILLER_26_253 ();
 FILLCELL_X16 FILLER_26_257 ();
 FILLCELL_X8 FILLER_26_273 ();
 FILLCELL_X2 FILLER_26_281 ();
 FILLCELL_X1 FILLER_26_283 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X16 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_89 ();
 FILLCELL_X4 FILLER_27_121 ();
 FILLCELL_X4 FILLER_27_135 ();
 FILLCELL_X1 FILLER_27_139 ();
 FILLCELL_X1 FILLER_27_142 ();
 FILLCELL_X8 FILLER_27_145 ();
 FILLCELL_X4 FILLER_27_153 ();
 FILLCELL_X32 FILLER_27_167 ();
 FILLCELL_X4 FILLER_27_199 ();
 FILLCELL_X2 FILLER_27_203 ();
 FILLCELL_X1 FILLER_27_205 ();
 FILLCELL_X16 FILLER_27_220 ();
 FILLCELL_X8 FILLER_27_236 ();
 FILLCELL_X4 FILLER_27_244 ();
 FILLCELL_X32 FILLER_27_250 ();
 FILLCELL_X2 FILLER_27_282 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X8 FILLER_28_65 ();
 FILLCELL_X4 FILLER_28_73 ();
 FILLCELL_X4 FILLER_28_88 ();
 FILLCELL_X16 FILLER_28_109 ();
 FILLCELL_X1 FILLER_28_125 ();
 FILLCELL_X1 FILLER_28_142 ();
 FILLCELL_X1 FILLER_28_150 ();
 FILLCELL_X8 FILLER_28_155 ();
 FILLCELL_X2 FILLER_28_163 ();
 FILLCELL_X1 FILLER_28_165 ();
 FILLCELL_X2 FILLER_28_197 ();
 FILLCELL_X1 FILLER_28_199 ();
 FILLCELL_X32 FILLER_28_216 ();
 FILLCELL_X32 FILLER_28_248 ();
 FILLCELL_X4 FILLER_28_280 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X16 FILLER_29_33 ();
 FILLCELL_X8 FILLER_29_49 ();
 FILLCELL_X1 FILLER_29_57 ();
 FILLCELL_X1 FILLER_29_81 ();
 FILLCELL_X32 FILLER_29_89 ();
 FILLCELL_X8 FILLER_29_121 ();
 FILLCELL_X1 FILLER_29_129 ();
 FILLCELL_X8 FILLER_29_158 ();
 FILLCELL_X2 FILLER_29_166 ();
 FILLCELL_X16 FILLER_29_184 ();
 FILLCELL_X8 FILLER_29_200 ();
 FILLCELL_X4 FILLER_29_208 ();
 FILLCELL_X1 FILLER_29_212 ();
 FILLCELL_X32 FILLER_29_215 ();
 FILLCELL_X32 FILLER_29_247 ();
 FILLCELL_X4 FILLER_29_279 ();
 FILLCELL_X1 FILLER_29_283 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X8 FILLER_30_129 ();
 FILLCELL_X4 FILLER_30_137 ();
 FILLCELL_X1 FILLER_30_141 ();
 FILLCELL_X8 FILLER_30_152 ();
 FILLCELL_X2 FILLER_30_160 ();
 FILLCELL_X32 FILLER_30_172 ();
 FILLCELL_X1 FILLER_30_204 ();
 FILLCELL_X32 FILLER_30_211 ();
 FILLCELL_X32 FILLER_30_243 ();
 FILLCELL_X8 FILLER_30_275 ();
 FILLCELL_X1 FILLER_30_283 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X8 FILLER_31_129 ();
 FILLCELL_X2 FILLER_31_137 ();
 FILLCELL_X1 FILLER_31_139 ();
 FILLCELL_X8 FILLER_31_159 ();
 FILLCELL_X16 FILLER_31_171 ();
 FILLCELL_X4 FILLER_31_187 ();
 FILLCELL_X1 FILLER_31_191 ();
 FILLCELL_X1 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_228 ();
 FILLCELL_X16 FILLER_31_260 ();
 FILLCELL_X8 FILLER_31_276 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X16 FILLER_32_97 ();
 FILLCELL_X8 FILLER_32_113 ();
 FILLCELL_X2 FILLER_32_121 ();
 FILLCELL_X1 FILLER_32_123 ();
 FILLCELL_X32 FILLER_32_141 ();
 FILLCELL_X16 FILLER_32_173 ();
 FILLCELL_X4 FILLER_32_189 ();
 FILLCELL_X2 FILLER_32_193 ();
 FILLCELL_X4 FILLER_32_202 ();
 FILLCELL_X2 FILLER_32_206 ();
 FILLCELL_X1 FILLER_32_208 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X16 FILLER_32_257 ();
 FILLCELL_X8 FILLER_32_273 ();
 FILLCELL_X2 FILLER_32_281 ();
 FILLCELL_X1 FILLER_32_283 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X16 FILLER_33_161 ();
 FILLCELL_X8 FILLER_33_177 ();
 FILLCELL_X8 FILLER_33_189 ();
 FILLCELL_X32 FILLER_33_204 ();
 FILLCELL_X32 FILLER_33_236 ();
 FILLCELL_X16 FILLER_33_268 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X16 FILLER_34_129 ();
 FILLCELL_X1 FILLER_34_145 ();
 FILLCELL_X4 FILLER_34_149 ();
 FILLCELL_X2 FILLER_34_153 ();
 FILLCELL_X8 FILLER_34_169 ();
 FILLCELL_X4 FILLER_34_177 ();
 FILLCELL_X2 FILLER_34_181 ();
 FILLCELL_X32 FILLER_34_202 ();
 FILLCELL_X32 FILLER_34_234 ();
 FILLCELL_X16 FILLER_34_266 ();
 FILLCELL_X2 FILLER_34_282 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X8 FILLER_35_129 ();
 FILLCELL_X1 FILLER_35_137 ();
 FILLCELL_X2 FILLER_35_158 ();
 FILLCELL_X4 FILLER_35_174 ();
 FILLCELL_X1 FILLER_35_178 ();
 FILLCELL_X32 FILLER_35_202 ();
 FILLCELL_X32 FILLER_35_234 ();
 FILLCELL_X16 FILLER_35_266 ();
 FILLCELL_X2 FILLER_35_282 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X4 FILLER_36_129 ();
 FILLCELL_X4 FILLER_36_139 ();
 FILLCELL_X1 FILLER_36_143 ();
 FILLCELL_X2 FILLER_36_147 ();
 FILLCELL_X1 FILLER_36_149 ();
 FILLCELL_X32 FILLER_36_156 ();
 FILLCELL_X32 FILLER_36_188 ();
 FILLCELL_X32 FILLER_36_220 ();
 FILLCELL_X32 FILLER_36_252 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X4 FILLER_37_129 ();
 FILLCELL_X1 FILLER_37_133 ();
 FILLCELL_X2 FILLER_37_137 ();
 FILLCELL_X2 FILLER_37_148 ();
 FILLCELL_X1 FILLER_37_150 ();
 FILLCELL_X8 FILLER_37_154 ();
 FILLCELL_X2 FILLER_37_162 ();
 FILLCELL_X32 FILLER_37_167 ();
 FILLCELL_X32 FILLER_37_199 ();
 FILLCELL_X32 FILLER_37_231 ();
 FILLCELL_X16 FILLER_37_263 ();
 FILLCELL_X4 FILLER_37_279 ();
 FILLCELL_X1 FILLER_37_283 ();
endmodule
