module dual_clock_fifo (almost_empty,
    almost_full,
    empty,
    full,
    rd_clk,
    rd_en,
    rd_rst_n,
    wr_clk,
    wr_en,
    wr_rst_n,
    fifo_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 output empty;
 output full;
 input rd_clk;
 input rd_en;
 input rd_rst_n;
 input wr_clk;
 input wr_en;
 input wr_rst_n;
 output [4:0] fifo_count;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr_bin[0] ;
 wire \rd_ptr_bin[1] ;
 wire \rd_ptr_bin[2] ;
 wire \rd_ptr_bin[3] ;
 wire \rd_ptr_bin[4] ;
 wire \rd_ptr_bin_wr_sync[4] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray[3] ;
 wire \rd_ptr_gray_wr_sync1[0] ;
 wire \rd_ptr_gray_wr_sync1[1] ;
 wire \rd_ptr_gray_wr_sync1[2] ;
 wire \rd_ptr_gray_wr_sync1[3] ;
 wire \rd_ptr_gray_wr_sync1[4] ;
 wire \rd_ptr_gray_wr_sync2[0] ;
 wire \rd_ptr_gray_wr_sync2[1] ;
 wire \rd_ptr_gray_wr_sync2[2] ;
 wire \rd_ptr_gray_wr_sync2[3] ;
 wire \wr_ptr_bin[0] ;
 wire \wr_ptr_bin[1] ;
 wire \wr_ptr_bin[2] ;
 wire \wr_ptr_bin[3] ;
 wire \wr_ptr_bin[4] ;
 wire \wr_ptr_bin_rd_sync[4] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray[3] ;
 wire \wr_ptr_gray_rd_sync1[0] ;
 wire \wr_ptr_gray_rd_sync1[1] ;
 wire \wr_ptr_gray_rd_sync1[2] ;
 wire \wr_ptr_gray_rd_sync1[3] ;
 wire \wr_ptr_gray_rd_sync1[4] ;
 wire \wr_ptr_gray_rd_sync2[0] ;
 wire \wr_ptr_gray_rd_sync2[1] ;
 wire \wr_ptr_gray_rd_sync2[2] ;
 wire \wr_ptr_gray_rd_sync2[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;

 sky130_fd_sc_hd__xor2_4 _205_ (.A(\wr_ptr_bin[4] ),
    .B(\rd_ptr_bin_wr_sync[4] ),
    .X(_046_));
 sky130_fd_sc_hd__xor2_1 _206_ (.A(\wr_ptr_gray[1] ),
    .B(\rd_ptr_gray_wr_sync2[1] ),
    .X(_047_));
 sky130_fd_sc_hd__xor2_1 _207_ (.A(\wr_ptr_gray[0] ),
    .B(\rd_ptr_gray_wr_sync2[0] ),
    .X(_048_));
 sky130_fd_sc_hd__xor2_1 _208_ (.A(\wr_ptr_gray[2] ),
    .B(\rd_ptr_gray_wr_sync2[2] ),
    .X(_049_));
 sky130_fd_sc_hd__xor2_1 _209_ (.A(\wr_ptr_gray[3] ),
    .B(\rd_ptr_gray_wr_sync2[3] ),
    .X(_050_));
 sky130_fd_sc_hd__nor4_4 _210_ (.A(_047_),
    .B(_048_),
    .C(_049_),
    .D(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__and2_2 _211_ (.A(_046_),
    .B(_051_),
    .X(_052_));
 sky130_fd_sc_hd__buf_6 _212_ (.A(_052_),
    .X(net23));
 sky130_fd_sc_hd__xor2_4 _213_ (.A(\wr_ptr_bin_rd_sync[4] ),
    .B(\rd_ptr_bin[4] ),
    .X(_053_));
 sky130_fd_sc_hd__xnor2_1 _214_ (.A(\wr_ptr_gray_rd_sync2[1] ),
    .B(\rd_ptr_gray[1] ),
    .Y(_054_));
 sky130_fd_sc_hd__xnor2_1 _215_ (.A(\wr_ptr_gray_rd_sync2[0] ),
    .B(\rd_ptr_gray[0] ),
    .Y(_055_));
 sky130_fd_sc_hd__xnor2_1 _216_ (.A(\wr_ptr_gray_rd_sync2[2] ),
    .B(\rd_ptr_gray[2] ),
    .Y(_056_));
 sky130_fd_sc_hd__xnor2_1 _217_ (.A(\wr_ptr_gray_rd_sync2[3] ),
    .B(\rd_ptr_gray[3] ),
    .Y(_057_));
 sky130_fd_sc_hd__nand4_4 _218_ (.A(_054_),
    .B(_055_),
    .C(_056_),
    .D(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _219_ (.A(_053_),
    .B(_058_),
    .Y(net17));
 sky130_fd_sc_hd__o21ai_4 _220_ (.A1(_053_),
    .A2(_058_),
    .B1(net2),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _221_ (.A(_059_),
    .Y(_008_));
 sky130_fd_sc_hd__xor2_1 _222_ (.A(\wr_ptr_gray_rd_sync2[3] ),
    .B(\wr_ptr_bin_rd_sync[4] ),
    .X(_172_));
 sky130_fd_sc_hd__xnor2_1 _223_ (.A(\wr_ptr_gray_rd_sync2[2] ),
    .B(_172_),
    .Y(_060_));
 sky130_fd_sc_hd__xor2_2 _224_ (.A(\wr_ptr_gray_rd_sync2[1] ),
    .B(_060_),
    .X(_169_));
 sky130_fd_sc_hd__nand2_1 _225_ (.A(_178_),
    .B(_182_),
    .Y(_061_));
 sky130_fd_sc_hd__a21oi_1 _226_ (.A1(_178_),
    .A2(_181_),
    .B1(_177_),
    .Y(_062_));
 sky130_fd_sc_hd__o21ai_0 _227_ (.A1(_168_),
    .A2(_061_),
    .B1(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__xor2_1 _228_ (.A(_174_),
    .B(_063_),
    .X(net21));
 sky130_fd_sc_hd__inv_1 _229_ (.A(_204_),
    .Y(net18));
 sky130_fd_sc_hd__nand2b_1 _230_ (.A_N(_170_),
    .B(_178_),
    .Y(_064_));
 sky130_fd_sc_hd__nor2_1 _231_ (.A(_173_),
    .B(_177_),
    .Y(_065_));
 sky130_fd_sc_hd__nor2_1 _232_ (.A(_174_),
    .B(_173_),
    .Y(_066_));
 sky130_fd_sc_hd__a21oi_1 _233_ (.A1(_064_),
    .A2(_065_),
    .B1(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__xnor2_1 _234_ (.A(_053_),
    .B(_067_),
    .Y(net22));
 sky130_fd_sc_hd__xnor2_2 _235_ (.A(\rd_ptr_bin_wr_sync[4] ),
    .B(\rd_ptr_gray_wr_sync2[3] ),
    .Y(_183_));
 sky130_fd_sc_hd__xor2_2 _236_ (.A(\rd_ptr_gray_wr_sync2[2] ),
    .B(_183_),
    .X(_186_));
 sky130_fd_sc_hd__xor2_2 _237_ (.A(\rd_ptr_gray_wr_sync2[1] ),
    .B(_186_),
    .X(_165_));
 sky130_fd_sc_hd__buf_6 _238_ (.A(\rd_ptr_bin[0] ),
    .X(_068_));
 sky130_fd_sc_hd__buf_8 _239_ (.A(_068_),
    .X(_069_));
 sky130_fd_sc_hd__clkbuf_4 _240_ (.A(\rd_ptr_bin[1] ),
    .X(_070_));
 sky130_fd_sc_hd__buf_4 _241_ (.A(_070_),
    .X(_071_));
 sky130_fd_sc_hd__mux4_2 _242_ (.A0(\mem[8][0] ),
    .A1(\mem[9][0] ),
    .A2(\mem[10][0] ),
    .A3(\mem[11][0] ),
    .S0(_069_),
    .S1(_071_),
    .X(_072_));
 sky130_fd_sc_hd__buf_8 _243_ (.A(_068_),
    .X(_073_));
 sky130_fd_sc_hd__buf_4 _244_ (.A(_070_),
    .X(_074_));
 sky130_fd_sc_hd__mux4_1 _245_ (.A0(\mem[0][0] ),
    .A1(\mem[1][0] ),
    .A2(\mem[2][0] ),
    .A3(\mem[3][0] ),
    .S0(_073_),
    .S1(_074_),
    .X(_075_));
 sky130_fd_sc_hd__mux4_1 _246_ (.A0(\mem[12][0] ),
    .A1(\mem[13][0] ),
    .A2(\mem[14][0] ),
    .A3(\mem[15][0] ),
    .S0(_073_),
    .S1(_074_),
    .X(_076_));
 sky130_fd_sc_hd__buf_6 _247_ (.A(_068_),
    .X(_077_));
 sky130_fd_sc_hd__clkbuf_4 _248_ (.A(_070_),
    .X(_078_));
 sky130_fd_sc_hd__mux4_1 _249_ (.A0(\mem[4][0] ),
    .A1(\mem[5][0] ),
    .A2(\mem[6][0] ),
    .A3(\mem[7][0] ),
    .S0(_077_),
    .S1(_078_),
    .X(_079_));
 sky130_fd_sc_hd__buf_2 _250_ (.A(\rd_ptr_bin[3] ),
    .X(_080_));
 sky130_fd_sc_hd__inv_6 _251_ (.A(_080_),
    .Y(_171_));
 sky130_fd_sc_hd__buf_4 _252_ (.A(\rd_ptr_bin[2] ),
    .X(_081_));
 sky130_fd_sc_hd__mux4_1 _253_ (.A0(_072_),
    .A1(_075_),
    .A2(_076_),
    .A3(_079_),
    .S0(_171_),
    .S1(_081_),
    .X(_000_));
 sky130_fd_sc_hd__mux4_1 _254_ (.A0(\mem[8][1] ),
    .A1(\mem[9][1] ),
    .A2(\mem[10][1] ),
    .A3(\mem[11][1] ),
    .S0(_069_),
    .S1(_071_),
    .X(_082_));
 sky130_fd_sc_hd__mux4_1 _255_ (.A0(\mem[0][1] ),
    .A1(\mem[1][1] ),
    .A2(\mem[2][1] ),
    .A3(\mem[3][1] ),
    .S0(_073_),
    .S1(_074_),
    .X(_083_));
 sky130_fd_sc_hd__mux4_1 _256_ (.A0(\mem[12][1] ),
    .A1(\mem[13][1] ),
    .A2(\mem[14][1] ),
    .A3(\mem[15][1] ),
    .S0(_073_),
    .S1(_074_),
    .X(_084_));
 sky130_fd_sc_hd__mux4_1 _257_ (.A0(\mem[4][1] ),
    .A1(\mem[5][1] ),
    .A2(\mem[6][1] ),
    .A3(\mem[7][1] ),
    .S0(_077_),
    .S1(_078_),
    .X(_085_));
 sky130_fd_sc_hd__mux4_1 _258_ (.A0(_082_),
    .A1(_083_),
    .A2(_084_),
    .A3(_085_),
    .S0(_171_),
    .S1(_081_),
    .X(_001_));
 sky130_fd_sc_hd__mux4_1 _259_ (.A0(\mem[8][2] ),
    .A1(\mem[9][2] ),
    .A2(\mem[10][2] ),
    .A3(\mem[11][2] ),
    .S0(_069_),
    .S1(_071_),
    .X(_086_));
 sky130_fd_sc_hd__mux4_1 _260_ (.A0(\mem[0][2] ),
    .A1(\mem[1][2] ),
    .A2(\mem[2][2] ),
    .A3(\mem[3][2] ),
    .S0(_068_),
    .S1(_070_),
    .X(_087_));
 sky130_fd_sc_hd__mux4_2 _261_ (.A0(\mem[12][2] ),
    .A1(\mem[13][2] ),
    .A2(\mem[14][2] ),
    .A3(\mem[15][2] ),
    .S0(_073_),
    .S1(_074_),
    .X(_088_));
 sky130_fd_sc_hd__mux4_1 _262_ (.A0(\mem[4][2] ),
    .A1(\mem[5][2] ),
    .A2(\mem[6][2] ),
    .A3(\mem[7][2] ),
    .S0(_077_),
    .S1(_078_),
    .X(_089_));
 sky130_fd_sc_hd__mux4_1 _263_ (.A0(_086_),
    .A1(_087_),
    .A2(_088_),
    .A3(_089_),
    .S0(_171_),
    .S1(_081_),
    .X(_002_));
 sky130_fd_sc_hd__mux4_1 _264_ (.A0(\mem[8][3] ),
    .A1(\mem[9][3] ),
    .A2(\mem[10][3] ),
    .A3(\mem[11][3] ),
    .S0(_069_),
    .S1(_071_),
    .X(_090_));
 sky130_fd_sc_hd__mux4_1 _265_ (.A0(\mem[0][3] ),
    .A1(\mem[1][3] ),
    .A2(\mem[2][3] ),
    .A3(\mem[3][3] ),
    .S0(_068_),
    .S1(_070_),
    .X(_091_));
 sky130_fd_sc_hd__mux4_2 _266_ (.A0(\mem[12][3] ),
    .A1(\mem[13][3] ),
    .A2(\mem[14][3] ),
    .A3(\mem[15][3] ),
    .S0(_073_),
    .S1(_074_),
    .X(_092_));
 sky130_fd_sc_hd__mux4_1 _267_ (.A0(\mem[4][3] ),
    .A1(\mem[5][3] ),
    .A2(\mem[6][3] ),
    .A3(\mem[7][3] ),
    .S0(_077_),
    .S1(_078_),
    .X(_093_));
 sky130_fd_sc_hd__mux4_1 _268_ (.A0(_090_),
    .A1(_091_),
    .A2(_092_),
    .A3(_093_),
    .S0(_171_),
    .S1(_081_),
    .X(_003_));
 sky130_fd_sc_hd__mux4_1 _269_ (.A0(\mem[8][4] ),
    .A1(\mem[9][4] ),
    .A2(\mem[10][4] ),
    .A3(\mem[11][4] ),
    .S0(_069_),
    .S1(_071_),
    .X(_094_));
 sky130_fd_sc_hd__mux4_1 _270_ (.A0(\mem[0][4] ),
    .A1(\mem[1][4] ),
    .A2(\mem[2][4] ),
    .A3(\mem[3][4] ),
    .S0(_068_),
    .S1(_070_),
    .X(_095_));
 sky130_fd_sc_hd__mux4_2 _271_ (.A0(\mem[12][4] ),
    .A1(\mem[13][4] ),
    .A2(\mem[14][4] ),
    .A3(\mem[15][4] ),
    .S0(_073_),
    .S1(_074_),
    .X(_096_));
 sky130_fd_sc_hd__mux4_1 _272_ (.A0(\mem[4][4] ),
    .A1(\mem[5][4] ),
    .A2(\mem[6][4] ),
    .A3(\mem[7][4] ),
    .S0(_077_),
    .S1(_078_),
    .X(_097_));
 sky130_fd_sc_hd__mux4_1 _273_ (.A0(_094_),
    .A1(_095_),
    .A2(_096_),
    .A3(_097_),
    .S0(_171_),
    .S1(_081_),
    .X(_004_));
 sky130_fd_sc_hd__mux4_1 _274_ (.A0(\mem[8][5] ),
    .A1(\mem[9][5] ),
    .A2(\mem[10][5] ),
    .A3(\mem[11][5] ),
    .S0(_069_),
    .S1(_071_),
    .X(_098_));
 sky130_fd_sc_hd__mux4_1 _275_ (.A0(\mem[0][5] ),
    .A1(\mem[1][5] ),
    .A2(\mem[2][5] ),
    .A3(\mem[3][5] ),
    .S0(_068_),
    .S1(_070_),
    .X(_099_));
 sky130_fd_sc_hd__mux4_2 _276_ (.A0(\mem[12][5] ),
    .A1(\mem[13][5] ),
    .A2(\mem[14][5] ),
    .A3(\mem[15][5] ),
    .S0(_073_),
    .S1(_074_),
    .X(_100_));
 sky130_fd_sc_hd__mux4_1 _277_ (.A0(\mem[4][5] ),
    .A1(\mem[5][5] ),
    .A2(\mem[6][5] ),
    .A3(\mem[7][5] ),
    .S0(_077_),
    .S1(_078_),
    .X(_101_));
 sky130_fd_sc_hd__mux4_1 _278_ (.A0(_098_),
    .A1(_099_),
    .A2(_100_),
    .A3(_101_),
    .S0(_171_),
    .S1(_081_),
    .X(_005_));
 sky130_fd_sc_hd__mux4_1 _279_ (.A0(\mem[8][6] ),
    .A1(\mem[9][6] ),
    .A2(\mem[10][6] ),
    .A3(\mem[11][6] ),
    .S0(_069_),
    .S1(_071_),
    .X(_102_));
 sky130_fd_sc_hd__mux4_1 _280_ (.A0(\mem[0][6] ),
    .A1(\mem[1][6] ),
    .A2(\mem[2][6] ),
    .A3(\mem[3][6] ),
    .S0(_068_),
    .S1(_070_),
    .X(_103_));
 sky130_fd_sc_hd__mux4_1 _281_ (.A0(\mem[12][6] ),
    .A1(\mem[13][6] ),
    .A2(\mem[14][6] ),
    .A3(\mem[15][6] ),
    .S0(_073_),
    .S1(_074_),
    .X(_104_));
 sky130_fd_sc_hd__mux4_1 _282_ (.A0(\mem[4][6] ),
    .A1(\mem[5][6] ),
    .A2(\mem[6][6] ),
    .A3(\mem[7][6] ),
    .S0(_069_),
    .S1(_071_),
    .X(_105_));
 sky130_fd_sc_hd__mux4_2 _283_ (.A0(_102_),
    .A1(_103_),
    .A2(_104_),
    .A3(_105_),
    .S0(_171_),
    .S1(_081_),
    .X(_006_));
 sky130_fd_sc_hd__mux4_1 _284_ (.A0(\mem[8][7] ),
    .A1(\mem[9][7] ),
    .A2(\mem[10][7] ),
    .A3(\mem[11][7] ),
    .S0(_069_),
    .S1(_071_),
    .X(_106_));
 sky130_fd_sc_hd__mux4_1 _285_ (.A0(\mem[0][7] ),
    .A1(\mem[1][7] ),
    .A2(\mem[2][7] ),
    .A3(\mem[3][7] ),
    .S0(_068_),
    .S1(_070_),
    .X(_107_));
 sky130_fd_sc_hd__mux4_1 _286_ (.A0(\mem[12][7] ),
    .A1(\mem[13][7] ),
    .A2(\mem[14][7] ),
    .A3(\mem[15][7] ),
    .S0(_073_),
    .S1(_074_),
    .X(_108_));
 sky130_fd_sc_hd__mux4_1 _287_ (.A0(\mem[4][7] ),
    .A1(\mem[5][7] ),
    .A2(\mem[6][7] ),
    .A3(\mem[7][7] ),
    .S0(_069_),
    .S1(_071_),
    .X(_109_));
 sky130_fd_sc_hd__mux4_1 _288_ (.A0(_106_),
    .A1(_107_),
    .A2(_108_),
    .A3(_109_),
    .S0(_171_),
    .S1(_081_),
    .X(_007_));
 sky130_fd_sc_hd__buf_4 _289_ (.A(\wr_ptr_bin[2] ),
    .X(_110_));
 sky130_fd_sc_hd__buf_4 _290_ (.A(\wr_ptr_bin[3] ),
    .X(_111_));
 sky130_fd_sc_hd__nand2b_4 _291_ (.A_N(_110_),
    .B(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__nand2_2 _292_ (.A(net13),
    .B(_196_),
    .Y(_113_));
 sky130_fd_sc_hd__nor3_4 _293_ (.A(net23),
    .B(_112_),
    .C(_113_),
    .Y(_023_));
 sky130_fd_sc_hd__nand2_2 _294_ (.A(net13),
    .B(_199_),
    .Y(_114_));
 sky130_fd_sc_hd__nor3_4 _295_ (.A(net23),
    .B(_112_),
    .C(_114_),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_2 _296_ (.A(net13),
    .B(_197_),
    .Y(_115_));
 sky130_fd_sc_hd__nor3_4 _297_ (.A(net23),
    .B(_112_),
    .C(_115_),
    .Y(_010_));
 sky130_fd_sc_hd__nand2_4 _298_ (.A(net13),
    .B(_201_),
    .Y(_116_));
 sky130_fd_sc_hd__nor3_4 _299_ (.A(net23),
    .B(_112_),
    .C(_116_),
    .Y(_011_));
 sky130_fd_sc_hd__a21boi_4 _300_ (.A1(_046_),
    .A2(_051_),
    .B1_N(net13),
    .Y(_117_));
 sky130_fd_sc_hd__and2_0 _301_ (.A(_111_),
    .B(\wr_ptr_bin[2] ),
    .X(_118_));
 sky130_fd_sc_hd__and3_4 _302_ (.A(_196_),
    .B(_117_),
    .C(_118_),
    .X(_012_));
 sky130_fd_sc_hd__and3_4 _303_ (.A(_199_),
    .B(_117_),
    .C(_118_),
    .X(_013_));
 sky130_fd_sc_hd__and3_4 _304_ (.A(_197_),
    .B(_117_),
    .C(_118_),
    .X(_014_));
 sky130_fd_sc_hd__nand3_1 _305_ (.A(net13),
    .B(_201_),
    .C(_118_),
    .Y(_119_));
 sky130_fd_sc_hd__a21oi_4 _306_ (.A1(_046_),
    .A2(_051_),
    .B1(_119_),
    .Y(_015_));
 sky130_fd_sc_hd__inv_1 _307_ (.A(\rd_ptr_bin[2] ),
    .Y(_175_));
 sky130_fd_sc_hd__nor4_4 _308_ (.A(_111_),
    .B(_110_),
    .C(net23),
    .D(_113_),
    .Y(_009_));
 sky130_fd_sc_hd__nor4_4 _309_ (.A(_111_),
    .B(_110_),
    .C(_052_),
    .D(_116_),
    .Y(_018_));
 sky130_fd_sc_hd__nand2b_4 _310_ (.A_N(_111_),
    .B(_110_),
    .Y(_120_));
 sky130_fd_sc_hd__nor3_4 _311_ (.A(net23),
    .B(_114_),
    .C(_120_),
    .Y(_020_));
 sky130_fd_sc_hd__nor3_4 _312_ (.A(net23),
    .B(_115_),
    .C(_120_),
    .Y(_021_));
 sky130_fd_sc_hd__nor3_4 _313_ (.A(net23),
    .B(_116_),
    .C(_120_),
    .Y(_022_));
 sky130_fd_sc_hd__nor4_4 _314_ (.A(_111_),
    .B(_110_),
    .C(_052_),
    .D(_115_),
    .Y(_017_));
 sky130_fd_sc_hd__nor3_4 _315_ (.A(net23),
    .B(_113_),
    .C(_120_),
    .Y(_019_));
 sky130_fd_sc_hd__nor4_4 _316_ (.A(_111_),
    .B(_110_),
    .C(_052_),
    .D(_114_),
    .Y(_016_));
 sky130_fd_sc_hd__inv_1 _317_ (.A(_078_),
    .Y(_179_));
 sky130_fd_sc_hd__inv_1 _318_ (.A(_192_),
    .Y(_164_));
 sky130_fd_sc_hd__inv_1 _319_ (.A(\wr_ptr_bin[0] ),
    .Y(_025_));
 sky130_fd_sc_hd__inv_1 _320_ (.A(_060_),
    .Y(_176_));
 sky130_fd_sc_hd__inv_1 _321_ (.A(_169_),
    .Y(_180_));
 sky130_fd_sc_hd__xnor2_1 _322_ (.A(\rd_ptr_gray_wr_sync2[0] ),
    .B(_165_),
    .Y(_191_));
 sky130_fd_sc_hd__inv_1 _323_ (.A(\wr_ptr_bin[1] ),
    .Y(_195_));
 sky130_fd_sc_hd__xor2_1 _324_ (.A(\wr_ptr_gray_rd_sync2[0] ),
    .B(_169_),
    .X(_203_));
 sky130_fd_sc_hd__xnor2_1 _325_ (.A(_077_),
    .B(_059_),
    .Y(_028_));
 sky130_fd_sc_hd__mux2_1 _326_ (.A0(_027_),
    .A1(_078_),
    .S(_059_),
    .X(_029_));
 sky130_fd_sc_hd__o211ai_1 _327_ (.A1(_053_),
    .A2(_058_),
    .B1(net2),
    .C1(_194_),
    .Y(_121_));
 sky130_fd_sc_hd__xnor2_1 _328_ (.A(_081_),
    .B(_121_),
    .Y(_030_));
 sky130_fd_sc_hd__nand2_1 _329_ (.A(_077_),
    .B(_078_),
    .Y(_122_));
 sky130_fd_sc_hd__nor2_1 _330_ (.A(_175_),
    .B(_122_),
    .Y(_123_));
 sky130_fd_sc_hd__o211ai_1 _331_ (.A1(_053_),
    .A2(_058_),
    .B1(_123_),
    .C1(net2),
    .Y(_124_));
 sky130_fd_sc_hd__xnor2_1 _332_ (.A(_080_),
    .B(_124_),
    .Y(_031_));
 sky130_fd_sc_hd__xnor2_1 _333_ (.A(_077_),
    .B(_027_),
    .Y(_125_));
 sky130_fd_sc_hd__mux2_1 _334_ (.A0(_125_),
    .A1(\rd_ptr_gray[0] ),
    .S(_059_),
    .X(_032_));
 sky130_fd_sc_hd__xnor2_1 _335_ (.A(_194_),
    .B(_027_),
    .Y(_126_));
 sky130_fd_sc_hd__xnor2_1 _336_ (.A(_081_),
    .B(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__mux2_1 _337_ (.A0(_127_),
    .A1(\rd_ptr_gray[1] ),
    .S(_059_),
    .X(_033_));
 sky130_fd_sc_hd__xor2_1 _338_ (.A(_080_),
    .B(_194_),
    .X(_128_));
 sky130_fd_sc_hd__nand2_1 _339_ (.A(\rd_ptr_bin[2] ),
    .B(_122_),
    .Y(_129_));
 sky130_fd_sc_hd__xnor2_1 _340_ (.A(_128_),
    .B(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__mux2_1 _341_ (.A0(_130_),
    .A1(\rd_ptr_gray[2] ),
    .S(_059_),
    .X(_034_));
 sky130_fd_sc_hd__a21boi_0 _342_ (.A1(\rd_ptr_bin[2] ),
    .A2(_194_),
    .B1_N(_080_),
    .Y(_131_));
 sky130_fd_sc_hd__nand3b_1 _343_ (.A_N(_194_),
    .B(_080_),
    .C(\rd_ptr_bin[2] ),
    .Y(_132_));
 sky130_fd_sc_hd__o211a_1 _344_ (.A1(\rd_ptr_bin[2] ),
    .A2(_080_),
    .B1(_077_),
    .C1(_078_),
    .X(_133_));
 sky130_fd_sc_hd__a22oi_1 _345_ (.A1(_122_),
    .A2(_131_),
    .B1(_132_),
    .B2(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__xnor2_1 _346_ (.A(\rd_ptr_bin[4] ),
    .B(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__mux2_1 _347_ (.A0(_135_),
    .A1(\rd_ptr_gray[3] ),
    .S(_059_),
    .X(_035_));
 sky130_fd_sc_hd__nor2_1 _348_ (.A(_175_),
    .B(_171_),
    .Y(_136_));
 sky130_fd_sc_hd__o2111ai_1 _349_ (.A1(_053_),
    .A2(_058_),
    .B1(_136_),
    .C1(_194_),
    .D1(net2),
    .Y(_137_));
 sky130_fd_sc_hd__xnor2_1 _350_ (.A(\rd_ptr_bin[4] ),
    .B(_137_),
    .Y(_036_));
 sky130_fd_sc_hd__xnor2_1 _351_ (.A(_025_),
    .B(_117_),
    .Y(_037_));
 sky130_fd_sc_hd__mux2_1 _352_ (.A0(\wr_ptr_bin[1] ),
    .A1(_026_),
    .S(_117_),
    .X(_038_));
 sky130_fd_sc_hd__a21oi_1 _353_ (.A1(_046_),
    .A2(_051_),
    .B1(_116_),
    .Y(_138_));
 sky130_fd_sc_hd__xor2_1 _354_ (.A(_110_),
    .B(_138_),
    .X(_039_));
 sky130_fd_sc_hd__nand4_1 _355_ (.A(net13),
    .B(_110_),
    .C(\wr_ptr_bin[1] ),
    .D(\wr_ptr_bin[0] ),
    .Y(_139_));
 sky130_fd_sc_hd__a21oi_1 _356_ (.A1(_046_),
    .A2(_051_),
    .B1(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__xor2_1 _357_ (.A(_111_),
    .B(_140_),
    .X(_040_));
 sky130_fd_sc_hd__xnor2_1 _358_ (.A(\wr_ptr_bin[0] ),
    .B(_026_),
    .Y(_141_));
 sky130_fd_sc_hd__mux2_1 _359_ (.A0(\wr_ptr_gray[0] ),
    .A1(_141_),
    .S(_117_),
    .X(_041_));
 sky130_fd_sc_hd__xnor2_1 _360_ (.A(_201_),
    .B(_026_),
    .Y(_142_));
 sky130_fd_sc_hd__xnor2_1 _361_ (.A(_110_),
    .B(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__mux2_1 _362_ (.A0(\wr_ptr_gray[1] ),
    .A1(_143_),
    .S(_117_),
    .X(_042_));
 sky130_fd_sc_hd__xor2_1 _363_ (.A(_111_),
    .B(_201_),
    .X(_144_));
 sky130_fd_sc_hd__nand2_1 _364_ (.A(\wr_ptr_bin[1] ),
    .B(\wr_ptr_bin[0] ),
    .Y(_145_));
 sky130_fd_sc_hd__nand2_1 _365_ (.A(_110_),
    .B(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__xnor2_1 _366_ (.A(_144_),
    .B(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__mux2_1 _367_ (.A0(\wr_ptr_gray[2] ),
    .A1(_147_),
    .S(_117_),
    .X(_043_));
 sky130_fd_sc_hd__a21boi_0 _368_ (.A1(\wr_ptr_bin[2] ),
    .A2(_201_),
    .B1_N(\wr_ptr_bin[3] ),
    .Y(_148_));
 sky130_fd_sc_hd__nand3b_1 _369_ (.A_N(_201_),
    .B(\wr_ptr_bin[2] ),
    .C(_111_),
    .Y(_149_));
 sky130_fd_sc_hd__o211a_1 _370_ (.A1(\wr_ptr_bin[3] ),
    .A2(\wr_ptr_bin[2] ),
    .B1(\wr_ptr_bin[1] ),
    .C1(\wr_ptr_bin[0] ),
    .X(_150_));
 sky130_fd_sc_hd__a22oi_1 _371_ (.A1(_145_),
    .A2(_148_),
    .B1(_149_),
    .B2(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__xnor2_1 _372_ (.A(\wr_ptr_bin[4] ),
    .B(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__mux2_1 _373_ (.A0(\wr_ptr_gray[3] ),
    .A1(_152_),
    .S(_117_),
    .X(_044_));
 sky130_fd_sc_hd__xor2_1 _374_ (.A(\wr_ptr_bin[4] ),
    .B(_015_),
    .X(_045_));
 sky130_fd_sc_hd__xnor2_1 _375_ (.A(_170_),
    .B(_178_),
    .Y(net20));
 sky130_fd_sc_hd__o21a_1 _376_ (.A1(net19),
    .A2(net18),
    .B1(net20),
    .X(_153_));
 sky130_fd_sc_hd__o32ai_1 _377_ (.A1(net21),
    .A2(net22),
    .A3(_153_),
    .B1(_058_),
    .B2(_053_),
    .Y(net15));
 sky130_fd_sc_hd__inv_1 _378_ (.A(_187_),
    .Y(_154_));
 sky130_fd_sc_hd__nor2b_1 _379_ (.A(_192_),
    .B_N(_190_),
    .Y(_155_));
 sky130_fd_sc_hd__o21ai_0 _380_ (.A1(_189_),
    .A2(_155_),
    .B1(_188_),
    .Y(_156_));
 sky130_fd_sc_hd__a21boi_0 _381_ (.A1(_154_),
    .A2(_156_),
    .B1_N(_185_),
    .Y(_157_));
 sky130_fd_sc_hd__nor3b_1 _382_ (.A(_185_),
    .B(_187_),
    .C_N(_156_),
    .Y(_158_));
 sky130_fd_sc_hd__a21o_1 _383_ (.A1(_188_),
    .A2(_166_),
    .B1(_187_),
    .X(_159_));
 sky130_fd_sc_hd__a21oi_1 _384_ (.A1(_185_),
    .A2(_159_),
    .B1(_184_),
    .Y(_160_));
 sky130_fd_sc_hd__xnor2_1 _385_ (.A(_046_),
    .B(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__xor2_1 _386_ (.A(_188_),
    .B(_166_),
    .X(_162_));
 sky130_fd_sc_hd__a21oi_1 _387_ (.A1(_046_),
    .A2(_051_),
    .B1(_162_),
    .Y(_163_));
 sky130_fd_sc_hd__o211ai_1 _388_ (.A1(_157_),
    .A2(_158_),
    .B1(_161_),
    .C1(_163_),
    .Y(net16));
 sky130_fd_sc_hd__fa_1 _389_ (.A(\wr_ptr_bin[1] ),
    .B(_164_),
    .CIN(_165_),
    .COUT(_166_),
    .SUM(_167_));
 sky130_fd_sc_hd__fa_1 _390_ (.A(\rd_ptr_bin[1] ),
    .B(_168_),
    .CIN(_169_),
    .COUT(_170_),
    .SUM(net19));
 sky130_fd_sc_hd__ha_1 _391_ (.A(_171_),
    .B(_172_),
    .COUT(_173_),
    .SUM(_174_));
 sky130_fd_sc_hd__ha_1 _392_ (.A(_175_),
    .B(_176_),
    .COUT(_177_),
    .SUM(_178_));
 sky130_fd_sc_hd__ha_1 _393_ (.A(_179_),
    .B(_180_),
    .COUT(_181_),
    .SUM(_182_));
 sky130_fd_sc_hd__ha_1 _394_ (.A(\wr_ptr_bin[3] ),
    .B(_183_),
    .COUT(_184_),
    .SUM(_185_));
 sky130_fd_sc_hd__ha_1 _395_ (.A(\wr_ptr_bin[2] ),
    .B(_186_),
    .COUT(_187_),
    .SUM(_188_));
 sky130_fd_sc_hd__ha_1 _396_ (.A(\wr_ptr_bin[1] ),
    .B(_165_),
    .COUT(_189_),
    .SUM(_190_));
 sky130_fd_sc_hd__ha_1 _397_ (.A(_025_),
    .B(_191_),
    .COUT(_192_),
    .SUM(_193_));
 sky130_fd_sc_hd__ha_2 _398_ (.A(\rd_ptr_bin[0] ),
    .B(\rd_ptr_bin[1] ),
    .COUT(_194_),
    .SUM(_027_));
 sky130_fd_sc_hd__ha_1 _399_ (.A(_025_),
    .B(_195_),
    .COUT(_196_),
    .SUM(_026_));
 sky130_fd_sc_hd__ha_1 _400_ (.A(_025_),
    .B(\wr_ptr_bin[1] ),
    .COUT(_197_),
    .SUM(_198_));
 sky130_fd_sc_hd__ha_1 _401_ (.A(\wr_ptr_bin[0] ),
    .B(_195_),
    .COUT(_199_),
    .SUM(_200_));
 sky130_fd_sc_hd__ha_2 _402_ (.A(\wr_ptr_bin[0] ),
    .B(\wr_ptr_bin[1] ),
    .COUT(_201_),
    .SUM(_202_));
 sky130_fd_sc_hd__ha_1 _403_ (.A(\rd_ptr_bin[0] ),
    .B(_203_),
    .COUT(_168_),
    .SUM(_204_));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net5),
    .DE(_009_),
    .Q(\mem[0][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net6),
    .DE(_009_),
    .Q(\mem[0][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net7),
    .DE(_009_),
    .Q(\mem[0][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net8),
    .DE(_009_),
    .Q(\mem[0][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net9),
    .DE(_009_),
    .Q(\mem[0][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net10),
    .DE(_009_),
    .Q(\mem[0][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net11),
    .DE(_009_),
    .Q(\mem[0][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net12),
    .DE(_009_),
    .Q(\mem[0][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net5),
    .DE(_010_),
    .Q(\mem[10][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net6),
    .DE(_010_),
    .Q(\mem[10][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net7),
    .DE(_010_),
    .Q(\mem[10][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net8),
    .DE(_010_),
    .Q(\mem[10][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net9),
    .DE(_010_),
    .Q(\mem[10][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net10),
    .DE(_010_),
    .Q(\mem[10][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net11),
    .DE(_010_),
    .Q(\mem[10][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net12),
    .DE(_010_),
    .Q(\mem[10][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\mem[11][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\mem[11][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\mem[11][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\mem[11][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\mem[11][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net10),
    .DE(_011_),
    .Q(\mem[11][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net11),
    .DE(_011_),
    .Q(\mem[11][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net12),
    .DE(_011_),
    .Q(\mem[11][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\mem[12][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\mem[12][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\mem[12][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\mem[12][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\mem[12][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net10),
    .DE(_012_),
    .Q(\mem[12][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net11),
    .DE(_012_),
    .Q(\mem[12][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net12),
    .DE(_012_),
    .Q(\mem[12][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\mem[13][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\mem[13][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\mem[13][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\mem[13][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\mem[13][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net10),
    .DE(_013_),
    .Q(\mem[13][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net11),
    .DE(_013_),
    .Q(\mem[13][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net12),
    .DE(_013_),
    .Q(\mem[13][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\mem[14][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\mem[14][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\mem[14][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\mem[14][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\mem[14][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net10),
    .DE(_014_),
    .Q(\mem[14][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net11),
    .DE(_014_),
    .Q(\mem[14][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net12),
    .DE(_014_),
    .Q(\mem[14][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\mem[15][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\mem[15][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\mem[15][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\mem[15][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\mem[15][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net10),
    .DE(_015_),
    .Q(\mem[15][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net11),
    .DE(_015_),
    .Q(\mem[15][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net12),
    .DE(_015_),
    .Q(\mem[15][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net5),
    .DE(_016_),
    .Q(\mem[1][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net6),
    .DE(_016_),
    .Q(\mem[1][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net7),
    .DE(_016_),
    .Q(\mem[1][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net8),
    .DE(_016_),
    .Q(\mem[1][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net9),
    .DE(_016_),
    .Q(\mem[1][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net10),
    .DE(_016_),
    .Q(\mem[1][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net11),
    .DE(_016_),
    .Q(\mem[1][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net12),
    .DE(_016_),
    .Q(\mem[1][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net5),
    .DE(_017_),
    .Q(\mem[2][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net6),
    .DE(_017_),
    .Q(\mem[2][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net7),
    .DE(_017_),
    .Q(\mem[2][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net8),
    .DE(_017_),
    .Q(\mem[2][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net9),
    .DE(_017_),
    .Q(\mem[2][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net10),
    .DE(_017_),
    .Q(\mem[2][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net11),
    .DE(_017_),
    .Q(\mem[2][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net12),
    .DE(_017_),
    .Q(\mem[2][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net5),
    .DE(_018_),
    .Q(\mem[3][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net6),
    .DE(_018_),
    .Q(\mem[3][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net7),
    .DE(_018_),
    .Q(\mem[3][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net8),
    .DE(_018_),
    .Q(\mem[3][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net9),
    .DE(_018_),
    .Q(\mem[3][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net10),
    .DE(_018_),
    .Q(\mem[3][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net11),
    .DE(_018_),
    .Q(\mem[3][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net12),
    .DE(_018_),
    .Q(\mem[3][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net5),
    .DE(_019_),
    .Q(\mem[4][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net6),
    .DE(_019_),
    .Q(\mem[4][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net7),
    .DE(_019_),
    .Q(\mem[4][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net8),
    .DE(_019_),
    .Q(\mem[4][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net9),
    .DE(_019_),
    .Q(\mem[4][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net10),
    .DE(_019_),
    .Q(\mem[4][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net11),
    .DE(_019_),
    .Q(\mem[4][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net12),
    .DE(_019_),
    .Q(\mem[4][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net5),
    .DE(_020_),
    .Q(\mem[5][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net6),
    .DE(_020_),
    .Q(\mem[5][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net7),
    .DE(_020_),
    .Q(\mem[5][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net8),
    .DE(_020_),
    .Q(\mem[5][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net9),
    .DE(_020_),
    .Q(\mem[5][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net10),
    .DE(_020_),
    .Q(\mem[5][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net11),
    .DE(_020_),
    .Q(\mem[5][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net12),
    .DE(_020_),
    .Q(\mem[5][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net5),
    .DE(_021_),
    .Q(\mem[6][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net6),
    .DE(_021_),
    .Q(\mem[6][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net7),
    .DE(_021_),
    .Q(\mem[6][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net8),
    .DE(_021_),
    .Q(\mem[6][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net9),
    .DE(_021_),
    .Q(\mem[6][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net10),
    .DE(_021_),
    .Q(\mem[6][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net11),
    .DE(_021_),
    .Q(\mem[6][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net12),
    .DE(_021_),
    .Q(\mem[6][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net5),
    .DE(_022_),
    .Q(\mem[7][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net6),
    .DE(_022_),
    .Q(\mem[7][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net7),
    .DE(_022_),
    .Q(\mem[7][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net8),
    .DE(_022_),
    .Q(\mem[7][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net9),
    .DE(_022_),
    .Q(\mem[7][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net10),
    .DE(_022_),
    .Q(\mem[7][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net11),
    .DE(_022_),
    .Q(\mem[7][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net12),
    .DE(_022_),
    .Q(\mem[7][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net5),
    .DE(_023_),
    .Q(\mem[8][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net6),
    .DE(_023_),
    .Q(\mem[8][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net7),
    .DE(_023_),
    .Q(\mem[8][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net8),
    .DE(_023_),
    .Q(\mem[8][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net9),
    .DE(_023_),
    .Q(\mem[8][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net10),
    .DE(_023_),
    .Q(\mem[8][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net11),
    .DE(_023_),
    .Q(\mem[8][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net12),
    .DE(_023_),
    .Q(\mem[8][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net5),
    .DE(_024_),
    .Q(\mem[9][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net6),
    .DE(_024_),
    .Q(\mem[9][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net7),
    .DE(_024_),
    .Q(\mem[9][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net8),
    .DE(_024_),
    .Q(\mem[9][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net9),
    .DE(_024_),
    .Q(\mem[9][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net10),
    .DE(_024_),
    .Q(\mem[9][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net11),
    .DE(_024_),
    .Q(\mem[9][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net12),
    .DE(_024_),
    .Q(\mem[9][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[0]$_DFFE_PP_  (.D(_000_),
    .DE(_008_),
    .Q(net24),
    .CLK(net1));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[1]$_DFFE_PP_  (.D(_001_),
    .DE(_008_),
    .Q(net25),
    .CLK(net1));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[2]$_DFFE_PP_  (.D(_002_),
    .DE(_008_),
    .Q(net26),
    .CLK(net1));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[3]$_DFFE_PP_  (.D(_003_),
    .DE(_008_),
    .Q(net27),
    .CLK(net1));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[4]$_DFFE_PP_  (.D(_004_),
    .DE(_008_),
    .Q(net28),
    .CLK(net1));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[5]$_DFFE_PP_  (.D(_005_),
    .DE(_008_),
    .Q(net29),
    .CLK(net1));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[6]$_DFFE_PP_  (.D(_006_),
    .DE(_008_),
    .Q(net30),
    .CLK(net1));
 sky130_fd_sc_hd__edfxtp_1 \rd_data_reg[7]$_DFFE_PP_  (.D(_007_),
    .DE(_008_),
    .Q(net31),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[0]$_DFFE_PN0P_  (.D(_028_),
    .Q(\rd_ptr_bin[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[1]$_DFFE_PN0P_  (.D(_029_),
    .Q(\rd_ptr_bin[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[2]$_DFFE_PN0P_  (.D(_030_),
    .Q(\rd_ptr_bin[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[3]$_DFFE_PN0P_  (.D(_031_),
    .Q(\rd_ptr_bin[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[0]$_DFFE_PN0P_  (.D(_032_),
    .Q(\rd_ptr_gray[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[1]$_DFFE_PN0P_  (.D(_033_),
    .Q(\rd_ptr_gray[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[2]$_DFFE_PN0P_  (.D(_034_),
    .Q(\rd_ptr_gray[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[3]$_DFFE_PN0P_  (.D(_035_),
    .Q(\rd_ptr_gray[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_4 \rd_ptr_gray[4]$_DFFE_PN0P_  (.D(_036_),
    .Q(\rd_ptr_bin[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_wr_sync1[0]$_DFF_PN0_  (.D(\rd_ptr_gray[0] ),
    .Q(\rd_ptr_gray_wr_sync1[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_wr_sync1[1]$_DFF_PN0_  (.D(\rd_ptr_gray[1] ),
    .Q(\rd_ptr_gray_wr_sync1[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_wr_sync1[2]$_DFF_PN0_  (.D(\rd_ptr_gray[2] ),
    .Q(\rd_ptr_gray_wr_sync1[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_wr_sync1[3]$_DFF_PN0_  (.D(\rd_ptr_gray[3] ),
    .Q(\rd_ptr_gray_wr_sync1[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_wr_sync1[4]$_DFF_PN0_  (.D(\rd_ptr_bin[4] ),
    .Q(\rd_ptr_gray_wr_sync1[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_wr_sync2[0]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[0] ),
    .Q(\rd_ptr_gray_wr_sync2[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr_gray_wr_sync2[1]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[1] ),
    .Q(\rd_ptr_gray_wr_sync2[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_wr_sync2[2]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[2] ),
    .Q(\rd_ptr_gray_wr_sync2[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_wr_sync2[3]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[3] ),
    .Q(\rd_ptr_gray_wr_sync2[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr_gray_wr_sync2[4]$_DFF_PN0_  (.D(\rd_ptr_gray_wr_sync1[4] ),
    .Q(\rd_ptr_bin_wr_sync[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr_bin[0]$_DFFE_PN0P_  (.D(_037_),
    .Q(\wr_ptr_bin[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr_bin[1]$_DFFE_PN0P_  (.D(_038_),
    .Q(\wr_ptr_bin[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_bin[2]$_DFFE_PN0P_  (.D(_039_),
    .Q(\wr_ptr_bin[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_bin[3]$_DFFE_PN0P_  (.D(_040_),
    .Q(\wr_ptr_bin[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[0]$_DFFE_PN0P_  (.D(_041_),
    .Q(\wr_ptr_gray[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[1]$_DFFE_PN0P_  (.D(_042_),
    .Q(\wr_ptr_gray[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[2]$_DFFE_PN0P_  (.D(_043_),
    .Q(\wr_ptr_gray[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[3]$_DFFE_PN0P_  (.D(_044_),
    .Q(\wr_ptr_gray[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr_gray[4]$_DFFE_PN0P_  (.D(_045_),
    .Q(\wr_ptr_bin[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_rd_sync1[0]$_DFF_PN0_  (.D(\wr_ptr_gray[0] ),
    .Q(\wr_ptr_gray_rd_sync1[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_rd_sync1[1]$_DFF_PN0_  (.D(\wr_ptr_gray[1] ),
    .Q(\wr_ptr_gray_rd_sync1[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_rd_sync1[2]$_DFF_PN0_  (.D(\wr_ptr_gray[2] ),
    .Q(\wr_ptr_gray_rd_sync1[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_rd_sync1[3]$_DFF_PN0_  (.D(\wr_ptr_gray[3] ),
    .Q(\wr_ptr_gray_rd_sync1[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_rd_sync1[4]$_DFF_PN0_  (.D(\wr_ptr_bin[4] ),
    .Q(\wr_ptr_gray_rd_sync1[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_rd_sync2[0]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[0] ),
    .Q(\wr_ptr_gray_rd_sync2[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_rd_sync2[1]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[1] ),
    .Q(\wr_ptr_gray_rd_sync2[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_rd_sync2[2]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[2] ),
    .Q(\wr_ptr_gray_rd_sync2[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_rd_sync2[3]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[3] ),
    .Q(\wr_ptr_gray_rd_sync2[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr_gray_rd_sync2[4]$_DFF_PN0_  (.D(\wr_ptr_gray_rd_sync1[4] ),
    .Q(\wr_ptr_bin_rd_sync[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_171 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(rd_clk),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(rd_en),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(rd_rst_n),
    .X(net3));
 sky130_fd_sc_hd__buf_16 input4 (.A(wr_clk),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(wr_data[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(wr_data[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(wr_data[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(wr_data[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(wr_data[4]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input10 (.A(wr_data[5]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(wr_data[6]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(wr_data[7]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(wr_en),
    .X(net13));
 sky130_fd_sc_hd__buf_6 input14 (.A(wr_rst_n),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(fifo_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(fifo_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(fifo_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(fifo_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(fifo_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .X(rd_data[7]));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_241 ();
endmodule
