module parameterized_loadable_counter (clk,
    enable,
    load,
    rst_n,
    count,
    data_in);
 input clk;
 input enable;
 input load;
 input rst_n;
 output [7:0] count;
 input [7:0] data_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X2 _055_ (.A(rst_n),
    .Z(_009_));
 INV_X1 _056_ (.A(_009_),
    .ZN(_010_));
 BUF_X2 _057_ (.A(load),
    .Z(_011_));
 INV_X1 _058_ (.A(_011_),
    .ZN(_012_));
 CLKBUF_X3 _059_ (.A(_012_),
    .Z(_013_));
 NOR2_X1 _060_ (.A1(_013_),
    .A2(net1),
    .ZN(_014_));
 BUF_X4 _061_ (.A(enable),
    .Z(_015_));
 MUX2_X1 _062_ (.A(net9),
    .B(_000_),
    .S(_015_),
    .Z(_016_));
 NOR2_X1 _063_ (.A1(_011_),
    .A2(_016_),
    .ZN(_017_));
 NOR3_X1 _064_ (.A1(_010_),
    .A2(_014_),
    .A3(_017_),
    .ZN(_001_));
 NOR2_X1 _065_ (.A1(_013_),
    .A2(net2),
    .ZN(_018_));
 MUX2_X1 _066_ (.A(net10),
    .B(_054_),
    .S(_015_),
    .Z(_019_));
 NOR2_X1 _067_ (.A1(_011_),
    .A2(_019_),
    .ZN(_020_));
 NOR3_X1 _068_ (.A1(_010_),
    .A2(_018_),
    .A3(_020_),
    .ZN(_002_));
 NOR2_X1 _069_ (.A1(_013_),
    .A2(net3),
    .ZN(_021_));
 BUF_X4 _070_ (.A(net11),
    .Z(_022_));
 NAND2_X1 _071_ (.A1(_015_),
    .A2(_053_),
    .ZN(_023_));
 XNOR2_X1 _072_ (.A(_022_),
    .B(_023_),
    .ZN(_024_));
 NOR2_X1 _073_ (.A1(_011_),
    .A2(_024_),
    .ZN(_025_));
 NOR3_X1 _074_ (.A1(_010_),
    .A2(_021_),
    .A3(_025_),
    .ZN(_003_));
 OAI21_X1 _075_ (.A(_009_),
    .B1(net4),
    .B2(_013_),
    .ZN(_026_));
 NAND4_X1 _076_ (.A1(_015_),
    .A2(_022_),
    .A3(net10),
    .A4(net9),
    .ZN(_027_));
 XOR2_X1 _077_ (.A(net12),
    .B(_027_),
    .Z(_028_));
 AOI21_X1 _078_ (.A(_026_),
    .B1(_028_),
    .B2(_013_),
    .ZN(_004_));
 OAI21_X1 _079_ (.A(_009_),
    .B1(net5),
    .B2(_013_),
    .ZN(_029_));
 NAND4_X1 _080_ (.A1(_015_),
    .A2(_053_),
    .A3(_022_),
    .A4(net12),
    .ZN(_030_));
 XOR2_X1 _081_ (.A(net13),
    .B(_030_),
    .Z(_031_));
 AOI21_X1 _082_ (.A(_029_),
    .B1(_031_),
    .B2(_013_),
    .ZN(_005_));
 OAI21_X1 _083_ (.A(_009_),
    .B1(net6),
    .B2(_012_),
    .ZN(_032_));
 AND3_X1 _084_ (.A1(_022_),
    .A2(net12),
    .A3(net13),
    .ZN(_033_));
 NAND4_X1 _085_ (.A1(_015_),
    .A2(net10),
    .A3(net9),
    .A4(_033_),
    .ZN(_034_));
 XOR2_X1 _086_ (.A(net14),
    .B(_034_),
    .Z(_035_));
 AOI21_X1 _087_ (.A(_032_),
    .B1(_035_),
    .B2(_013_),
    .ZN(_006_));
 OAI21_X1 _088_ (.A(_009_),
    .B1(net7),
    .B2(_012_),
    .ZN(_036_));
 NAND4_X1 _089_ (.A1(_022_),
    .A2(net12),
    .A3(net13),
    .A4(net14),
    .ZN(_037_));
 NOR2_X1 _090_ (.A1(_023_),
    .A2(_037_),
    .ZN(_038_));
 XNOR2_X1 _091_ (.A(net15),
    .B(_038_),
    .ZN(_039_));
 AOI21_X1 _092_ (.A(_036_),
    .B1(_039_),
    .B2(_013_),
    .ZN(_007_));
 NOR2_X1 _093_ (.A1(_011_),
    .A2(_015_),
    .ZN(_040_));
 AOI22_X1 _094_ (.A1(_011_),
    .A2(net8),
    .B1(_040_),
    .B2(net16),
    .ZN(_041_));
 NAND3_X1 _095_ (.A1(_013_),
    .A2(_015_),
    .A3(_009_),
    .ZN(_042_));
 NAND3_X1 _096_ (.A1(net10),
    .A2(net9),
    .A3(net15),
    .ZN(_043_));
 NOR2_X1 _097_ (.A1(_037_),
    .A2(_043_),
    .ZN(_044_));
 XNOR2_X1 _098_ (.A(net16),
    .B(_044_),
    .ZN(_045_));
 OAI22_X1 _099_ (.A1(_010_),
    .A2(_041_),
    .B1(_042_),
    .B2(_045_),
    .ZN(_008_));
 HA_X1 _100_ (.A(net9),
    .B(net10),
    .CO(_053_),
    .S(_054_));
 DFF_X2 \counter_reg[0]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net9),
    .QN(_000_));
 DFF_X2 \counter_reg[1]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net10),
    .QN(_052_));
 DFF_X1 \counter_reg[2]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net11),
    .QN(_051_));
 DFF_X2 \counter_reg[3]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net12),
    .QN(_050_));
 DFF_X2 \counter_reg[4]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net13),
    .QN(_049_));
 DFF_X1 \counter_reg[5]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net14),
    .QN(_048_));
 DFF_X1 \counter_reg[6]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net15),
    .QN(_047_));
 DFF_X1 \counter_reg[7]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net16),
    .QN(_046_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_63 ();
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[2]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[3]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[5]),
    .Z(net6));
 BUF_X1 input7 (.A(data_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[7]),
    .Z(net8));
 BUF_X1 output9 (.A(net9),
    .Z(count[0]));
 BUF_X1 output10 (.A(net10),
    .Z(count[1]));
 BUF_X1 output11 (.A(net11),
    .Z(count[2]));
 BUF_X1 output12 (.A(net12),
    .Z(count[3]));
 BUF_X1 output13 (.A(net13),
    .Z(count[4]));
 BUF_X1 output14 (.A(net14),
    .Z(count[5]));
 BUF_X1 output15 (.A(net15),
    .Z(count[6]));
 BUF_X1 output16 (.A(net16),
    .Z(count[7]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X8 FILLER_0_97 ();
 FILLCELL_X4 FILLER_0_105 ();
 FILLCELL_X8 FILLER_0_115 ();
 FILLCELL_X32 FILLER_0_126 ();
 FILLCELL_X32 FILLER_0_158 ();
 FILLCELL_X32 FILLER_0_190 ();
 FILLCELL_X8 FILLER_0_222 ();
 FILLCELL_X4 FILLER_0_230 ();
 FILLCELL_X2 FILLER_0_234 ();
 FILLCELL_X1 FILLER_0_236 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X8 FILLER_1_97 ();
 FILLCELL_X2 FILLER_1_105 ();
 FILLCELL_X16 FILLER_1_110 ();
 FILLCELL_X2 FILLER_1_126 ();
 FILLCELL_X32 FILLER_1_131 ();
 FILLCELL_X32 FILLER_1_163 ();
 FILLCELL_X32 FILLER_1_195 ();
 FILLCELL_X8 FILLER_1_227 ();
 FILLCELL_X2 FILLER_1_235 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X8 FILLER_2_225 ();
 FILLCELL_X4 FILLER_2_233 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X8 FILLER_3_225 ();
 FILLCELL_X4 FILLER_3_233 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X8 FILLER_4_225 ();
 FILLCELL_X4 FILLER_4_233 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_102 ();
 FILLCELL_X32 FILLER_5_134 ();
 FILLCELL_X32 FILLER_5_166 ();
 FILLCELL_X32 FILLER_5_198 ();
 FILLCELL_X4 FILLER_5_230 ();
 FILLCELL_X2 FILLER_5_234 ();
 FILLCELL_X1 FILLER_5_236 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X8 FILLER_6_97 ();
 FILLCELL_X1 FILLER_6_105 ();
 FILLCELL_X32 FILLER_6_109 ();
 FILLCELL_X32 FILLER_6_141 ();
 FILLCELL_X32 FILLER_6_173 ();
 FILLCELL_X32 FILLER_6_205 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_65 ();
 FILLCELL_X8 FILLER_7_81 ();
 FILLCELL_X4 FILLER_7_89 ();
 FILLCELL_X4 FILLER_7_119 ();
 FILLCELL_X4 FILLER_7_145 ();
 FILLCELL_X1 FILLER_7_149 ();
 FILLCELL_X32 FILLER_7_157 ();
 FILLCELL_X32 FILLER_7_189 ();
 FILLCELL_X16 FILLER_7_221 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X4 FILLER_8_97 ();
 FILLCELL_X2 FILLER_8_101 ();
 FILLCELL_X1 FILLER_8_103 ();
 FILLCELL_X8 FILLER_8_111 ();
 FILLCELL_X4 FILLER_8_119 ();
 FILLCELL_X2 FILLER_8_127 ();
 FILLCELL_X1 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_133 ();
 FILLCELL_X32 FILLER_8_165 ();
 FILLCELL_X32 FILLER_8_197 ();
 FILLCELL_X8 FILLER_8_229 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X16 FILLER_9_97 ();
 FILLCELL_X2 FILLER_9_113 ();
 FILLCELL_X1 FILLER_9_115 ();
 FILLCELL_X32 FILLER_9_126 ();
 FILLCELL_X32 FILLER_9_158 ();
 FILLCELL_X32 FILLER_9_190 ();
 FILLCELL_X8 FILLER_9_222 ();
 FILLCELL_X4 FILLER_9_230 ();
 FILLCELL_X2 FILLER_9_234 ();
 FILLCELL_X1 FILLER_9_236 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X16 FILLER_10_97 ();
 FILLCELL_X1 FILLER_10_113 ();
 FILLCELL_X1 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_151 ();
 FILLCELL_X32 FILLER_10_183 ();
 FILLCELL_X16 FILLER_10_215 ();
 FILLCELL_X4 FILLER_10_231 ();
 FILLCELL_X2 FILLER_10_235 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X1 FILLER_11_97 ();
 FILLCELL_X2 FILLER_11_110 ();
 FILLCELL_X1 FILLER_11_112 ();
 FILLCELL_X8 FILLER_11_115 ();
 FILLCELL_X2 FILLER_11_123 ();
 FILLCELL_X1 FILLER_11_125 ();
 FILLCELL_X4 FILLER_11_129 ();
 FILLCELL_X1 FILLER_11_133 ();
 FILLCELL_X32 FILLER_11_141 ();
 FILLCELL_X16 FILLER_11_173 ();
 FILLCELL_X8 FILLER_11_189 ();
 FILLCELL_X4 FILLER_11_197 ();
 FILLCELL_X32 FILLER_11_204 ();
 FILLCELL_X1 FILLER_11_236 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_36 ();
 FILLCELL_X16 FILLER_12_68 ();
 FILLCELL_X4 FILLER_12_84 ();
 FILLCELL_X8 FILLER_12_110 ();
 FILLCELL_X4 FILLER_12_118 ();
 FILLCELL_X1 FILLER_12_122 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X8 FILLER_12_225 ();
 FILLCELL_X4 FILLER_12_233 ();
 FILLCELL_X32 FILLER_13_4 ();
 FILLCELL_X32 FILLER_13_36 ();
 FILLCELL_X32 FILLER_13_68 ();
 FILLCELL_X1 FILLER_13_100 ();
 FILLCELL_X16 FILLER_13_107 ();
 FILLCELL_X2 FILLER_13_123 ();
 FILLCELL_X1 FILLER_13_125 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X8 FILLER_13_225 ();
 FILLCELL_X4 FILLER_13_233 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X4 FILLER_14_97 ();
 FILLCELL_X2 FILLER_14_101 ();
 FILLCELL_X1 FILLER_14_103 ();
 FILLCELL_X16 FILLER_14_108 ();
 FILLCELL_X2 FILLER_14_124 ();
 FILLCELL_X1 FILLER_14_126 ();
 FILLCELL_X32 FILLER_14_147 ();
 FILLCELL_X32 FILLER_14_179 ();
 FILLCELL_X16 FILLER_14_211 ();
 FILLCELL_X8 FILLER_14_227 ();
 FILLCELL_X2 FILLER_14_235 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X4 FILLER_15_97 ();
 FILLCELL_X2 FILLER_15_101 ();
 FILLCELL_X1 FILLER_15_103 ();
 FILLCELL_X8 FILLER_15_107 ();
 FILLCELL_X2 FILLER_15_115 ();
 FILLCELL_X2 FILLER_15_125 ();
 FILLCELL_X32 FILLER_15_138 ();
 FILLCELL_X32 FILLER_15_170 ();
 FILLCELL_X32 FILLER_15_202 ();
 FILLCELL_X2 FILLER_15_234 ();
 FILLCELL_X1 FILLER_15_236 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X4 FILLER_16_97 ();
 FILLCELL_X1 FILLER_16_101 ();
 FILLCELL_X32 FILLER_16_104 ();
 FILLCELL_X32 FILLER_16_136 ();
 FILLCELL_X32 FILLER_16_168 ();
 FILLCELL_X32 FILLER_16_203 ();
 FILLCELL_X2 FILLER_16_235 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X16 FILLER_17_65 ();
 FILLCELL_X8 FILLER_17_81 ();
 FILLCELL_X2 FILLER_17_89 ();
 FILLCELL_X16 FILLER_17_97 ();
 FILLCELL_X8 FILLER_17_113 ();
 FILLCELL_X2 FILLER_17_121 ();
 FILLCELL_X32 FILLER_17_146 ();
 FILLCELL_X32 FILLER_17_178 ();
 FILLCELL_X16 FILLER_17_210 ();
 FILLCELL_X8 FILLER_17_226 ();
 FILLCELL_X2 FILLER_17_234 ();
 FILLCELL_X1 FILLER_17_236 ();
 FILLCELL_X16 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_17 ();
 FILLCELL_X1 FILLER_18_19 ();
 FILLCELL_X16 FILLER_18_23 ();
 FILLCELL_X8 FILLER_18_39 ();
 FILLCELL_X1 FILLER_18_47 ();
 FILLCELL_X32 FILLER_18_52 ();
 FILLCELL_X4 FILLER_18_84 ();
 FILLCELL_X2 FILLER_18_88 ();
 FILLCELL_X1 FILLER_18_90 ();
 FILLCELL_X8 FILLER_18_108 ();
 FILLCELL_X4 FILLER_18_116 ();
 FILLCELL_X2 FILLER_18_120 ();
 FILLCELL_X2 FILLER_18_126 ();
 FILLCELL_X1 FILLER_18_128 ();
 FILLCELL_X32 FILLER_18_141 ();
 FILLCELL_X32 FILLER_18_173 ();
 FILLCELL_X32 FILLER_18_205 ();
 FILLCELL_X16 FILLER_19_1 ();
 FILLCELL_X8 FILLER_19_17 ();
 FILLCELL_X1 FILLER_19_25 ();
 FILLCELL_X32 FILLER_19_29 ();
 FILLCELL_X16 FILLER_19_61 ();
 FILLCELL_X8 FILLER_19_77 ();
 FILLCELL_X4 FILLER_19_85 ();
 FILLCELL_X8 FILLER_19_106 ();
 FILLCELL_X1 FILLER_19_114 ();
 FILLCELL_X4 FILLER_19_119 ();
 FILLCELL_X32 FILLER_19_136 ();
 FILLCELL_X32 FILLER_19_168 ();
 FILLCELL_X32 FILLER_19_200 ();
 FILLCELL_X4 FILLER_19_232 ();
 FILLCELL_X1 FILLER_19_236 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X16 FILLER_20_97 ();
 FILLCELL_X8 FILLER_20_113 ();
 FILLCELL_X4 FILLER_20_121 ();
 FILLCELL_X2 FILLER_20_125 ();
 FILLCELL_X1 FILLER_20_127 ();
 FILLCELL_X32 FILLER_20_147 ();
 FILLCELL_X32 FILLER_20_179 ();
 FILLCELL_X16 FILLER_20_211 ();
 FILLCELL_X8 FILLER_20_227 ();
 FILLCELL_X2 FILLER_20_235 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X16 FILLER_21_97 ();
 FILLCELL_X1 FILLER_21_113 ();
 FILLCELL_X32 FILLER_21_131 ();
 FILLCELL_X32 FILLER_21_163 ();
 FILLCELL_X32 FILLER_21_195 ();
 FILLCELL_X8 FILLER_21_227 ();
 FILLCELL_X2 FILLER_21_235 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X8 FILLER_22_225 ();
 FILLCELL_X4 FILLER_22_233 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X8 FILLER_23_225 ();
 FILLCELL_X4 FILLER_23_233 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X8 FILLER_24_225 ();
 FILLCELL_X4 FILLER_24_233 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X8 FILLER_25_225 ();
 FILLCELL_X4 FILLER_25_233 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X8 FILLER_26_225 ();
 FILLCELL_X4 FILLER_26_233 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X8 FILLER_27_225 ();
 FILLCELL_X4 FILLER_27_233 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X8 FILLER_28_225 ();
 FILLCELL_X4 FILLER_28_233 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X8 FILLER_29_225 ();
 FILLCELL_X4 FILLER_29_233 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X4 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_136 ();
 FILLCELL_X32 FILLER_30_168 ();
 FILLCELL_X32 FILLER_30_200 ();
 FILLCELL_X4 FILLER_30_232 ();
 FILLCELL_X1 FILLER_30_236 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X4 FILLER_31_97 ();
 FILLCELL_X2 FILLER_31_101 ();
 FILLCELL_X8 FILLER_31_106 ();
 FILLCELL_X4 FILLER_31_114 ();
 FILLCELL_X2 FILLER_31_118 ();
 FILLCELL_X1 FILLER_31_120 ();
 FILLCELL_X16 FILLER_31_127 ();
 FILLCELL_X4 FILLER_31_143 ();
 FILLCELL_X32 FILLER_31_150 ();
 FILLCELL_X32 FILLER_31_182 ();
 FILLCELL_X16 FILLER_31_214 ();
 FILLCELL_X4 FILLER_31_230 ();
 FILLCELL_X2 FILLER_31_234 ();
 FILLCELL_X1 FILLER_31_236 ();
endmodule
