module pwm_generator (clk,
    enable,
    pwm_out,
    rst_n,
    duty_cycle,
    period);
 input clk;
 input enable;
 output pwm_out;
 input rst_n;
 input [7:0] duty_cycle;
 input [7:0] period;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \duty_reg[0] ;
 wire \duty_reg[1] ;
 wire \duty_reg[2] ;
 wire \duty_reg[3] ;
 wire \duty_reg[4] ;
 wire \duty_reg[5] ;
 wire \duty_reg[6] ;
 wire \duty_reg[7] ;
 wire \period_reg[0] ;
 wire \period_reg[1] ;
 wire \period_reg[2] ;
 wire \period_reg[3] ;
 wire \period_reg[4] ;
 wire \period_reg[5] ;
 wire \period_reg[6] ;
 wire \period_reg[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X1 _188_ (.A(rst_n),
    .Z(_025_));
 INV_X1 _189_ (.A(_025_),
    .ZN(_026_));
 CLKBUF_X3 _190_ (.A(_026_),
    .Z(_027_));
 BUF_X4 _191_ (.A(enable),
    .Z(_028_));
 INV_X2 _192_ (.A(_028_),
    .ZN(_029_));
 AOI21_X1 _193_ (.A(_154_),
    .B1(_157_),
    .B2(_155_),
    .ZN(_030_));
 AOI21_X1 _194_ (.A(_160_),
    .B1(_163_),
    .B2(_161_),
    .ZN(_031_));
 NAND2_X1 _195_ (.A1(_155_),
    .A2(_158_),
    .ZN(_032_));
 OAI21_X1 _196_ (.A(_030_),
    .B1(_031_),
    .B2(_032_),
    .ZN(_033_));
 NOR3_X1 _197_ (.A1(\counter[0] ),
    .A2(_029_),
    .A3(_033_),
    .ZN(_034_));
 INV_X1 _198_ (.A(_148_),
    .ZN(_035_));
 NAND4_X4 _199_ (.A1(_146_),
    .A2(_149_),
    .A3(_143_),
    .A4(_152_),
    .ZN(_036_));
 NAND2_X1 _200_ (.A1(_035_),
    .A2(_036_),
    .ZN(_037_));
 OAI21_X1 _201_ (.A(_149_),
    .B1(_152_),
    .B2(_151_),
    .ZN(_038_));
 INV_X1 _202_ (.A(_038_),
    .ZN(_039_));
 NOR2_X1 _203_ (.A1(_145_),
    .A2(_151_),
    .ZN(_040_));
 INV_X1 _204_ (.A(_146_),
    .ZN(_041_));
 OAI21_X2 _205_ (.A(_040_),
    .B1(_142_),
    .B2(_041_),
    .ZN(_042_));
 AOI21_X4 _206_ (.A(_037_),
    .B1(_039_),
    .B2(_042_),
    .ZN(_043_));
 NAND4_X4 _207_ (.A1(_155_),
    .A2(_164_),
    .A3(_161_),
    .A4(_158_),
    .ZN(_044_));
 OAI21_X1 _208_ (.A(_034_),
    .B1(_043_),
    .B2(_044_),
    .ZN(_045_));
 NAND2_X1 _209_ (.A1(\counter[0] ),
    .A2(_029_),
    .ZN(_046_));
 AOI21_X1 _210_ (.A(_027_),
    .B1(_045_),
    .B2(_046_),
    .ZN(_000_));
 NAND2_X1 _211_ (.A1(\counter[1] ),
    .A2(_029_),
    .ZN(_047_));
 INV_X1 _212_ (.A(_166_),
    .ZN(_048_));
 NOR3_X1 _213_ (.A1(_048_),
    .A2(_029_),
    .A3(_033_),
    .ZN(_049_));
 OAI21_X1 _214_ (.A(_049_),
    .B1(_043_),
    .B2(_044_),
    .ZN(_050_));
 AOI21_X1 _215_ (.A(_027_),
    .B1(_047_),
    .B2(_050_),
    .ZN(_001_));
 NAND2_X1 _216_ (.A1(\counter[2] ),
    .A2(_029_),
    .ZN(_051_));
 OR2_X1 _217_ (.A1(_032_),
    .A2(_031_),
    .ZN(_052_));
 AND2_X1 _218_ (.A1(_052_),
    .A2(_030_),
    .ZN(_053_));
 INV_X1 _219_ (.A(\counter[2] ),
    .ZN(_054_));
 AND3_X1 _220_ (.A1(_165_),
    .A2(_054_),
    .A3(_028_),
    .ZN(_055_));
 NOR2_X1 _221_ (.A1(_165_),
    .A2(_054_),
    .ZN(_056_));
 OAI221_X1 _222_ (.A(_053_),
    .B1(_055_),
    .B2(_056_),
    .C1(_043_),
    .C2(_044_),
    .ZN(_057_));
 AOI21_X1 _223_ (.A(_027_),
    .B1(_051_),
    .B2(_057_),
    .ZN(_002_));
 BUF_X2 _224_ (.A(\counter[3] ),
    .Z(_058_));
 NAND2_X1 _225_ (.A1(_058_),
    .A2(_029_),
    .ZN(_059_));
 NAND3_X1 _226_ (.A1(\counter[0] ),
    .A2(\counter[2] ),
    .A3(\counter[1] ),
    .ZN(_060_));
 NOR3_X1 _227_ (.A1(_058_),
    .A2(_029_),
    .A3(_060_),
    .ZN(_061_));
 AND2_X1 _228_ (.A1(_058_),
    .A2(_060_),
    .ZN(_062_));
 OAI221_X1 _229_ (.A(_053_),
    .B1(_061_),
    .B2(_062_),
    .C1(_043_),
    .C2(_044_),
    .ZN(_063_));
 AOI21_X1 _230_ (.A(_027_),
    .B1(_059_),
    .B2(_063_),
    .ZN(_003_));
 CLKBUF_X3 _231_ (.A(_025_),
    .Z(_064_));
 NAND4_X2 _232_ (.A1(_165_),
    .A2(\counter[2] ),
    .A3(_058_),
    .A4(_028_),
    .ZN(_065_));
 XNOR2_X1 _233_ (.A(\counter[4] ),
    .B(_065_),
    .ZN(_066_));
 NAND2_X1 _234_ (.A1(_064_),
    .A2(_066_),
    .ZN(_067_));
 OAI21_X2 _235_ (.A(_053_),
    .B1(_043_),
    .B2(_044_),
    .ZN(_068_));
 AOI21_X1 _236_ (.A(_067_),
    .B1(_068_),
    .B2(_028_),
    .ZN(_004_));
 NAND3_X1 _237_ (.A1(_058_),
    .A2(\counter[4] ),
    .A3(_028_),
    .ZN(_069_));
 NOR2_X1 _238_ (.A1(_060_),
    .A2(_069_),
    .ZN(_070_));
 XOR2_X1 _239_ (.A(\counter[5] ),
    .B(_070_),
    .Z(_071_));
 NAND2_X1 _240_ (.A1(_025_),
    .A2(_071_),
    .ZN(_072_));
 AOI21_X1 _241_ (.A(_072_),
    .B1(_068_),
    .B2(_028_),
    .ZN(_005_));
 NAND2_X1 _242_ (.A1(\counter[4] ),
    .A2(\counter[5] ),
    .ZN(_073_));
 NOR2_X1 _243_ (.A1(_065_),
    .A2(_073_),
    .ZN(_074_));
 XNOR2_X1 _244_ (.A(\counter[6] ),
    .B(_074_),
    .ZN(_075_));
 OR2_X1 _245_ (.A1(_026_),
    .A2(_075_),
    .ZN(_076_));
 AOI21_X1 _246_ (.A(_076_),
    .B1(_068_),
    .B2(_028_),
    .ZN(_006_));
 NAND3_X1 _247_ (.A1(\counter[5] ),
    .A2(\counter[6] ),
    .A3(_070_),
    .ZN(_077_));
 XOR2_X2 _248_ (.A(\counter[7] ),
    .B(_077_),
    .Z(_078_));
 AOI211_X2 _249_ (.A(_026_),
    .B(_078_),
    .C1(_068_),
    .C2(_028_),
    .ZN(_007_));
 NOR2_X4 _250_ (.A1(_044_),
    .A2(_036_),
    .ZN(_079_));
 CLKBUF_X3 _251_ (.A(_079_),
    .Z(_080_));
 NAND2_X1 _252_ (.A1(net1),
    .A2(_080_),
    .ZN(_081_));
 OR2_X1 _253_ (.A1(_044_),
    .A2(_036_),
    .ZN(_082_));
 BUF_X2 _254_ (.A(_082_),
    .Z(_083_));
 BUF_X4 _255_ (.A(_083_),
    .Z(_084_));
 NAND2_X1 _256_ (.A1(\duty_reg[0] ),
    .A2(_084_),
    .ZN(_085_));
 AOI21_X1 _257_ (.A(_027_),
    .B1(_081_),
    .B2(_085_),
    .ZN(_008_));
 NAND2_X1 _258_ (.A1(net2),
    .A2(_079_),
    .ZN(_086_));
 NAND2_X1 _259_ (.A1(\duty_reg[1] ),
    .A2(_083_),
    .ZN(_087_));
 AOI21_X1 _260_ (.A(_027_),
    .B1(_086_),
    .B2(_087_),
    .ZN(_009_));
 NAND2_X1 _261_ (.A1(net3),
    .A2(_079_),
    .ZN(_088_));
 NAND2_X1 _262_ (.A1(\duty_reg[2] ),
    .A2(_083_),
    .ZN(_089_));
 AOI21_X1 _263_ (.A(_027_),
    .B1(_088_),
    .B2(_089_),
    .ZN(_010_));
 NAND2_X1 _264_ (.A1(net4),
    .A2(_079_),
    .ZN(_090_));
 NAND2_X1 _265_ (.A1(\duty_reg[3] ),
    .A2(_083_),
    .ZN(_091_));
 AOI21_X1 _266_ (.A(_027_),
    .B1(_090_),
    .B2(_091_),
    .ZN(_011_));
 NAND2_X1 _267_ (.A1(net5),
    .A2(_079_),
    .ZN(_092_));
 NAND2_X1 _268_ (.A1(\duty_reg[4] ),
    .A2(_083_),
    .ZN(_093_));
 AOI21_X1 _269_ (.A(_027_),
    .B1(_092_),
    .B2(_093_),
    .ZN(_012_));
 NAND2_X1 _270_ (.A1(net6),
    .A2(_079_),
    .ZN(_094_));
 NAND2_X1 _271_ (.A1(\duty_reg[5] ),
    .A2(_083_),
    .ZN(_095_));
 AOI21_X1 _272_ (.A(_027_),
    .B1(_094_),
    .B2(_095_),
    .ZN(_013_));
 NAND2_X1 _273_ (.A1(net7),
    .A2(_079_),
    .ZN(_096_));
 NAND2_X1 _274_ (.A1(\duty_reg[6] ),
    .A2(_083_),
    .ZN(_097_));
 AOI21_X1 _275_ (.A(_026_),
    .B1(_096_),
    .B2(_097_),
    .ZN(_014_));
 NAND2_X1 _276_ (.A1(\duty_reg[7] ),
    .A2(_084_),
    .ZN(_098_));
 NAND2_X1 _277_ (.A1(net8),
    .A2(_080_),
    .ZN(_099_));
 NAND3_X1 _278_ (.A1(_064_),
    .A2(_098_),
    .A3(_099_),
    .ZN(_015_));
 NAND2_X1 _279_ (.A1(\period_reg[0] ),
    .A2(_084_),
    .ZN(_100_));
 NAND2_X1 _280_ (.A1(net9),
    .A2(_080_),
    .ZN(_101_));
 NAND3_X1 _281_ (.A1(_064_),
    .A2(_100_),
    .A3(_101_),
    .ZN(_016_));
 NAND2_X1 _282_ (.A1(\period_reg[1] ),
    .A2(_084_),
    .ZN(_102_));
 NAND2_X1 _283_ (.A1(net10),
    .A2(_080_),
    .ZN(_103_));
 NAND3_X1 _284_ (.A1(_064_),
    .A2(_102_),
    .A3(_103_),
    .ZN(_017_));
 NAND2_X1 _285_ (.A1(\period_reg[2] ),
    .A2(_084_),
    .ZN(_104_));
 NAND2_X1 _286_ (.A1(net11),
    .A2(_080_),
    .ZN(_105_));
 NAND3_X1 _287_ (.A1(_064_),
    .A2(_104_),
    .A3(_105_),
    .ZN(_018_));
 NAND2_X1 _288_ (.A1(\period_reg[3] ),
    .A2(_084_),
    .ZN(_106_));
 NAND2_X1 _289_ (.A1(net12),
    .A2(_080_),
    .ZN(_107_));
 NAND3_X1 _290_ (.A1(_064_),
    .A2(_106_),
    .A3(_107_),
    .ZN(_019_));
 NAND2_X1 _291_ (.A1(\period_reg[4] ),
    .A2(_084_),
    .ZN(_108_));
 NAND2_X1 _292_ (.A1(net13),
    .A2(_080_),
    .ZN(_109_));
 NAND3_X1 _293_ (.A1(_064_),
    .A2(_108_),
    .A3(_109_),
    .ZN(_020_));
 NAND2_X1 _294_ (.A1(\period_reg[5] ),
    .A2(_084_),
    .ZN(_110_));
 NAND2_X1 _295_ (.A1(net14),
    .A2(_080_),
    .ZN(_111_));
 NAND3_X1 _296_ (.A1(_064_),
    .A2(_110_),
    .A3(_111_),
    .ZN(_021_));
 NAND2_X1 _297_ (.A1(\period_reg[6] ),
    .A2(_084_),
    .ZN(_112_));
 NAND2_X1 _298_ (.A1(net15),
    .A2(_080_),
    .ZN(_113_));
 NAND3_X1 _299_ (.A1(_064_),
    .A2(_112_),
    .A3(_113_),
    .ZN(_022_));
 NAND2_X1 _300_ (.A1(\period_reg[7] ),
    .A2(_084_),
    .ZN(_114_));
 NAND2_X1 _301_ (.A1(net16),
    .A2(_080_),
    .ZN(_115_));
 NAND3_X1 _302_ (.A1(_064_),
    .A2(_114_),
    .A3(_115_),
    .ZN(_023_));
 NAND3_X1 _303_ (.A1(_181_),
    .A2(_175_),
    .A3(_178_),
    .ZN(_116_));
 INV_X1 _304_ (.A(_187_),
    .ZN(_117_));
 INV_X1 _305_ (.A(\counter[0] ),
    .ZN(_118_));
 AOI21_X1 _306_ (.A(_117_),
    .B1(\duty_reg[0] ),
    .B2(_118_),
    .ZN(_119_));
 OAI21_X1 _307_ (.A(_184_),
    .B1(_186_),
    .B2(_119_),
    .ZN(_120_));
 INV_X1 _308_ (.A(_183_),
    .ZN(_121_));
 AOI21_X1 _309_ (.A(_116_),
    .B1(_120_),
    .B2(_121_),
    .ZN(_122_));
 NAND2_X1 _310_ (.A1(_028_),
    .A2(_025_),
    .ZN(_123_));
 NOR4_X1 _311_ (.A1(_168_),
    .A2(_171_),
    .A3(_174_),
    .A4(_123_),
    .ZN(_124_));
 AOI21_X1 _312_ (.A(_177_),
    .B1(_178_),
    .B2(_180_),
    .ZN(_125_));
 INV_X1 _313_ (.A(_175_),
    .ZN(_126_));
 OAI21_X1 _314_ (.A(_124_),
    .B1(_125_),
    .B2(_126_),
    .ZN(_127_));
 OAI21_X1 _315_ (.A(_169_),
    .B1(_172_),
    .B2(_171_),
    .ZN(_128_));
 NOR2_X1 _316_ (.A1(_168_),
    .A2(_029_),
    .ZN(_129_));
 AOI22_X1 _317_ (.A1(_029_),
    .A2(net17),
    .B1(_128_),
    .B2(_129_),
    .ZN(_130_));
 OAI22_X1 _318_ (.A1(_122_),
    .A2(_127_),
    .B1(_130_),
    .B2(_026_),
    .ZN(_024_));
 HA_X1 _319_ (.A(_141_),
    .B(\period_reg[0] ),
    .CO(_142_),
    .S(_143_));
 HA_X1 _320_ (.A(\counter[1] ),
    .B(_144_),
    .CO(_145_),
    .S(_146_));
 HA_X1 _321_ (.A(\counter[3] ),
    .B(_147_),
    .CO(_148_),
    .S(_149_));
 HA_X1 _322_ (.A(\counter[2] ),
    .B(_150_),
    .CO(_151_),
    .S(_152_));
 HA_X1 _323_ (.A(\counter[7] ),
    .B(_153_),
    .CO(_154_),
    .S(_155_));
 HA_X1 _324_ (.A(\counter[6] ),
    .B(_156_),
    .CO(_157_),
    .S(_158_));
 HA_X1 _325_ (.A(\counter[5] ),
    .B(_159_),
    .CO(_160_),
    .S(_161_));
 HA_X1 _326_ (.A(\counter[4] ),
    .B(_162_),
    .CO(_163_),
    .S(_164_));
 HA_X1 _327_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .CO(_165_),
    .S(_166_));
 HA_X1 _328_ (.A(\counter[7] ),
    .B(_167_),
    .CO(_168_),
    .S(_169_));
 HA_X1 _329_ (.A(\counter[6] ),
    .B(_170_),
    .CO(_171_),
    .S(_172_));
 HA_X1 _330_ (.A(\counter[5] ),
    .B(_173_),
    .CO(_174_),
    .S(_175_));
 HA_X1 _331_ (.A(\counter[4] ),
    .B(_176_),
    .CO(_177_),
    .S(_178_));
 HA_X1 _332_ (.A(\counter[3] ),
    .B(_179_),
    .CO(_180_),
    .S(_181_));
 HA_X1 _333_ (.A(\counter[2] ),
    .B(_182_),
    .CO(_183_),
    .S(_184_));
 HA_X1 _334_ (.A(\counter[1] ),
    .B(_185_),
    .CO(_186_),
    .S(_187_));
 DFF_X2 \counter[0]$_SDFFE_PN0P_  (.D(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\counter[0] ),
    .QN(_141_));
 DFF_X2 \counter[1]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\counter[1] ),
    .QN(_140_));
 DFF_X2 \counter[2]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[2] ),
    .QN(_139_));
 DFF_X2 \counter[3]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[3] ),
    .QN(_138_));
 DFF_X2 \counter[4]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[4] ),
    .QN(_137_));
 DFF_X2 \counter[5]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[5] ),
    .QN(_136_));
 DFF_X2 \counter[6]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[6] ),
    .QN(_135_));
 DFF_X2 \counter[7]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[7] ),
    .QN(_134_));
 DFF_X1 \duty_reg[0]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[0] ),
    .QN(_133_));
 DFF_X1 \duty_reg[1]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[1] ),
    .QN(_185_));
 DFF_X1 \duty_reg[2]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[2] ),
    .QN(_182_));
 DFF_X1 \duty_reg[3]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[3] ),
    .QN(_179_));
 DFF_X1 \duty_reg[4]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[4] ),
    .QN(_176_));
 DFF_X1 \duty_reg[5]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[5] ),
    .QN(_173_));
 DFF_X1 \duty_reg[6]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[6] ),
    .QN(_170_));
 DFF_X1 \duty_reg[7]$_SDFFE_PN1P_  (.D(_015_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\duty_reg[7] ),
    .QN(_167_));
 DFF_X1 \period_reg[0]$_SDFFE_PN1P_  (.D(_016_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\period_reg[0] ),
    .QN(_132_));
 DFF_X1 \period_reg[1]$_SDFFE_PN1P_  (.D(_017_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\period_reg[1] ),
    .QN(_144_));
 DFF_X1 \period_reg[2]$_SDFFE_PN1P_  (.D(_018_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\period_reg[2] ),
    .QN(_150_));
 DFF_X1 \period_reg[3]$_SDFFE_PN1P_  (.D(_019_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\period_reg[3] ),
    .QN(_147_));
 DFF_X1 \period_reg[4]$_SDFFE_PN1P_  (.D(_020_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\period_reg[4] ),
    .QN(_162_));
 DFF_X1 \period_reg[5]$_SDFFE_PN1P_  (.D(_021_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\period_reg[5] ),
    .QN(_159_));
 DFF_X1 \period_reg[6]$_SDFFE_PN1P_  (.D(_022_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\period_reg[6] ),
    .QN(_156_));
 DFF_X1 \period_reg[7]$_SDFFE_PN1P_  (.D(_023_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\period_reg[7] ),
    .QN(_153_));
 DFF_X1 \pwm_out$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net17),
    .QN(_131_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_107 ();
 BUF_X1 input1 (.A(duty_cycle[0]),
    .Z(net1));
 BUF_X1 input2 (.A(duty_cycle[1]),
    .Z(net2));
 BUF_X1 input3 (.A(duty_cycle[2]),
    .Z(net3));
 BUF_X1 input4 (.A(duty_cycle[3]),
    .Z(net4));
 BUF_X1 input5 (.A(duty_cycle[4]),
    .Z(net5));
 BUF_X1 input6 (.A(duty_cycle[5]),
    .Z(net6));
 BUF_X1 input7 (.A(duty_cycle[6]),
    .Z(net7));
 BUF_X1 input8 (.A(duty_cycle[7]),
    .Z(net8));
 BUF_X1 input9 (.A(period[0]),
    .Z(net9));
 BUF_X1 input10 (.A(period[1]),
    .Z(net10));
 BUF_X1 input11 (.A(period[2]),
    .Z(net11));
 BUF_X1 input12 (.A(period[3]),
    .Z(net12));
 BUF_X1 input13 (.A(period[4]),
    .Z(net13));
 BUF_X1 input14 (.A(period[5]),
    .Z(net14));
 BUF_X1 input15 (.A(period[6]),
    .Z(net15));
 BUF_X1 input16 (.A(period[7]),
    .Z(net16));
 BUF_X1 output17 (.A(net17),
    .Z(pwm_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 INV_X2 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X16 FILLER_0_129 ();
 FILLCELL_X8 FILLER_0_145 ();
 FILLCELL_X2 FILLER_0_153 ();
 FILLCELL_X1 FILLER_0_155 ();
 FILLCELL_X8 FILLER_0_159 ();
 FILLCELL_X2 FILLER_0_167 ();
 FILLCELL_X1 FILLER_0_169 ();
 FILLCELL_X32 FILLER_0_173 ();
 FILLCELL_X32 FILLER_0_205 ();
 FILLCELL_X32 FILLER_0_237 ();
 FILLCELL_X32 FILLER_0_269 ();
 FILLCELL_X32 FILLER_0_301 ();
 FILLCELL_X32 FILLER_0_333 ();
 FILLCELL_X32 FILLER_0_365 ();
 FILLCELL_X4 FILLER_0_397 ();
 FILLCELL_X2 FILLER_0_401 ();
 FILLCELL_X1 FILLER_0_403 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X16 FILLER_1_385 ();
 FILLCELL_X2 FILLER_1_401 ();
 FILLCELL_X1 FILLER_1_403 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X16 FILLER_2_385 ();
 FILLCELL_X2 FILLER_2_401 ();
 FILLCELL_X1 FILLER_2_403 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X16 FILLER_3_385 ();
 FILLCELL_X2 FILLER_3_401 ();
 FILLCELL_X1 FILLER_3_403 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X16 FILLER_4_385 ();
 FILLCELL_X2 FILLER_4_401 ();
 FILLCELL_X1 FILLER_4_403 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X16 FILLER_5_385 ();
 FILLCELL_X2 FILLER_5_401 ();
 FILLCELL_X1 FILLER_5_403 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X16 FILLER_6_385 ();
 FILLCELL_X2 FILLER_6_401 ();
 FILLCELL_X1 FILLER_6_403 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X16 FILLER_7_385 ();
 FILLCELL_X2 FILLER_7_401 ();
 FILLCELL_X1 FILLER_7_403 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X16 FILLER_8_385 ();
 FILLCELL_X2 FILLER_8_401 ();
 FILLCELL_X1 FILLER_8_403 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X16 FILLER_9_385 ();
 FILLCELL_X2 FILLER_9_401 ();
 FILLCELL_X1 FILLER_9_403 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X16 FILLER_10_385 ();
 FILLCELL_X2 FILLER_10_401 ();
 FILLCELL_X1 FILLER_10_403 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X16 FILLER_11_385 ();
 FILLCELL_X2 FILLER_11_401 ();
 FILLCELL_X1 FILLER_11_403 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X16 FILLER_12_385 ();
 FILLCELL_X2 FILLER_12_401 ();
 FILLCELL_X1 FILLER_12_403 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X16 FILLER_13_385 ();
 FILLCELL_X2 FILLER_13_401 ();
 FILLCELL_X1 FILLER_13_403 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X16 FILLER_14_385 ();
 FILLCELL_X2 FILLER_14_401 ();
 FILLCELL_X1 FILLER_14_403 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X16 FILLER_15_385 ();
 FILLCELL_X2 FILLER_15_401 ();
 FILLCELL_X1 FILLER_15_403 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X16 FILLER_16_385 ();
 FILLCELL_X2 FILLER_16_401 ();
 FILLCELL_X1 FILLER_16_403 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X8 FILLER_17_225 ();
 FILLCELL_X2 FILLER_17_233 ();
 FILLCELL_X32 FILLER_17_242 ();
 FILLCELL_X32 FILLER_17_274 ();
 FILLCELL_X32 FILLER_17_306 ();
 FILLCELL_X32 FILLER_17_338 ();
 FILLCELL_X32 FILLER_17_370 ();
 FILLCELL_X2 FILLER_17_402 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X16 FILLER_18_385 ();
 FILLCELL_X2 FILLER_18_401 ();
 FILLCELL_X1 FILLER_18_403 ();
 FILLCELL_X16 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_17 ();
 FILLCELL_X2 FILLER_19_21 ();
 FILLCELL_X1 FILLER_19_23 ();
 FILLCELL_X32 FILLER_19_27 ();
 FILLCELL_X32 FILLER_19_59 ();
 FILLCELL_X32 FILLER_19_91 ();
 FILLCELL_X16 FILLER_19_123 ();
 FILLCELL_X8 FILLER_19_139 ();
 FILLCELL_X4 FILLER_19_147 ();
 FILLCELL_X1 FILLER_19_151 ();
 FILLCELL_X8 FILLER_19_155 ();
 FILLCELL_X4 FILLER_19_163 ();
 FILLCELL_X1 FILLER_19_167 ();
 FILLCELL_X32 FILLER_19_171 ();
 FILLCELL_X32 FILLER_19_203 ();
 FILLCELL_X32 FILLER_19_235 ();
 FILLCELL_X32 FILLER_19_267 ();
 FILLCELL_X32 FILLER_19_299 ();
 FILLCELL_X32 FILLER_19_331 ();
 FILLCELL_X32 FILLER_19_363 ();
 FILLCELL_X8 FILLER_19_395 ();
 FILLCELL_X1 FILLER_19_403 ();
 FILLCELL_X8 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_9 ();
 FILLCELL_X2 FILLER_20_16 ();
 FILLCELL_X1 FILLER_20_18 ();
 FILLCELL_X32 FILLER_20_22 ();
 FILLCELL_X4 FILLER_20_54 ();
 FILLCELL_X2 FILLER_20_61 ();
 FILLCELL_X1 FILLER_20_63 ();
 FILLCELL_X32 FILLER_20_67 ();
 FILLCELL_X32 FILLER_20_99 ();
 FILLCELL_X16 FILLER_20_131 ();
 FILLCELL_X4 FILLER_20_147 ();
 FILLCELL_X8 FILLER_20_155 ();
 FILLCELL_X2 FILLER_20_163 ();
 FILLCELL_X1 FILLER_20_165 ();
 FILLCELL_X8 FILLER_20_173 ();
 FILLCELL_X4 FILLER_20_181 ();
 FILLCELL_X1 FILLER_20_185 ();
 FILLCELL_X16 FILLER_20_203 ();
 FILLCELL_X4 FILLER_20_219 ();
 FILLCELL_X1 FILLER_20_223 ();
 FILLCELL_X32 FILLER_20_262 ();
 FILLCELL_X32 FILLER_20_294 ();
 FILLCELL_X32 FILLER_20_326 ();
 FILLCELL_X32 FILLER_20_358 ();
 FILLCELL_X8 FILLER_20_390 ();
 FILLCELL_X4 FILLER_20_398 ();
 FILLCELL_X2 FILLER_20_402 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X16 FILLER_21_33 ();
 FILLCELL_X8 FILLER_21_49 ();
 FILLCELL_X4 FILLER_21_57 ();
 FILLCELL_X1 FILLER_21_61 ();
 FILLCELL_X4 FILLER_21_66 ();
 FILLCELL_X1 FILLER_21_76 ();
 FILLCELL_X16 FILLER_21_98 ();
 FILLCELL_X8 FILLER_21_114 ();
 FILLCELL_X1 FILLER_21_122 ();
 FILLCELL_X8 FILLER_21_153 ();
 FILLCELL_X16 FILLER_21_187 ();
 FILLCELL_X4 FILLER_21_203 ();
 FILLCELL_X2 FILLER_21_222 ();
 FILLCELL_X1 FILLER_21_224 ();
 FILLCELL_X32 FILLER_21_242 ();
 FILLCELL_X32 FILLER_21_274 ();
 FILLCELL_X32 FILLER_21_306 ();
 FILLCELL_X32 FILLER_21_338 ();
 FILLCELL_X32 FILLER_21_370 ();
 FILLCELL_X2 FILLER_21_402 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X16 FILLER_22_33 ();
 FILLCELL_X8 FILLER_22_49 ();
 FILLCELL_X2 FILLER_22_57 ();
 FILLCELL_X16 FILLER_22_103 ();
 FILLCELL_X8 FILLER_22_119 ();
 FILLCELL_X1 FILLER_22_127 ();
 FILLCELL_X16 FILLER_22_148 ();
 FILLCELL_X8 FILLER_22_164 ();
 FILLCELL_X4 FILLER_22_172 ();
 FILLCELL_X2 FILLER_22_176 ();
 FILLCELL_X16 FILLER_22_190 ();
 FILLCELL_X2 FILLER_22_210 ();
 FILLCELL_X32 FILLER_22_231 ();
 FILLCELL_X32 FILLER_22_263 ();
 FILLCELL_X32 FILLER_22_295 ();
 FILLCELL_X32 FILLER_22_327 ();
 FILLCELL_X32 FILLER_22_359 ();
 FILLCELL_X8 FILLER_22_391 ();
 FILLCELL_X4 FILLER_22_399 ();
 FILLCELL_X1 FILLER_22_403 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_97 ();
 FILLCELL_X4 FILLER_23_113 ();
 FILLCELL_X1 FILLER_23_117 ();
 FILLCELL_X2 FILLER_23_139 ();
 FILLCELL_X1 FILLER_23_141 ();
 FILLCELL_X32 FILLER_23_146 ();
 FILLCELL_X8 FILLER_23_178 ();
 FILLCELL_X2 FILLER_23_186 ();
 FILLCELL_X1 FILLER_23_188 ();
 FILLCELL_X8 FILLER_23_194 ();
 FILLCELL_X1 FILLER_23_202 ();
 FILLCELL_X2 FILLER_23_212 ();
 FILLCELL_X8 FILLER_23_218 ();
 FILLCELL_X4 FILLER_23_226 ();
 FILLCELL_X2 FILLER_23_230 ();
 FILLCELL_X1 FILLER_23_232 ();
 FILLCELL_X2 FILLER_23_243 ();
 FILLCELL_X1 FILLER_23_245 ();
 FILLCELL_X32 FILLER_23_249 ();
 FILLCELL_X32 FILLER_23_281 ();
 FILLCELL_X32 FILLER_23_313 ();
 FILLCELL_X32 FILLER_23_345 ();
 FILLCELL_X16 FILLER_23_377 ();
 FILLCELL_X8 FILLER_23_393 ();
 FILLCELL_X2 FILLER_23_401 ();
 FILLCELL_X1 FILLER_23_403 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X16 FILLER_24_97 ();
 FILLCELL_X8 FILLER_24_113 ();
 FILLCELL_X1 FILLER_24_143 ();
 FILLCELL_X32 FILLER_24_148 ();
 FILLCELL_X32 FILLER_24_180 ();
 FILLCELL_X16 FILLER_24_212 ();
 FILLCELL_X4 FILLER_24_228 ();
 FILLCELL_X1 FILLER_24_232 ();
 FILLCELL_X2 FILLER_24_235 ();
 FILLCELL_X32 FILLER_24_240 ();
 FILLCELL_X32 FILLER_24_272 ();
 FILLCELL_X32 FILLER_24_304 ();
 FILLCELL_X32 FILLER_24_336 ();
 FILLCELL_X32 FILLER_24_368 ();
 FILLCELL_X4 FILLER_24_400 ();
 FILLCELL_X16 FILLER_25_1 ();
 FILLCELL_X8 FILLER_25_17 ();
 FILLCELL_X4 FILLER_25_25 ();
 FILLCELL_X32 FILLER_25_32 ();
 FILLCELL_X32 FILLER_25_64 ();
 FILLCELL_X32 FILLER_25_96 ();
 FILLCELL_X32 FILLER_25_128 ();
 FILLCELL_X16 FILLER_25_160 ();
 FILLCELL_X1 FILLER_25_176 ();
 FILLCELL_X32 FILLER_25_184 ();
 FILLCELL_X16 FILLER_25_216 ();
 FILLCELL_X8 FILLER_25_232 ();
 FILLCELL_X2 FILLER_25_240 ();
 FILLCELL_X32 FILLER_25_256 ();
 FILLCELL_X32 FILLER_25_288 ();
 FILLCELL_X32 FILLER_25_320 ();
 FILLCELL_X8 FILLER_25_352 ();
 FILLCELL_X4 FILLER_25_360 ();
 FILLCELL_X2 FILLER_25_364 ();
 FILLCELL_X32 FILLER_25_369 ();
 FILLCELL_X2 FILLER_25_401 ();
 FILLCELL_X1 FILLER_25_403 ();
 FILLCELL_X8 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_9 ();
 FILLCELL_X1 FILLER_26_11 ();
 FILLCELL_X32 FILLER_26_15 ();
 FILLCELL_X8 FILLER_26_47 ();
 FILLCELL_X1 FILLER_26_55 ();
 FILLCELL_X32 FILLER_26_86 ();
 FILLCELL_X32 FILLER_26_118 ();
 FILLCELL_X8 FILLER_26_150 ();
 FILLCELL_X4 FILLER_26_158 ();
 FILLCELL_X1 FILLER_26_162 ();
 FILLCELL_X1 FILLER_26_177 ();
 FILLCELL_X16 FILLER_26_194 ();
 FILLCELL_X8 FILLER_26_213 ();
 FILLCELL_X4 FILLER_26_221 ();
 FILLCELL_X2 FILLER_26_225 ();
 FILLCELL_X1 FILLER_26_227 ();
 FILLCELL_X32 FILLER_26_251 ();
 FILLCELL_X32 FILLER_26_283 ();
 FILLCELL_X32 FILLER_26_315 ();
 FILLCELL_X32 FILLER_26_347 ();
 FILLCELL_X16 FILLER_26_379 ();
 FILLCELL_X8 FILLER_26_395 ();
 FILLCELL_X1 FILLER_26_403 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X16 FILLER_27_33 ();
 FILLCELL_X8 FILLER_27_49 ();
 FILLCELL_X4 FILLER_27_57 ();
 FILLCELL_X8 FILLER_27_65 ();
 FILLCELL_X16 FILLER_27_76 ();
 FILLCELL_X4 FILLER_27_92 ();
 FILLCELL_X2 FILLER_27_96 ();
 FILLCELL_X1 FILLER_27_98 ();
 FILLCELL_X16 FILLER_27_109 ();
 FILLCELL_X4 FILLER_27_125 ();
 FILLCELL_X4 FILLER_27_147 ();
 FILLCELL_X1 FILLER_27_151 ();
 FILLCELL_X1 FILLER_27_165 ();
 FILLCELL_X2 FILLER_27_186 ();
 FILLCELL_X32 FILLER_27_191 ();
 FILLCELL_X8 FILLER_27_223 ();
 FILLCELL_X4 FILLER_27_231 ();
 FILLCELL_X2 FILLER_27_235 ();
 FILLCELL_X1 FILLER_27_237 ();
 FILLCELL_X1 FILLER_27_247 ();
 FILLCELL_X32 FILLER_27_265 ();
 FILLCELL_X32 FILLER_27_297 ();
 FILLCELL_X32 FILLER_27_329 ();
 FILLCELL_X32 FILLER_27_361 ();
 FILLCELL_X8 FILLER_27_393 ();
 FILLCELL_X2 FILLER_27_401 ();
 FILLCELL_X1 FILLER_27_403 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X16 FILLER_28_33 ();
 FILLCELL_X8 FILLER_28_49 ();
 FILLCELL_X1 FILLER_28_57 ();
 FILLCELL_X16 FILLER_28_75 ();
 FILLCELL_X8 FILLER_28_91 ();
 FILLCELL_X1 FILLER_28_99 ();
 FILLCELL_X4 FILLER_28_116 ();
 FILLCELL_X1 FILLER_28_120 ();
 FILLCELL_X8 FILLER_28_123 ();
 FILLCELL_X4 FILLER_28_131 ();
 FILLCELL_X1 FILLER_28_135 ();
 FILLCELL_X16 FILLER_28_144 ();
 FILLCELL_X2 FILLER_28_160 ();
 FILLCELL_X8 FILLER_28_171 ();
 FILLCELL_X2 FILLER_28_179 ();
 FILLCELL_X4 FILLER_28_185 ();
 FILLCELL_X2 FILLER_28_193 ();
 FILLCELL_X16 FILLER_28_200 ();
 FILLCELL_X8 FILLER_28_216 ();
 FILLCELL_X4 FILLER_28_224 ();
 FILLCELL_X2 FILLER_28_228 ();
 FILLCELL_X1 FILLER_28_230 ();
 FILLCELL_X2 FILLER_28_233 ();
 FILLCELL_X32 FILLER_28_240 ();
 FILLCELL_X32 FILLER_28_272 ();
 FILLCELL_X32 FILLER_28_304 ();
 FILLCELL_X32 FILLER_28_336 ();
 FILLCELL_X32 FILLER_28_368 ();
 FILLCELL_X4 FILLER_28_400 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X16 FILLER_29_65 ();
 FILLCELL_X8 FILLER_29_81 ();
 FILLCELL_X4 FILLER_29_89 ();
 FILLCELL_X1 FILLER_29_95 ();
 FILLCELL_X2 FILLER_29_134 ();
 FILLCELL_X8 FILLER_29_146 ();
 FILLCELL_X1 FILLER_29_154 ();
 FILLCELL_X16 FILLER_29_174 ();
 FILLCELL_X2 FILLER_29_190 ();
 FILLCELL_X1 FILLER_29_192 ();
 FILLCELL_X8 FILLER_29_212 ();
 FILLCELL_X4 FILLER_29_220 ();
 FILLCELL_X8 FILLER_29_238 ();
 FILLCELL_X1 FILLER_29_246 ();
 FILLCELL_X32 FILLER_29_251 ();
 FILLCELL_X32 FILLER_29_283 ();
 FILLCELL_X32 FILLER_29_315 ();
 FILLCELL_X32 FILLER_29_347 ();
 FILLCELL_X16 FILLER_29_379 ();
 FILLCELL_X8 FILLER_29_395 ();
 FILLCELL_X1 FILLER_29_403 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X1 FILLER_30_65 ();
 FILLCELL_X4 FILLER_30_86 ();
 FILLCELL_X2 FILLER_30_90 ();
 FILLCELL_X1 FILLER_30_115 ();
 FILLCELL_X1 FILLER_30_119 ();
 FILLCELL_X4 FILLER_30_143 ();
 FILLCELL_X1 FILLER_30_147 ();
 FILLCELL_X1 FILLER_30_157 ();
 FILLCELL_X32 FILLER_30_162 ();
 FILLCELL_X16 FILLER_30_194 ();
 FILLCELL_X8 FILLER_30_210 ();
 FILLCELL_X4 FILLER_30_218 ();
 FILLCELL_X4 FILLER_30_236 ();
 FILLCELL_X1 FILLER_30_240 ();
 FILLCELL_X32 FILLER_30_258 ();
 FILLCELL_X32 FILLER_30_290 ();
 FILLCELL_X32 FILLER_30_322 ();
 FILLCELL_X32 FILLER_30_354 ();
 FILLCELL_X16 FILLER_30_386 ();
 FILLCELL_X2 FILLER_30_402 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X16 FILLER_31_33 ();
 FILLCELL_X8 FILLER_31_49 ();
 FILLCELL_X4 FILLER_31_57 ();
 FILLCELL_X1 FILLER_31_61 ();
 FILLCELL_X32 FILLER_31_86 ();
 FILLCELL_X8 FILLER_31_118 ();
 FILLCELL_X4 FILLER_31_126 ();
 FILLCELL_X1 FILLER_31_130 ();
 FILLCELL_X8 FILLER_31_150 ();
 FILLCELL_X4 FILLER_31_158 ();
 FILLCELL_X1 FILLER_31_162 ();
 FILLCELL_X1 FILLER_31_167 ();
 FILLCELL_X16 FILLER_31_170 ();
 FILLCELL_X8 FILLER_31_186 ();
 FILLCELL_X1 FILLER_31_194 ();
 FILLCELL_X2 FILLER_31_205 ();
 FILLCELL_X32 FILLER_31_213 ();
 FILLCELL_X2 FILLER_31_245 ();
 FILLCELL_X1 FILLER_31_247 ();
 FILLCELL_X32 FILLER_31_254 ();
 FILLCELL_X32 FILLER_31_286 ();
 FILLCELL_X32 FILLER_31_318 ();
 FILLCELL_X16 FILLER_31_350 ();
 FILLCELL_X32 FILLER_31_369 ();
 FILLCELL_X2 FILLER_31_401 ();
 FILLCELL_X1 FILLER_31_403 ();
 FILLCELL_X16 FILLER_32_1 ();
 FILLCELL_X1 FILLER_32_20 ();
 FILLCELL_X32 FILLER_32_24 ();
 FILLCELL_X8 FILLER_32_56 ();
 FILLCELL_X2 FILLER_32_64 ();
 FILLCELL_X1 FILLER_32_66 ();
 FILLCELL_X4 FILLER_32_74 ();
 FILLCELL_X2 FILLER_32_78 ();
 FILLCELL_X32 FILLER_32_83 ();
 FILLCELL_X32 FILLER_32_115 ();
 FILLCELL_X16 FILLER_32_147 ();
 FILLCELL_X2 FILLER_32_176 ();
 FILLCELL_X4 FILLER_32_188 ();
 FILLCELL_X32 FILLER_32_196 ();
 FILLCELL_X32 FILLER_32_228 ();
 FILLCELL_X32 FILLER_32_260 ();
 FILLCELL_X32 FILLER_32_292 ();
 FILLCELL_X32 FILLER_32_324 ();
 FILLCELL_X32 FILLER_32_356 ();
 FILLCELL_X16 FILLER_32_388 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X2 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_166 ();
 FILLCELL_X32 FILLER_33_198 ();
 FILLCELL_X2 FILLER_33_230 ();
 FILLCELL_X1 FILLER_33_232 ();
 FILLCELL_X32 FILLER_33_250 ();
 FILLCELL_X32 FILLER_33_282 ();
 FILLCELL_X32 FILLER_33_314 ();
 FILLCELL_X32 FILLER_33_346 ();
 FILLCELL_X16 FILLER_33_378 ();
 FILLCELL_X8 FILLER_33_394 ();
 FILLCELL_X2 FILLER_33_402 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X16 FILLER_34_129 ();
 FILLCELL_X8 FILLER_34_145 ();
 FILLCELL_X1 FILLER_34_153 ();
 FILLCELL_X1 FILLER_34_159 ();
 FILLCELL_X32 FILLER_34_177 ();
 FILLCELL_X8 FILLER_34_209 ();
 FILLCELL_X4 FILLER_34_217 ();
 FILLCELL_X2 FILLER_34_221 ();
 FILLCELL_X2 FILLER_34_240 ();
 FILLCELL_X32 FILLER_34_252 ();
 FILLCELL_X32 FILLER_34_284 ();
 FILLCELL_X32 FILLER_34_316 ();
 FILLCELL_X16 FILLER_34_348 ();
 FILLCELL_X8 FILLER_34_364 ();
 FILLCELL_X16 FILLER_34_375 ();
 FILLCELL_X8 FILLER_34_391 ();
 FILLCELL_X4 FILLER_34_399 ();
 FILLCELL_X1 FILLER_34_403 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X4 FILLER_35_161 ();
 FILLCELL_X4 FILLER_35_189 ();
 FILLCELL_X2 FILLER_35_217 ();
 FILLCELL_X1 FILLER_35_219 ();
 FILLCELL_X32 FILLER_35_243 ();
 FILLCELL_X32 FILLER_35_275 ();
 FILLCELL_X32 FILLER_35_307 ();
 FILLCELL_X32 FILLER_35_339 ();
 FILLCELL_X32 FILLER_35_371 ();
 FILLCELL_X1 FILLER_35_403 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X4 FILLER_36_161 ();
 FILLCELL_X2 FILLER_36_165 ();
 FILLCELL_X1 FILLER_36_167 ();
 FILLCELL_X4 FILLER_36_171 ();
 FILLCELL_X2 FILLER_36_175 ();
 FILLCELL_X1 FILLER_36_177 ();
 FILLCELL_X32 FILLER_36_182 ();
 FILLCELL_X16 FILLER_36_214 ();
 FILLCELL_X2 FILLER_36_230 ();
 FILLCELL_X2 FILLER_36_236 ();
 FILLCELL_X32 FILLER_36_245 ();
 FILLCELL_X32 FILLER_36_277 ();
 FILLCELL_X32 FILLER_36_309 ();
 FILLCELL_X32 FILLER_36_341 ();
 FILLCELL_X16 FILLER_36_373 ();
 FILLCELL_X8 FILLER_36_389 ();
 FILLCELL_X4 FILLER_36_397 ();
 FILLCELL_X2 FILLER_36_401 ();
 FILLCELL_X1 FILLER_36_403 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X16 FILLER_37_161 ();
 FILLCELL_X4 FILLER_37_177 ();
 FILLCELL_X32 FILLER_37_184 ();
 FILLCELL_X8 FILLER_37_219 ();
 FILLCELL_X4 FILLER_37_227 ();
 FILLCELL_X2 FILLER_37_231 ();
 FILLCELL_X1 FILLER_37_233 ();
 FILLCELL_X32 FILLER_37_237 ();
 FILLCELL_X32 FILLER_37_269 ();
 FILLCELL_X32 FILLER_37_301 ();
 FILLCELL_X32 FILLER_37_333 ();
 FILLCELL_X32 FILLER_37_365 ();
 FILLCELL_X4 FILLER_37_397 ();
 FILLCELL_X2 FILLER_37_401 ();
 FILLCELL_X1 FILLER_37_403 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X16 FILLER_38_385 ();
 FILLCELL_X2 FILLER_38_401 ();
 FILLCELL_X1 FILLER_38_403 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X16 FILLER_39_385 ();
 FILLCELL_X2 FILLER_39_401 ();
 FILLCELL_X1 FILLER_39_403 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X16 FILLER_40_385 ();
 FILLCELL_X2 FILLER_40_401 ();
 FILLCELL_X1 FILLER_40_403 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X16 FILLER_41_385 ();
 FILLCELL_X2 FILLER_41_401 ();
 FILLCELL_X1 FILLER_41_403 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X16 FILLER_42_385 ();
 FILLCELL_X2 FILLER_42_401 ();
 FILLCELL_X1 FILLER_42_403 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X16 FILLER_43_385 ();
 FILLCELL_X2 FILLER_43_401 ();
 FILLCELL_X1 FILLER_43_403 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X16 FILLER_44_385 ();
 FILLCELL_X2 FILLER_44_401 ();
 FILLCELL_X1 FILLER_44_403 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X16 FILLER_45_385 ();
 FILLCELL_X2 FILLER_45_401 ();
 FILLCELL_X1 FILLER_45_403 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X16 FILLER_46_385 ();
 FILLCELL_X2 FILLER_46_401 ();
 FILLCELL_X1 FILLER_46_403 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X16 FILLER_47_385 ();
 FILLCELL_X2 FILLER_47_401 ();
 FILLCELL_X1 FILLER_47_403 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X16 FILLER_48_385 ();
 FILLCELL_X2 FILLER_48_401 ();
 FILLCELL_X1 FILLER_48_403 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X16 FILLER_49_385 ();
 FILLCELL_X2 FILLER_49_401 ();
 FILLCELL_X1 FILLER_49_403 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X16 FILLER_50_385 ();
 FILLCELL_X2 FILLER_50_401 ();
 FILLCELL_X1 FILLER_50_403 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X16 FILLER_51_385 ();
 FILLCELL_X2 FILLER_51_401 ();
 FILLCELL_X1 FILLER_51_403 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X16 FILLER_52_385 ();
 FILLCELL_X2 FILLER_52_401 ();
 FILLCELL_X1 FILLER_52_403 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X8 FILLER_53_161 ();
 FILLCELL_X4 FILLER_53_169 ();
 FILLCELL_X2 FILLER_53_173 ();
 FILLCELL_X1 FILLER_53_175 ();
 FILLCELL_X4 FILLER_53_179 ();
 FILLCELL_X32 FILLER_53_186 ();
 FILLCELL_X16 FILLER_53_221 ();
 FILLCELL_X2 FILLER_53_237 ();
 FILLCELL_X32 FILLER_53_245 ();
 FILLCELL_X32 FILLER_53_277 ();
 FILLCELL_X32 FILLER_53_309 ();
 FILLCELL_X32 FILLER_53_341 ();
 FILLCELL_X16 FILLER_53_373 ();
 FILLCELL_X8 FILLER_53_389 ();
 FILLCELL_X4 FILLER_53_397 ();
 FILLCELL_X2 FILLER_53_401 ();
 FILLCELL_X1 FILLER_53_403 ();
endmodule
