module performance_counter (clear,
    clk,
    enable,
    rst_n,
    all_counts,
    count_value,
    counter_sel,
    event_inc);
 input clear;
 input clk;
 input enable;
 input rst_n;
 output [255:0] all_counts;
 output [31:0] count_value;
 input [7:0] counter_sel;
 input [7:0] event_inc;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire \prev_event_inc[0] ;
 wire \prev_event_inc[1] ;
 wire \prev_event_inc[2] ;
 wire \prev_event_inc[3] ;
 wire \prev_event_inc[4] ;
 wire \prev_event_inc[5] ;
 wire \prev_event_inc[6] ;
 wire \prev_event_inc[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;

 sky130_fd_sc_hd__clkbuf_2 _1554_ (.A(clear),
    .X(_1215_));
 sky130_fd_sc_hd__buf_6 _1555_ (.A(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__buf_4 _1556_ (.A(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__clkbuf_4 _1557_ (.A(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__buf_4 _1558_ (.A(net4),
    .X(_1219_));
 sky130_fd_sc_hd__clkbuf_8 _1559_ (.A(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__and3b_1 _1560_ (.A_N(\prev_event_inc[0] ),
    .B(net5),
    .C(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__xnor2_1 _1561_ (.A(net14),
    .B(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__nor2_1 _1562_ (.A(_1218_),
    .B(_1222_),
    .Y(_0000_));
 sky130_fd_sc_hd__and4b_2 _1563_ (.A_N(\prev_event_inc[3] ),
    .B(net267),
    .C(_1219_),
    .D(net8),
    .X(_1223_));
 sky130_fd_sc_hd__and2_0 _1564_ (.A(net268),
    .B(_1550_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_2 _1565_ (.A(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__nand2_2 _1566_ (.A(_1223_),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__xor2_1 _1567_ (.A(net15),
    .B(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__nor2_1 _1568_ (.A(_1218_),
    .B(_1227_),
    .Y(_0001_));
 sky130_fd_sc_hd__buf_2 _1569_ (.A(_1223_),
    .X(_1228_));
 sky130_fd_sc_hd__and3_1 _1570_ (.A(net265),
    .B(net266),
    .C(net268),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_2 _1571_ (.A(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__nand3_1 _1572_ (.A(net15),
    .B(_1228_),
    .C(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__xor2_1 _1573_ (.A(net16),
    .B(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__nor2_1 _1574_ (.A(_1218_),
    .B(_1232_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand4_1 _1575_ (.A(net15),
    .B(net16),
    .C(_1228_),
    .D(_1225_),
    .Y(_1233_));
 sky130_fd_sc_hd__xor2_1 _1576_ (.A(net17),
    .B(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__nor2_1 _1577_ (.A(_1218_),
    .B(_1234_),
    .Y(_0003_));
 sky130_fd_sc_hd__and3_1 _1578_ (.A(net15),
    .B(net16),
    .C(net17),
    .X(_1235_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1579_ (.A(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__nand3_1 _1580_ (.A(_1228_),
    .B(_1230_),
    .C(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__xor2_1 _1581_ (.A(net18),
    .B(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__nor2_1 _1582_ (.A(_1218_),
    .B(_1238_),
    .Y(_0004_));
 sky130_fd_sc_hd__nand4_1 _1583_ (.A(net18),
    .B(_1228_),
    .C(_1225_),
    .D(_1236_),
    .Y(_1239_));
 sky130_fd_sc_hd__xor2_1 _1584_ (.A(net19),
    .B(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__nor2_1 _1585_ (.A(_1218_),
    .B(_1240_),
    .Y(_0005_));
 sky130_fd_sc_hd__and2_0 _1586_ (.A(net18),
    .B(net19),
    .X(_1241_));
 sky130_fd_sc_hd__and4_1 _1587_ (.A(_1228_),
    .B(_1230_),
    .C(_1236_),
    .D(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__xnor2_1 _1588_ (.A(net20),
    .B(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__nor2_1 _1589_ (.A(_1218_),
    .B(_1243_),
    .Y(_0006_));
 sky130_fd_sc_hd__and3_1 _1590_ (.A(net18),
    .B(net19),
    .C(net20),
    .X(_1244_));
 sky130_fd_sc_hd__nand4_1 _1591_ (.A(_1228_),
    .B(_1225_),
    .C(_1236_),
    .D(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__xor2_1 _1592_ (.A(net21),
    .B(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__nor2_1 _1593_ (.A(_1218_),
    .B(_1246_),
    .Y(_0007_));
 sky130_fd_sc_hd__and4_2 _1594_ (.A(net18),
    .B(net19),
    .C(net20),
    .D(net21),
    .X(_1247_));
 sky130_fd_sc_hd__nand4_1 _1595_ (.A(_1228_),
    .B(_1230_),
    .C(_1236_),
    .D(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__xor2_1 _1596_ (.A(net22),
    .B(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__nor2_1 _1597_ (.A(_1218_),
    .B(_1249_),
    .Y(_0008_));
 sky130_fd_sc_hd__nand3_1 _1598_ (.A(_1228_),
    .B(_1225_),
    .C(_1236_),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2_1 _1599_ (.A(net22),
    .B(_1247_),
    .Y(_1251_));
 sky130_fd_sc_hd__o21ai_0 _1600_ (.A1(_1250_),
    .A2(_1251_),
    .B1(net23),
    .Y(_1252_));
 sky130_fd_sc_hd__or3_1 _1601_ (.A(net23),
    .B(_1250_),
    .C(_1251_),
    .X(_1253_));
 sky130_fd_sc_hd__buf_4 _1602_ (.A(_1215_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_4 _1603_ (.A(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__a21oi_1 _1604_ (.A1(_1252_),
    .A2(_1253_),
    .B1(_1255_),
    .Y(_0009_));
 sky130_fd_sc_hd__and2_1 _1605_ (.A(net22),
    .B(net23),
    .X(_1256_));
 sky130_fd_sc_hd__nand2_2 _1606_ (.A(_1247_),
    .B(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__o21ai_0 _1607_ (.A1(_1237_),
    .A2(_1257_),
    .B1(net24),
    .Y(_1258_));
 sky130_fd_sc_hd__or3_1 _1608_ (.A(net24),
    .B(_1237_),
    .C(_1257_),
    .X(_1259_));
 sky130_fd_sc_hd__a21oi_1 _1609_ (.A1(_1258_),
    .A2(_1259_),
    .B1(_1255_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_1 _1610_ (.A(net269),
    .Y(_1260_));
 sky130_fd_sc_hd__inv_1 _1611_ (.A(_1540_),
    .Y(_1261_));
 sky130_fd_sc_hd__nand4b_2 _1612_ (.A_N(\prev_event_inc[0] ),
    .B(net192),
    .C(net4),
    .D(net5),
    .Y(_1262_));
 sky130_fd_sc_hd__nand4_2 _1613_ (.A(net203),
    .B(net214),
    .C(net225),
    .D(net236),
    .Y(_1263_));
 sky130_fd_sc_hd__nand2_1 _1614_ (.A(net247),
    .B(net258),
    .Y(_1264_));
 sky130_fd_sc_hd__or4_1 _1615_ (.A(_1261_),
    .B(_1262_),
    .C(_1263_),
    .D(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__clkbuf_4 _1616_ (.A(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__o21ai_0 _1617_ (.A1(_1260_),
    .A2(_1266_),
    .B1(net25),
    .Y(_1267_));
 sky130_fd_sc_hd__or3_1 _1618_ (.A(_1260_),
    .B(net25),
    .C(_1266_),
    .X(_1268_));
 sky130_fd_sc_hd__a21oi_1 _1619_ (.A1(_1267_),
    .A2(_1268_),
    .B1(_1255_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_1 _1620_ (.A(net24),
    .Y(_1269_));
 sky130_fd_sc_hd__o31ai_1 _1621_ (.A1(_1269_),
    .A2(_1250_),
    .A3(_1257_),
    .B1(net26),
    .Y(_1270_));
 sky130_fd_sc_hd__or4_1 _1622_ (.A(_1269_),
    .B(net26),
    .C(_1250_),
    .D(_1257_),
    .X(_1271_));
 sky130_fd_sc_hd__a21oi_1 _1623_ (.A1(_1270_),
    .A2(_1271_),
    .B1(_1255_),
    .Y(_0012_));
 sky130_fd_sc_hd__nand2_1 _1624_ (.A(_1228_),
    .B(_1230_),
    .Y(_1272_));
 sky130_fd_sc_hd__and4_2 _1625_ (.A(net15),
    .B(net16),
    .C(net17),
    .D(net26),
    .X(_1273_));
 sky130_fd_sc_hd__nand4_4 _1626_ (.A(net24),
    .B(_1247_),
    .C(_1256_),
    .D(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__o21ai_0 _1627_ (.A1(_1272_),
    .A2(_1274_),
    .B1(net27),
    .Y(_1275_));
 sky130_fd_sc_hd__or3_1 _1628_ (.A(net27),
    .B(_1272_),
    .C(_1274_),
    .X(_1276_));
 sky130_fd_sc_hd__a21oi_1 _1629_ (.A1(_1275_),
    .A2(_1276_),
    .B1(_1255_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_1 _1630_ (.A(net27),
    .Y(_1277_));
 sky130_fd_sc_hd__nand4_2 _1631_ (.A(net24),
    .B(_1223_),
    .C(_1225_),
    .D(_1273_),
    .Y(_1278_));
 sky130_fd_sc_hd__buf_2 _1632_ (.A(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__o31ai_1 _1633_ (.A1(_1277_),
    .A2(_1257_),
    .A3(_1279_),
    .B1(net28),
    .Y(_1280_));
 sky130_fd_sc_hd__or4_1 _1634_ (.A(_1277_),
    .B(net28),
    .C(_1257_),
    .D(_1279_),
    .X(_1281_));
 sky130_fd_sc_hd__a21oi_1 _1635_ (.A1(_1280_),
    .A2(_1281_),
    .B1(_1255_),
    .Y(_0014_));
 sky130_fd_sc_hd__nand4_4 _1636_ (.A(net24),
    .B(_1223_),
    .C(_1230_),
    .D(_1273_),
    .Y(_1282_));
 sky130_fd_sc_hd__buf_2 _1637_ (.A(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__nand2_1 _1638_ (.A(net27),
    .B(net28),
    .Y(_1284_));
 sky130_fd_sc_hd__o31ai_1 _1639_ (.A1(_1257_),
    .A2(_1283_),
    .A3(_1284_),
    .B1(net29),
    .Y(_1285_));
 sky130_fd_sc_hd__or4_1 _1640_ (.A(net29),
    .B(_1257_),
    .C(_1283_),
    .D(_1284_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_4 _1641_ (.A(_1216_),
    .X(_1287_));
 sky130_fd_sc_hd__buf_4 _1642_ (.A(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__a21oi_1 _1643_ (.A1(_1285_),
    .A2(_1286_),
    .B1(_1288_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand3_1 _1644_ (.A(net27),
    .B(net28),
    .C(net29),
    .Y(_1289_));
 sky130_fd_sc_hd__o31ai_1 _1645_ (.A1(_1226_),
    .A2(_1274_),
    .A3(_1289_),
    .B1(net30),
    .Y(_1290_));
 sky130_fd_sc_hd__or4_1 _1646_ (.A(net30),
    .B(_1226_),
    .C(_1274_),
    .D(_1289_),
    .X(_1291_));
 sky130_fd_sc_hd__a21oi_1 _1647_ (.A1(_1290_),
    .A2(_1291_),
    .B1(_1288_),
    .Y(_0016_));
 sky130_fd_sc_hd__nand4_1 _1648_ (.A(net27),
    .B(net28),
    .C(net29),
    .D(net30),
    .Y(_1292_));
 sky130_fd_sc_hd__o31ai_1 _1649_ (.A1(_1272_),
    .A2(_1274_),
    .A3(_1292_),
    .B1(net31),
    .Y(_1293_));
 sky130_fd_sc_hd__or4_1 _1650_ (.A(net31),
    .B(_1272_),
    .C(_1274_),
    .D(_1292_),
    .X(_1294_));
 sky130_fd_sc_hd__a21oi_1 _1651_ (.A1(_1293_),
    .A2(_1294_),
    .B1(_1288_),
    .Y(_0017_));
 sky130_fd_sc_hd__and4_1 _1652_ (.A(net27),
    .B(net28),
    .C(net29),
    .D(net30),
    .X(_1295_));
 sky130_fd_sc_hd__nand2_1 _1653_ (.A(net31),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__o31ai_1 _1654_ (.A1(_1226_),
    .A2(_1274_),
    .A3(_1296_),
    .B1(net32),
    .Y(_1297_));
 sky130_fd_sc_hd__or4_1 _1655_ (.A(net32),
    .B(_1226_),
    .C(_1274_),
    .D(_1296_),
    .X(_1298_));
 sky130_fd_sc_hd__a21oi_1 _1656_ (.A1(_1297_),
    .A2(_1298_),
    .B1(_1288_),
    .Y(_0018_));
 sky130_fd_sc_hd__and2_0 _1657_ (.A(net31),
    .B(net32),
    .X(_1299_));
 sky130_fd_sc_hd__nand4_2 _1658_ (.A(_1247_),
    .B(_1256_),
    .C(_1295_),
    .D(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__clkbuf_2 _1659_ (.A(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__buf_2 _1660_ (.A(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__o21ai_0 _1661_ (.A1(_1283_),
    .A2(_1302_),
    .B1(net33),
    .Y(_1303_));
 sky130_fd_sc_hd__or3_1 _1662_ (.A(net33),
    .B(_1283_),
    .C(_1301_),
    .X(_1304_));
 sky130_fd_sc_hd__a21oi_1 _1663_ (.A1(_1303_),
    .A2(_1304_),
    .B1(_1288_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_1 _1664_ (.A(net33),
    .Y(_1305_));
 sky130_fd_sc_hd__o31ai_1 _1665_ (.A1(_1305_),
    .A2(_1279_),
    .A3(_1302_),
    .B1(net34),
    .Y(_1306_));
 sky130_fd_sc_hd__or4_1 _1666_ (.A(_1305_),
    .B(net34),
    .C(_1279_),
    .D(_1301_),
    .X(_1307_));
 sky130_fd_sc_hd__a21oi_1 _1667_ (.A1(_1306_),
    .A2(_1307_),
    .B1(_1288_),
    .Y(_0020_));
 sky130_fd_sc_hd__nand2_1 _1668_ (.A(net33),
    .B(net34),
    .Y(_1308_));
 sky130_fd_sc_hd__o31ai_1 _1669_ (.A1(_1283_),
    .A2(_1302_),
    .A3(_1308_),
    .B1(net35),
    .Y(_1309_));
 sky130_fd_sc_hd__or4_1 _1670_ (.A(net35),
    .B(_1283_),
    .C(_1301_),
    .D(_1308_),
    .X(_1310_));
 sky130_fd_sc_hd__a21oi_1 _1671_ (.A1(_1309_),
    .A2(_1310_),
    .B1(_1288_),
    .Y(_0021_));
 sky130_fd_sc_hd__and4_1 _1672_ (.A(net203),
    .B(net214),
    .C(net225),
    .D(net236),
    .X(_1311_));
 sky130_fd_sc_hd__nand3_1 _1673_ (.A(net247),
    .B(net258),
    .C(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__nand2_1 _1674_ (.A(net269),
    .B(net25),
    .Y(_1313_));
 sky130_fd_sc_hd__and4b_1 _1675_ (.A_N(\prev_event_inc[0] ),
    .B(net192),
    .C(_1219_),
    .D(net5),
    .X(_1314_));
 sky130_fd_sc_hd__nand3_1 _1676_ (.A(net14),
    .B(net125),
    .C(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__o31ai_1 _1677_ (.A1(_1312_),
    .A2(_1313_),
    .A3(_1315_),
    .B1(net36),
    .Y(_1316_));
 sky130_fd_sc_hd__or4_1 _1678_ (.A(net36),
    .B(_1312_),
    .C(_1313_),
    .D(_1315_),
    .X(_1317_));
 sky130_fd_sc_hd__a21oi_1 _1679_ (.A1(_1316_),
    .A2(_1317_),
    .B1(_1288_),
    .Y(_0022_));
 sky130_fd_sc_hd__nand3_1 _1680_ (.A(net33),
    .B(net34),
    .C(net35),
    .Y(_1318_));
 sky130_fd_sc_hd__o31ai_1 _1681_ (.A1(_1279_),
    .A2(_1302_),
    .A3(_1318_),
    .B1(net37),
    .Y(_1319_));
 sky130_fd_sc_hd__or4_1 _1682_ (.A(net37),
    .B(_1279_),
    .C(_1301_),
    .D(_1318_),
    .X(_1320_));
 sky130_fd_sc_hd__a21oi_1 _1683_ (.A1(_1319_),
    .A2(_1320_),
    .B1(_1288_),
    .Y(_0023_));
 sky130_fd_sc_hd__nand4_1 _1684_ (.A(net33),
    .B(net34),
    .C(net35),
    .D(net37),
    .Y(_1321_));
 sky130_fd_sc_hd__o31ai_1 _1685_ (.A1(_1283_),
    .A2(_1302_),
    .A3(_1321_),
    .B1(net38),
    .Y(_1322_));
 sky130_fd_sc_hd__or4_1 _1686_ (.A(net38),
    .B(_1282_),
    .C(_1301_),
    .D(_1321_),
    .X(_1323_));
 sky130_fd_sc_hd__a21oi_1 _1687_ (.A1(_1322_),
    .A2(_1323_),
    .B1(_1288_),
    .Y(_0024_));
 sky130_fd_sc_hd__and4_1 _1688_ (.A(net33),
    .B(net34),
    .C(net35),
    .D(net37),
    .X(_1324_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1689_ (.A(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__nand2_1 _1690_ (.A(net38),
    .B(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__o31ai_1 _1691_ (.A1(_1279_),
    .A2(_1302_),
    .A3(_1326_),
    .B1(net39),
    .Y(_1327_));
 sky130_fd_sc_hd__or4_1 _1692_ (.A(net39),
    .B(_1279_),
    .C(_1301_),
    .D(_1326_),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_4 _1693_ (.A(_1287_),
    .X(_1329_));
 sky130_fd_sc_hd__a21oi_1 _1694_ (.A1(_1327_),
    .A2(_1328_),
    .B1(_1329_),
    .Y(_0025_));
 sky130_fd_sc_hd__nand3_1 _1695_ (.A(net38),
    .B(net39),
    .C(_1325_),
    .Y(_1330_));
 sky130_fd_sc_hd__o31ai_1 _1696_ (.A1(_1283_),
    .A2(_1302_),
    .A3(_1330_),
    .B1(net40),
    .Y(_1331_));
 sky130_fd_sc_hd__or4_1 _1697_ (.A(net40),
    .B(_1282_),
    .C(_1301_),
    .D(_1330_),
    .X(_1332_));
 sky130_fd_sc_hd__a21oi_1 _1698_ (.A1(_1331_),
    .A2(_1332_),
    .B1(_1329_),
    .Y(_0026_));
 sky130_fd_sc_hd__nand4_1 _1699_ (.A(net38),
    .B(net39),
    .C(net40),
    .D(_1325_),
    .Y(_1333_));
 sky130_fd_sc_hd__o31ai_1 _1700_ (.A1(_1279_),
    .A2(_1302_),
    .A3(_1333_),
    .B1(net41),
    .Y(_1334_));
 sky130_fd_sc_hd__or4_1 _1701_ (.A(net41),
    .B(_1278_),
    .C(_1301_),
    .D(_1333_),
    .X(_1335_));
 sky130_fd_sc_hd__a21oi_1 _1702_ (.A1(_1334_),
    .A2(_1335_),
    .B1(_1329_),
    .Y(_0027_));
 sky130_fd_sc_hd__and4_1 _1703_ (.A(net38),
    .B(net39),
    .C(net40),
    .D(net41),
    .X(_1336_));
 sky130_fd_sc_hd__nand2_1 _1704_ (.A(_1325_),
    .B(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__o31ai_1 _1705_ (.A1(_1283_),
    .A2(_1302_),
    .A3(_1337_),
    .B1(net42),
    .Y(_1338_));
 sky130_fd_sc_hd__or4_1 _1706_ (.A(net42),
    .B(_1282_),
    .C(_1300_),
    .D(_1337_),
    .X(_1339_));
 sky130_fd_sc_hd__a21oi_1 _1707_ (.A1(_1338_),
    .A2(_1339_),
    .B1(_1329_),
    .Y(_0028_));
 sky130_fd_sc_hd__nand3_1 _1708_ (.A(net42),
    .B(_1325_),
    .C(_1336_),
    .Y(_1340_));
 sky130_fd_sc_hd__o31ai_1 _1709_ (.A1(_1279_),
    .A2(_1302_),
    .A3(_1340_),
    .B1(net43),
    .Y(_1341_));
 sky130_fd_sc_hd__or4_1 _1710_ (.A(net43),
    .B(_1278_),
    .C(_1300_),
    .D(_1340_),
    .X(_1342_));
 sky130_fd_sc_hd__a21oi_1 _1711_ (.A1(_1341_),
    .A2(_1342_),
    .B1(_1329_),
    .Y(_0029_));
 sky130_fd_sc_hd__nand4_1 _1712_ (.A(net42),
    .B(net43),
    .C(_1325_),
    .D(_1336_),
    .Y(_1343_));
 sky130_fd_sc_hd__o31ai_1 _1713_ (.A1(_1283_),
    .A2(_1301_),
    .A3(_1343_),
    .B1(net44),
    .Y(_1344_));
 sky130_fd_sc_hd__or4_1 _1714_ (.A(net44),
    .B(_1282_),
    .C(_1300_),
    .D(_1343_),
    .X(_1345_));
 sky130_fd_sc_hd__a21oi_1 _1715_ (.A1(_1344_),
    .A2(_1345_),
    .B1(_1329_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_1 _1716_ (.A(net45),
    .Y(_1346_));
 sky130_fd_sc_hd__nand3b_1 _1717_ (.A_N(\prev_event_inc[4] ),
    .B(net9),
    .C(_1220_),
    .Y(_1347_));
 sky130_fd_sc_hd__xnor2_1 _1718_ (.A(_1346_),
    .B(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__nor2_1 _1719_ (.A(_1218_),
    .B(_1348_),
    .Y(_0031_));
 sky130_fd_sc_hd__clkbuf_4 _1720_ (.A(_1217_),
    .X(_1349_));
 sky130_fd_sc_hd__mux2i_1 _1721_ (.A0(_1549_),
    .A1(net46),
    .S(_1347_),
    .Y(_1350_));
 sky130_fd_sc_hd__nor2_1 _1722_ (.A(_1349_),
    .B(_1350_),
    .Y(_0032_));
 sky130_fd_sc_hd__nand3_4 _1723_ (.A(net269),
    .B(net25),
    .C(net36),
    .Y(_1351_));
 sky130_fd_sc_hd__clkbuf_4 _1724_ (.A(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__o21ai_0 _1725_ (.A1(_1266_),
    .A2(_1352_),
    .B1(net47),
    .Y(_1353_));
 sky130_fd_sc_hd__clkbuf_4 _1726_ (.A(_1265_),
    .X(_1354_));
 sky130_fd_sc_hd__or3_1 _1727_ (.A(net47),
    .B(_1354_),
    .C(_1352_),
    .X(_1355_));
 sky130_fd_sc_hd__a21oi_1 _1728_ (.A1(_1353_),
    .A2(_1355_),
    .B1(_1329_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_1 _1729_ (.A(net48),
    .Y(_1356_));
 sky130_fd_sc_hd__nand4b_1 _1730_ (.A_N(\prev_event_inc[4] ),
    .B(_1548_),
    .C(_1220_),
    .D(net9),
    .Y(_1357_));
 sky130_fd_sc_hd__xnor2_1 _1731_ (.A(_1356_),
    .B(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__nor2_1 _1732_ (.A(_1349_),
    .B(_1358_),
    .Y(_0034_));
 sky130_fd_sc_hd__nand2_1 _1733_ (.A(net45),
    .B(net46),
    .Y(_1359_));
 sky130_fd_sc_hd__nand4b_1 _1734_ (.A_N(\prev_event_inc[4] ),
    .B(net48),
    .C(_1220_),
    .D(net9),
    .Y(_1360_));
 sky130_fd_sc_hd__o21ai_0 _1735_ (.A1(_1359_),
    .A2(_1360_),
    .B1(net49),
    .Y(_1361_));
 sky130_fd_sc_hd__inv_1 _1736_ (.A(net49),
    .Y(_1362_));
 sky130_fd_sc_hd__and2_1 _1737_ (.A(net45),
    .B(net46),
    .X(_1363_));
 sky130_fd_sc_hd__and4b_1 _1738_ (.A_N(\prev_event_inc[4] ),
    .B(net48),
    .C(net4),
    .D(net9),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_4 _1739_ (.A(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__nand3_1 _1740_ (.A(_1362_),
    .B(_1363_),
    .C(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__a21oi_1 _1741_ (.A1(_1361_),
    .A2(_1366_),
    .B1(_1329_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_1 _1742_ (.A(net50),
    .Y(_1367_));
 sky130_fd_sc_hd__nand3_1 _1743_ (.A(net49),
    .B(_1548_),
    .C(_1365_),
    .Y(_1368_));
 sky130_fd_sc_hd__xnor2_1 _1744_ (.A(_1367_),
    .B(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__nor2_1 _1745_ (.A(_1349_),
    .B(_1369_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_1 _1746_ (.A(net51),
    .Y(_1370_));
 sky130_fd_sc_hd__nand4_1 _1747_ (.A(net49),
    .B(net50),
    .C(_1363_),
    .D(_1365_),
    .Y(_1371_));
 sky130_fd_sc_hd__xnor2_1 _1748_ (.A(_1370_),
    .B(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__nor2_1 _1749_ (.A(_1349_),
    .B(_1372_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_1 _1750_ (.A(net52),
    .Y(_1373_));
 sky130_fd_sc_hd__and3_2 _1751_ (.A(net49),
    .B(net50),
    .C(net51),
    .X(_1374_));
 sky130_fd_sc_hd__nand3_1 _1752_ (.A(_1548_),
    .B(_1365_),
    .C(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__xnor2_1 _1753_ (.A(_1373_),
    .B(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__nor2_1 _1754_ (.A(_1349_),
    .B(_1376_),
    .Y(_0038_));
 sky130_fd_sc_hd__nand4_2 _1755_ (.A(net49),
    .B(net50),
    .C(net51),
    .D(net52),
    .Y(_1377_));
 sky130_fd_sc_hd__nor3_1 _1756_ (.A(_1359_),
    .B(_1360_),
    .C(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__xnor2_1 _1757_ (.A(net53),
    .B(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__nor2_1 _1758_ (.A(_1349_),
    .B(_1379_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_1 _1759_ (.A(net54),
    .Y(_1380_));
 sky130_fd_sc_hd__and4_1 _1760_ (.A(net49),
    .B(net50),
    .C(net51),
    .D(net52),
    .X(_1381_));
 sky130_fd_sc_hd__nand4_1 _1761_ (.A(net53),
    .B(_1548_),
    .C(_1365_),
    .D(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__xnor2_1 _1762_ (.A(_1380_),
    .B(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__nor2_1 _1763_ (.A(_1349_),
    .B(_1383_),
    .Y(_0040_));
 sky130_fd_sc_hd__nand2_1 _1764_ (.A(net53),
    .B(net54),
    .Y(_1384_));
 sky130_fd_sc_hd__nor4_1 _1765_ (.A(_1359_),
    .B(_1360_),
    .C(_1377_),
    .D(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__xnor2_1 _1766_ (.A(net55),
    .B(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__nor2_1 _1767_ (.A(_1349_),
    .B(_1386_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_1 _1768_ (.A(net56),
    .Y(_1387_));
 sky130_fd_sc_hd__and3_1 _1769_ (.A(net53),
    .B(net54),
    .C(net55),
    .X(_1388_));
 sky130_fd_sc_hd__nand4_1 _1770_ (.A(_1548_),
    .B(_1365_),
    .C(_1381_),
    .D(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__xnor2_1 _1771_ (.A(_1387_),
    .B(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__nor2_1 _1772_ (.A(_1349_),
    .B(_1390_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_1 _1773_ (.A(net57),
    .Y(_1391_));
 sky130_fd_sc_hd__and4_2 _1774_ (.A(net53),
    .B(net54),
    .C(net55),
    .D(net56),
    .X(_1392_));
 sky130_fd_sc_hd__nand4_4 _1775_ (.A(_1363_),
    .B(_1365_),
    .C(_1381_),
    .D(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__xnor2_1 _1776_ (.A(_1391_),
    .B(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__nor2_1 _1777_ (.A(_1349_),
    .B(_1394_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_1 _1778_ (.A(net47),
    .Y(_1395_));
 sky130_fd_sc_hd__nand4_1 _1779_ (.A(net14),
    .B(net125),
    .C(net247),
    .D(net258),
    .Y(_1396_));
 sky130_fd_sc_hd__or4_1 _1780_ (.A(_1262_),
    .B(_1263_),
    .C(_1351_),
    .D(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__buf_2 _1781_ (.A(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__buf_2 _1782_ (.A(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__o21ai_0 _1783_ (.A1(_1395_),
    .A2(_1399_),
    .B1(net58),
    .Y(_1400_));
 sky130_fd_sc_hd__or3_1 _1784_ (.A(_1395_),
    .B(net58),
    .C(_1399_),
    .X(_1401_));
 sky130_fd_sc_hd__a21oi_1 _1785_ (.A1(_1400_),
    .A2(_1401_),
    .B1(_1329_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand2_2 _1786_ (.A(_1548_),
    .B(_1365_),
    .Y(_1402_));
 sky130_fd_sc_hd__nand2_1 _1787_ (.A(net57),
    .B(_1392_),
    .Y(_1403_));
 sky130_fd_sc_hd__o31ai_1 _1788_ (.A1(_1402_),
    .A2(_1377_),
    .A3(_1403_),
    .B1(net59),
    .Y(_1404_));
 sky130_fd_sc_hd__or4_1 _1789_ (.A(net59),
    .B(_1402_),
    .C(_1377_),
    .D(_1403_),
    .X(_1405_));
 sky130_fd_sc_hd__a21oi_1 _1790_ (.A1(_1404_),
    .A2(_1405_),
    .B1(_1329_),
    .Y(_0045_));
 sky130_fd_sc_hd__nand2_1 _1791_ (.A(net57),
    .B(net59),
    .Y(_1406_));
 sky130_fd_sc_hd__o21ai_0 _1792_ (.A1(_1393_),
    .A2(_1406_),
    .B1(net60),
    .Y(_1407_));
 sky130_fd_sc_hd__or3_1 _1793_ (.A(net60),
    .B(_1393_),
    .C(_1406_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_4 _1794_ (.A(_1287_),
    .X(_1409_));
 sky130_fd_sc_hd__a21oi_1 _1795_ (.A1(_1407_),
    .A2(_1408_),
    .B1(_1409_),
    .Y(_0046_));
 sky130_fd_sc_hd__and4_1 _1796_ (.A(net52),
    .B(net57),
    .C(net59),
    .D(net60),
    .X(_1410_));
 sky130_fd_sc_hd__nand3_2 _1797_ (.A(_1374_),
    .B(_1392_),
    .C(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__o21ai_0 _1798_ (.A1(_1402_),
    .A2(_1411_),
    .B1(net61),
    .Y(_1412_));
 sky130_fd_sc_hd__or3_1 _1799_ (.A(net61),
    .B(_1402_),
    .C(_1411_),
    .X(_1413_));
 sky130_fd_sc_hd__a21oi_1 _1800_ (.A1(_1412_),
    .A2(_1413_),
    .B1(_1409_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_1 _1801_ (.A(net61),
    .Y(_1414_));
 sky130_fd_sc_hd__and3_1 _1802_ (.A(net57),
    .B(net59),
    .C(net60),
    .X(_1415_));
 sky130_fd_sc_hd__inv_1 _1803_ (.A(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__o31ai_1 _1804_ (.A1(_1414_),
    .A2(_1393_),
    .A3(_1416_),
    .B1(net62),
    .Y(_1417_));
 sky130_fd_sc_hd__or4_1 _1805_ (.A(_1414_),
    .B(net62),
    .C(_1393_),
    .D(_1416_),
    .X(_1418_));
 sky130_fd_sc_hd__a21oi_1 _1806_ (.A1(_1417_),
    .A2(_1418_),
    .B1(_1409_),
    .Y(_0048_));
 sky130_fd_sc_hd__nand2_1 _1807_ (.A(net61),
    .B(net62),
    .Y(_1419_));
 sky130_fd_sc_hd__o31ai_1 _1808_ (.A1(_1402_),
    .A2(_1411_),
    .A3(_1419_),
    .B1(net63),
    .Y(_1420_));
 sky130_fd_sc_hd__or4_1 _1809_ (.A(net63),
    .B(_1402_),
    .C(_1411_),
    .D(_1419_),
    .X(_1421_));
 sky130_fd_sc_hd__a21oi_1 _1810_ (.A1(_1420_),
    .A2(_1421_),
    .B1(_1409_),
    .Y(_0049_));
 sky130_fd_sc_hd__nand3_1 _1811_ (.A(net61),
    .B(net62),
    .C(net63),
    .Y(_1422_));
 sky130_fd_sc_hd__o31ai_1 _1812_ (.A1(_1393_),
    .A2(_1416_),
    .A3(_1422_),
    .B1(net64),
    .Y(_1423_));
 sky130_fd_sc_hd__or4_1 _1813_ (.A(net64),
    .B(_1393_),
    .C(_1416_),
    .D(_1422_),
    .X(_1424_));
 sky130_fd_sc_hd__a21oi_1 _1814_ (.A1(_1423_),
    .A2(_1424_),
    .B1(_1409_),
    .Y(_0050_));
 sky130_fd_sc_hd__nand4_1 _1815_ (.A(net61),
    .B(net62),
    .C(net63),
    .D(net64),
    .Y(_1425_));
 sky130_fd_sc_hd__o31ai_1 _1816_ (.A1(_1402_),
    .A2(_1411_),
    .A3(_1425_),
    .B1(net65),
    .Y(_1426_));
 sky130_fd_sc_hd__or4_1 _1817_ (.A(net65),
    .B(_1402_),
    .C(_1411_),
    .D(_1425_),
    .X(_1427_));
 sky130_fd_sc_hd__a21oi_1 _1818_ (.A1(_1426_),
    .A2(_1427_),
    .B1(_1409_),
    .Y(_0051_));
 sky130_fd_sc_hd__and4_1 _1819_ (.A(net61),
    .B(net62),
    .C(net63),
    .D(net64),
    .X(_1428_));
 sky130_fd_sc_hd__nand3_1 _1820_ (.A(net65),
    .B(_1415_),
    .C(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__o21ai_0 _1821_ (.A1(_1393_),
    .A2(_1429_),
    .B1(net66),
    .Y(_1430_));
 sky130_fd_sc_hd__or3_1 _1822_ (.A(net66),
    .B(_1393_),
    .C(_1429_),
    .X(_1431_));
 sky130_fd_sc_hd__a21oi_1 _1823_ (.A1(_1430_),
    .A2(_1431_),
    .B1(_1409_),
    .Y(_0052_));
 sky130_fd_sc_hd__nand4_2 _1824_ (.A(net65),
    .B(_1548_),
    .C(_1365_),
    .D(_1428_),
    .Y(_1432_));
 sky130_fd_sc_hd__clkbuf_2 _1825_ (.A(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__nand4_2 _1826_ (.A(net66),
    .B(_1374_),
    .C(_1392_),
    .D(_1410_),
    .Y(_1434_));
 sky130_fd_sc_hd__o21ai_0 _1827_ (.A1(_1433_),
    .A2(_1434_),
    .B1(net67),
    .Y(_1435_));
 sky130_fd_sc_hd__or3_1 _1828_ (.A(net67),
    .B(_1433_),
    .C(_1434_),
    .X(_1436_));
 sky130_fd_sc_hd__a21oi_1 _1829_ (.A1(_1435_),
    .A2(_1436_),
    .B1(_1409_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_1 _1830_ (.A(net67),
    .Y(_1437_));
 sky130_fd_sc_hd__nand4_1 _1831_ (.A(net65),
    .B(_1363_),
    .C(_1365_),
    .D(_1428_),
    .Y(_1438_));
 sky130_fd_sc_hd__buf_2 _1832_ (.A(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__o31ai_1 _1833_ (.A1(_1437_),
    .A2(_1434_),
    .A3(_1439_),
    .B1(net68),
    .Y(_1440_));
 sky130_fd_sc_hd__or4_1 _1834_ (.A(_1437_),
    .B(net68),
    .C(_1434_),
    .D(_1439_),
    .X(_1441_));
 sky130_fd_sc_hd__a21oi_1 _1835_ (.A1(_1440_),
    .A2(_1441_),
    .B1(_1409_),
    .Y(_0054_));
 sky130_fd_sc_hd__nand2_1 _1836_ (.A(net47),
    .B(net58),
    .Y(_1442_));
 sky130_fd_sc_hd__o31ai_1 _1837_ (.A1(_1266_),
    .A2(_1352_),
    .A3(_1442_),
    .B1(net69),
    .Y(_1443_));
 sky130_fd_sc_hd__or4_1 _1838_ (.A(net69),
    .B(_1354_),
    .C(_1351_),
    .D(_1442_),
    .X(_1444_));
 sky130_fd_sc_hd__a21oi_1 _1839_ (.A1(_1443_),
    .A2(_1444_),
    .B1(_1409_),
    .Y(_0055_));
 sky130_fd_sc_hd__nand2_1 _1840_ (.A(net67),
    .B(net68),
    .Y(_1445_));
 sky130_fd_sc_hd__o31ai_1 _1841_ (.A1(_1433_),
    .A2(_1434_),
    .A3(_1445_),
    .B1(net70),
    .Y(_1446_));
 sky130_fd_sc_hd__or4_1 _1842_ (.A(net70),
    .B(_1433_),
    .C(_1434_),
    .D(_1445_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_4 _1843_ (.A(_1287_),
    .X(_1448_));
 sky130_fd_sc_hd__a21oi_1 _1844_ (.A1(_1446_),
    .A2(_1447_),
    .B1(_1448_),
    .Y(_0056_));
 sky130_fd_sc_hd__and4_1 _1845_ (.A(net66),
    .B(net67),
    .C(net68),
    .D(net70),
    .X(_1449_));
 sky130_fd_sc_hd__nand4_4 _1846_ (.A(_1374_),
    .B(_1392_),
    .C(_1410_),
    .D(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__buf_2 _1847_ (.A(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__o21ai_0 _1848_ (.A1(_1439_),
    .A2(_1451_),
    .B1(net71),
    .Y(_1452_));
 sky130_fd_sc_hd__or3_1 _1849_ (.A(net71),
    .B(_1439_),
    .C(_1451_),
    .X(_1453_));
 sky130_fd_sc_hd__a21oi_1 _1850_ (.A1(_1452_),
    .A2(_1453_),
    .B1(_1448_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_1 _1851_ (.A(net71),
    .Y(_1454_));
 sky130_fd_sc_hd__o31ai_1 _1852_ (.A1(_1454_),
    .A2(_1433_),
    .A3(_1451_),
    .B1(net72),
    .Y(_1455_));
 sky130_fd_sc_hd__or4_1 _1853_ (.A(_1454_),
    .B(net72),
    .C(_1433_),
    .D(_1450_),
    .X(_1456_));
 sky130_fd_sc_hd__a21oi_1 _1854_ (.A1(_1455_),
    .A2(_1456_),
    .B1(_1448_),
    .Y(_0058_));
 sky130_fd_sc_hd__nand2_1 _1855_ (.A(net71),
    .B(net72),
    .Y(_1457_));
 sky130_fd_sc_hd__o31ai_1 _1856_ (.A1(_1439_),
    .A2(_1451_),
    .A3(_1457_),
    .B1(net73),
    .Y(_1458_));
 sky130_fd_sc_hd__or4_1 _1857_ (.A(net73),
    .B(_1439_),
    .C(_1450_),
    .D(_1457_),
    .X(_1459_));
 sky130_fd_sc_hd__a21oi_1 _1858_ (.A1(_1458_),
    .A2(_1459_),
    .B1(_1448_),
    .Y(_0059_));
 sky130_fd_sc_hd__nand3_1 _1859_ (.A(net71),
    .B(net72),
    .C(net73),
    .Y(_1460_));
 sky130_fd_sc_hd__o31ai_1 _1860_ (.A1(_1433_),
    .A2(_1451_),
    .A3(_1460_),
    .B1(net74),
    .Y(_1461_));
 sky130_fd_sc_hd__or4_1 _1861_ (.A(net74),
    .B(_1433_),
    .C(_1450_),
    .D(_1460_),
    .X(_1462_));
 sky130_fd_sc_hd__a21oi_1 _1862_ (.A1(_1461_),
    .A2(_1462_),
    .B1(_1448_),
    .Y(_0060_));
 sky130_fd_sc_hd__nand4_1 _1863_ (.A(net71),
    .B(net72),
    .C(net73),
    .D(net74),
    .Y(_1463_));
 sky130_fd_sc_hd__o31ai_1 _1864_ (.A1(_1439_),
    .A2(_1451_),
    .A3(_1463_),
    .B1(net75),
    .Y(_1464_));
 sky130_fd_sc_hd__or4_1 _1865_ (.A(net75),
    .B(_1439_),
    .C(_1450_),
    .D(_1463_),
    .X(_1465_));
 sky130_fd_sc_hd__a21oi_1 _1866_ (.A1(_1464_),
    .A2(_1465_),
    .B1(_1448_),
    .Y(_0061_));
 sky130_fd_sc_hd__and4_1 _1867_ (.A(net71),
    .B(net72),
    .C(net73),
    .D(net74),
    .X(_1466_));
 sky130_fd_sc_hd__nand2_1 _1868_ (.A(net75),
    .B(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__o31ai_1 _1869_ (.A1(_1433_),
    .A2(_1451_),
    .A3(_1467_),
    .B1(net76),
    .Y(_1468_));
 sky130_fd_sc_hd__or4_1 _1870_ (.A(net76),
    .B(_1432_),
    .C(_1450_),
    .D(_1467_),
    .X(_1469_));
 sky130_fd_sc_hd__a21oi_1 _1871_ (.A1(_1468_),
    .A2(_1469_),
    .B1(_1448_),
    .Y(_0062_));
 sky130_fd_sc_hd__nand3_1 _1872_ (.A(net75),
    .B(net76),
    .C(_1466_),
    .Y(_1470_));
 sky130_fd_sc_hd__o31ai_1 _1873_ (.A1(_1439_),
    .A2(_1451_),
    .A3(_1470_),
    .B1(net77),
    .Y(_1471_));
 sky130_fd_sc_hd__or4_1 _1874_ (.A(net77),
    .B(_1438_),
    .C(_1450_),
    .D(_1470_),
    .X(_1472_));
 sky130_fd_sc_hd__a21oi_1 _1875_ (.A1(_1471_),
    .A2(_1472_),
    .B1(_1448_),
    .Y(_0063_));
 sky130_fd_sc_hd__nand4_1 _1876_ (.A(net75),
    .B(net76),
    .C(net77),
    .D(_1466_),
    .Y(_1473_));
 sky130_fd_sc_hd__o31ai_1 _1877_ (.A1(_1433_),
    .A2(_1451_),
    .A3(_1473_),
    .B1(net78),
    .Y(_1474_));
 sky130_fd_sc_hd__or4_1 _1878_ (.A(net78),
    .B(_1432_),
    .C(_1450_),
    .D(_1473_),
    .X(_1475_));
 sky130_fd_sc_hd__a21oi_1 _1879_ (.A1(_1474_),
    .A2(_1475_),
    .B1(_1448_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_1 _1880_ (.A(net79),
    .Y(_1476_));
 sky130_fd_sc_hd__nor2_1 _1881_ (.A(_1254_),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__buf_4 _1882_ (.A(_1215_),
    .X(_1478_));
 sky130_fd_sc_hd__nor2_1 _1883_ (.A(_1478_),
    .B(net79),
    .Y(_1479_));
 sky130_fd_sc_hd__inv_1 _1884_ (.A(net78),
    .Y(_1480_));
 sky130_fd_sc_hd__nor4_1 _1885_ (.A(_1480_),
    .B(_1439_),
    .C(_1451_),
    .D(_1473_),
    .Y(_1481_));
 sky130_fd_sc_hd__mux2_1 _1886_ (.A0(_1477_),
    .A1(_1479_),
    .S(_1481_),
    .X(_0065_));
 sky130_fd_sc_hd__nand3_1 _1887_ (.A(net47),
    .B(net58),
    .C(net69),
    .Y(_1482_));
 sky130_fd_sc_hd__o21ai_0 _1888_ (.A1(_1399_),
    .A2(_1482_),
    .B1(net80),
    .Y(_1483_));
 sky130_fd_sc_hd__or3_1 _1889_ (.A(net80),
    .B(_1399_),
    .C(_1482_),
    .X(_1484_));
 sky130_fd_sc_hd__a21oi_1 _1890_ (.A1(_1483_),
    .A2(_1484_),
    .B1(_1448_),
    .Y(_0066_));
 sky130_fd_sc_hd__buf_2 _1891_ (.A(_1217_),
    .X(_1485_));
 sky130_fd_sc_hd__and3b_1 _1892_ (.A_N(\prev_event_inc[5] ),
    .B(net10),
    .C(_1220_),
    .X(_1486_));
 sky130_fd_sc_hd__xnor2_1 _1893_ (.A(net81),
    .B(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__nor2_1 _1894_ (.A(_1485_),
    .B(_1487_),
    .Y(_0067_));
 sky130_fd_sc_hd__mux2i_1 _1895_ (.A0(net82),
    .A1(_1547_),
    .S(_1486_),
    .Y(_1488_));
 sky130_fd_sc_hd__nor2_1 _1896_ (.A(_1485_),
    .B(_1488_),
    .Y(_0068_));
 sky130_fd_sc_hd__clkbuf_4 _1897_ (.A(_1546_),
    .X(_1489_));
 sky130_fd_sc_hd__nand2_1 _1898_ (.A(_1489_),
    .B(_1486_),
    .Y(_1490_));
 sky130_fd_sc_hd__xor2_1 _1899_ (.A(net83),
    .B(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__nor2_1 _1900_ (.A(_1485_),
    .B(_1491_),
    .Y(_0069_));
 sky130_fd_sc_hd__nand4b_4 _1901_ (.A_N(\prev_event_inc[5] ),
    .B(net83),
    .C(net4),
    .D(net10),
    .Y(_1492_));
 sky130_fd_sc_hd__nand2_2 _1902_ (.A(net81),
    .B(net82),
    .Y(_1493_));
 sky130_fd_sc_hd__o21ai_0 _1903_ (.A1(_1492_),
    .A2(_1493_),
    .B1(net84),
    .Y(_1494_));
 sky130_fd_sc_hd__or3_1 _1904_ (.A(net84),
    .B(_1492_),
    .C(_1493_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_4 _1905_ (.A(_1287_),
    .X(_1496_));
 sky130_fd_sc_hd__a21oi_1 _1906_ (.A1(_1494_),
    .A2(_1495_),
    .B1(_1496_),
    .Y(_0070_));
 sky130_fd_sc_hd__and4b_1 _1907_ (.A_N(\prev_event_inc[5] ),
    .B(net83),
    .C(_1219_),
    .D(net10),
    .X(_1497_));
 sky130_fd_sc_hd__buf_2 _1908_ (.A(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__nand3_1 _1909_ (.A(net84),
    .B(_1489_),
    .C(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__xor2_1 _1910_ (.A(net85),
    .B(_1499_),
    .X(_1500_));
 sky130_fd_sc_hd__nor2_1 _1911_ (.A(_1485_),
    .B(_1500_),
    .Y(_0071_));
 sky130_fd_sc_hd__nand2_1 _1912_ (.A(net84),
    .B(net85),
    .Y(_1501_));
 sky130_fd_sc_hd__nor3_1 _1913_ (.A(_1492_),
    .B(_1493_),
    .C(_1501_),
    .Y(_1502_));
 sky130_fd_sc_hd__xnor2_1 _1914_ (.A(net86),
    .B(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__nor2_1 _1915_ (.A(_1485_),
    .B(_1503_),
    .Y(_0072_));
 sky130_fd_sc_hd__and3_1 _1916_ (.A(net84),
    .B(net85),
    .C(net86),
    .X(_1504_));
 sky130_fd_sc_hd__nand3_1 _1917_ (.A(_1489_),
    .B(_1498_),
    .C(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__xor2_1 _1918_ (.A(net87),
    .B(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__nor2_1 _1919_ (.A(_1485_),
    .B(_1506_),
    .Y(_0073_));
 sky130_fd_sc_hd__nand4_2 _1920_ (.A(net84),
    .B(net85),
    .C(net86),
    .D(net87),
    .Y(_1507_));
 sky130_fd_sc_hd__nor3_1 _1921_ (.A(_1492_),
    .B(_1493_),
    .C(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__xnor2_1 _1922_ (.A(net88),
    .B(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__nor2_1 _1923_ (.A(_1485_),
    .B(_1509_),
    .Y(_0074_));
 sky130_fd_sc_hd__and4_1 _1924_ (.A(net84),
    .B(net85),
    .C(net86),
    .D(net87),
    .X(_1510_));
 sky130_fd_sc_hd__nand4_1 _1925_ (.A(net88),
    .B(_1489_),
    .C(_1498_),
    .D(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__xor2_1 _1926_ (.A(net89),
    .B(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__nor2_1 _1927_ (.A(_1485_),
    .B(_1512_),
    .Y(_0075_));
 sky130_fd_sc_hd__nand2_1 _1928_ (.A(net88),
    .B(net89),
    .Y(_1513_));
 sky130_fd_sc_hd__nor4_1 _1929_ (.A(_1492_),
    .B(_1493_),
    .C(_1507_),
    .D(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__xnor2_1 _1930_ (.A(net90),
    .B(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__nor2_1 _1931_ (.A(_1485_),
    .B(_1515_),
    .Y(_0076_));
 sky130_fd_sc_hd__nand4_1 _1932_ (.A(net47),
    .B(net58),
    .C(net69),
    .D(net80),
    .Y(_1516_));
 sky130_fd_sc_hd__o31ai_1 _1933_ (.A1(_1266_),
    .A2(_1352_),
    .A3(_1516_),
    .B1(net91),
    .Y(_1517_));
 sky130_fd_sc_hd__or4_1 _1934_ (.A(net91),
    .B(_1354_),
    .C(_1351_),
    .D(_1516_),
    .X(_1518_));
 sky130_fd_sc_hd__a21oi_1 _1935_ (.A1(_1517_),
    .A2(_1518_),
    .B1(_1496_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_1 _1936_ (.A(_1489_),
    .Y(_1519_));
 sky130_fd_sc_hd__nand3_1 _1937_ (.A(net88),
    .B(net89),
    .C(net90),
    .Y(_1520_));
 sky130_fd_sc_hd__nor4_1 _1938_ (.A(_1519_),
    .B(_1492_),
    .C(_1507_),
    .D(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__xnor2_1 _1939_ (.A(net92),
    .B(_1521_),
    .Y(_1522_));
 sky130_fd_sc_hd__nor2_1 _1940_ (.A(_1485_),
    .B(_1522_),
    .Y(_0078_));
 sky130_fd_sc_hd__buf_4 _1941_ (.A(_1217_),
    .X(_1523_));
 sky130_fd_sc_hd__and4_2 _1942_ (.A(net88),
    .B(net89),
    .C(net90),
    .D(net92),
    .X(_1524_));
 sky130_fd_sc_hd__or4b_1 _1943_ (.A(_1492_),
    .B(_1493_),
    .C(_1507_),
    .D_N(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__clkbuf_2 _1944_ (.A(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__xor2_1 _1945_ (.A(net93),
    .B(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__nor2_1 _1946_ (.A(_1523_),
    .B(_1527_),
    .Y(_0079_));
 sky130_fd_sc_hd__nand3_1 _1947_ (.A(_1489_),
    .B(_1498_),
    .C(_1510_),
    .Y(_1528_));
 sky130_fd_sc_hd__nand2_1 _1948_ (.A(net93),
    .B(_1524_),
    .Y(_1529_));
 sky130_fd_sc_hd__o21ai_0 _1949_ (.A1(_1528_),
    .A2(_1529_),
    .B1(net94),
    .Y(_1530_));
 sky130_fd_sc_hd__or3_1 _1950_ (.A(net94),
    .B(_1528_),
    .C(_1529_),
    .X(_1531_));
 sky130_fd_sc_hd__a21oi_1 _1951_ (.A1(_1530_),
    .A2(_1531_),
    .B1(_1496_),
    .Y(_0080_));
 sky130_fd_sc_hd__nand2_1 _1952_ (.A(net93),
    .B(net94),
    .Y(_1532_));
 sky130_fd_sc_hd__o21ai_0 _1953_ (.A1(_1526_),
    .A2(_1532_),
    .B1(net95),
    .Y(_1533_));
 sky130_fd_sc_hd__or3_1 _1954_ (.A(net95),
    .B(_1526_),
    .C(_1532_),
    .X(_1534_));
 sky130_fd_sc_hd__a21oi_1 _1955_ (.A1(_1533_),
    .A2(_1534_),
    .B1(_1496_),
    .Y(_0081_));
 sky130_fd_sc_hd__nand2_1 _1956_ (.A(_1489_),
    .B(_1498_),
    .Y(_1535_));
 sky130_fd_sc_hd__and3_2 _1957_ (.A(net93),
    .B(net94),
    .C(net95),
    .X(_1536_));
 sky130_fd_sc_hd__nand4_2 _1958_ (.A(net87),
    .B(_1504_),
    .C(_1524_),
    .D(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__o21ai_0 _1959_ (.A1(_1535_),
    .A2(_1537_),
    .B1(net96),
    .Y(_0264_));
 sky130_fd_sc_hd__or3_1 _1960_ (.A(net96),
    .B(_1535_),
    .C(_1537_),
    .X(_0265_));
 sky130_fd_sc_hd__a21oi_1 _1961_ (.A1(_0264_),
    .A2(_0265_),
    .B1(_1496_),
    .Y(_0082_));
 sky130_fd_sc_hd__nand2_1 _1962_ (.A(net96),
    .B(_1536_),
    .Y(_0266_));
 sky130_fd_sc_hd__o21ai_0 _1963_ (.A1(_1526_),
    .A2(_0266_),
    .B1(net97),
    .Y(_0267_));
 sky130_fd_sc_hd__or3_1 _1964_ (.A(net97),
    .B(_1526_),
    .C(_0266_),
    .X(_0268_));
 sky130_fd_sc_hd__a21oi_1 _1965_ (.A1(_0267_),
    .A2(_0268_),
    .B1(_1496_),
    .Y(_0083_));
 sky130_fd_sc_hd__nand2_1 _1966_ (.A(net96),
    .B(net97),
    .Y(_0269_));
 sky130_fd_sc_hd__o31ai_1 _1967_ (.A1(_1535_),
    .A2(_1537_),
    .A3(_0269_),
    .B1(net98),
    .Y(_0270_));
 sky130_fd_sc_hd__or4_1 _1968_ (.A(net98),
    .B(_1535_),
    .C(_1537_),
    .D(_0269_),
    .X(_0271_));
 sky130_fd_sc_hd__a21oi_1 _1969_ (.A1(_0270_),
    .A2(_0271_),
    .B1(_1496_),
    .Y(_0084_));
 sky130_fd_sc_hd__nand4_1 _1970_ (.A(net96),
    .B(net97),
    .C(net98),
    .D(_1536_),
    .Y(_0272_));
 sky130_fd_sc_hd__o21ai_0 _1971_ (.A1(_1526_),
    .A2(_0272_),
    .B1(net99),
    .Y(_0273_));
 sky130_fd_sc_hd__or3_1 _1972_ (.A(net99),
    .B(_1526_),
    .C(_0272_),
    .X(_0274_));
 sky130_fd_sc_hd__a21oi_1 _1973_ (.A1(_0273_),
    .A2(_0274_),
    .B1(_1496_),
    .Y(_0085_));
 sky130_fd_sc_hd__nand4_1 _1974_ (.A(net96),
    .B(net97),
    .C(net98),
    .D(net99),
    .Y(_0275_));
 sky130_fd_sc_hd__o31ai_1 _1975_ (.A1(_1535_),
    .A2(_1537_),
    .A3(_0275_),
    .B1(net100),
    .Y(_0276_));
 sky130_fd_sc_hd__or4_1 _1976_ (.A(net100),
    .B(_1535_),
    .C(_1537_),
    .D(_0275_),
    .X(_0277_));
 sky130_fd_sc_hd__a21oi_1 _1977_ (.A1(_0276_),
    .A2(_0277_),
    .B1(_1496_),
    .Y(_0086_));
 sky130_fd_sc_hd__and4_1 _1978_ (.A(net96),
    .B(net97),
    .C(net98),
    .D(net99),
    .X(_0278_));
 sky130_fd_sc_hd__nand3_1 _1979_ (.A(net100),
    .B(_1536_),
    .C(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__o21ai_0 _1980_ (.A1(_1526_),
    .A2(_0279_),
    .B1(net101),
    .Y(_0280_));
 sky130_fd_sc_hd__or3_1 _1981_ (.A(net101),
    .B(_1526_),
    .C(_0279_),
    .X(_0281_));
 sky130_fd_sc_hd__a21oi_1 _1982_ (.A1(_0280_),
    .A2(_0281_),
    .B1(_1496_),
    .Y(_0087_));
 sky130_fd_sc_hd__and4_1 _1983_ (.A(net47),
    .B(net58),
    .C(net69),
    .D(net80),
    .X(_0282_));
 sky130_fd_sc_hd__buf_2 _1984_ (.A(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_1 _1985_ (.A(net91),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_0 _1986_ (.A1(_1399_),
    .A2(_0284_),
    .B1(net102),
    .Y(_0285_));
 sky130_fd_sc_hd__or3_1 _1987_ (.A(net102),
    .B(_1398_),
    .C(_0284_),
    .X(_0286_));
 sky130_fd_sc_hd__buf_2 _1988_ (.A(_1287_),
    .X(_0287_));
 sky130_fd_sc_hd__a21oi_1 _1989_ (.A1(_0285_),
    .A2(_0286_),
    .B1(_0287_),
    .Y(_0088_));
 sky130_fd_sc_hd__and2_0 _1990_ (.A(net87),
    .B(net101),
    .X(_0288_));
 sky130_fd_sc_hd__nand4_4 _1991_ (.A(_1504_),
    .B(_1524_),
    .C(_1536_),
    .D(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__buf_2 _1992_ (.A(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__buf_2 _1993_ (.A(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__nand3_2 _1994_ (.A(net100),
    .B(_1498_),
    .C(_0278_),
    .Y(_0292_));
 sky130_fd_sc_hd__o31ai_1 _1995_ (.A1(_1519_),
    .A2(_0291_),
    .A3(_0292_),
    .B1(net103),
    .Y(_0293_));
 sky130_fd_sc_hd__or4_1 _1996_ (.A(net103),
    .B(_1519_),
    .C(_0290_),
    .D(_0292_),
    .X(_0294_));
 sky130_fd_sc_hd__a21oi_1 _1997_ (.A1(_0293_),
    .A2(_0294_),
    .B1(_0287_),
    .Y(_0089_));
 sky130_fd_sc_hd__nand3_1 _1998_ (.A(net81),
    .B(net82),
    .C(net103),
    .Y(_0295_));
 sky130_fd_sc_hd__o31ai_1 _1999_ (.A1(_0291_),
    .A2(_0292_),
    .A3(_0295_),
    .B1(net104),
    .Y(_0296_));
 sky130_fd_sc_hd__or4_1 _2000_ (.A(net104),
    .B(_0290_),
    .C(_0292_),
    .D(_0295_),
    .X(_0297_));
 sky130_fd_sc_hd__a21oi_1 _2001_ (.A1(_0296_),
    .A2(_0297_),
    .B1(_0287_),
    .Y(_0090_));
 sky130_fd_sc_hd__nand3_1 _2002_ (.A(net103),
    .B(net104),
    .C(_1489_),
    .Y(_0298_));
 sky130_fd_sc_hd__o31ai_1 _2003_ (.A1(_0291_),
    .A2(_0292_),
    .A3(_0298_),
    .B1(net105),
    .Y(_0299_));
 sky130_fd_sc_hd__or4_1 _2004_ (.A(net105),
    .B(_0290_),
    .C(_0292_),
    .D(_0298_),
    .X(_0300_));
 sky130_fd_sc_hd__a21oi_1 _2005_ (.A1(_0299_),
    .A2(_0300_),
    .B1(_0287_),
    .Y(_0091_));
 sky130_fd_sc_hd__and4_1 _2006_ (.A(net100),
    .B(net103),
    .C(net104),
    .D(net105),
    .X(_0301_));
 sky130_fd_sc_hd__or4b_1 _2007_ (.A(_1492_),
    .B(_1493_),
    .C(_0275_),
    .D_N(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_2 _2008_ (.A(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__o21ai_0 _2009_ (.A1(_0291_),
    .A2(_0303_),
    .B1(net106),
    .Y(_0304_));
 sky130_fd_sc_hd__or3_1 _2010_ (.A(net106),
    .B(_0290_),
    .C(_0303_),
    .X(_0305_));
 sky130_fd_sc_hd__a21oi_1 _2011_ (.A1(_0304_),
    .A2(_0305_),
    .B1(_0287_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_1 _2012_ (.A(net106),
    .Y(_0306_));
 sky130_fd_sc_hd__nand4_4 _2013_ (.A(_1489_),
    .B(_1498_),
    .C(_0278_),
    .D(_0301_),
    .Y(_0307_));
 sky130_fd_sc_hd__o31ai_1 _2014_ (.A1(_0306_),
    .A2(_0291_),
    .A3(_0307_),
    .B1(net107),
    .Y(_0308_));
 sky130_fd_sc_hd__or4_1 _2015_ (.A(_0306_),
    .B(net107),
    .C(_0290_),
    .D(_0307_),
    .X(_0309_));
 sky130_fd_sc_hd__a21oi_1 _2016_ (.A1(_0308_),
    .A2(_0309_),
    .B1(_0287_),
    .Y(_0093_));
 sky130_fd_sc_hd__nand2_1 _2017_ (.A(net106),
    .B(net107),
    .Y(_0310_));
 sky130_fd_sc_hd__o31ai_1 _2018_ (.A1(_0291_),
    .A2(_0303_),
    .A3(_0310_),
    .B1(net108),
    .Y(_0311_));
 sky130_fd_sc_hd__or4_1 _2019_ (.A(net108),
    .B(_0290_),
    .C(_0303_),
    .D(_0310_),
    .X(_0312_));
 sky130_fd_sc_hd__a21oi_1 _2020_ (.A1(_0311_),
    .A2(_0312_),
    .B1(_0287_),
    .Y(_0094_));
 sky130_fd_sc_hd__nand3_1 _2021_ (.A(net106),
    .B(net107),
    .C(net108),
    .Y(_0313_));
 sky130_fd_sc_hd__o31ai_1 _2022_ (.A1(_0291_),
    .A2(_0307_),
    .A3(_0313_),
    .B1(net109),
    .Y(_0314_));
 sky130_fd_sc_hd__or4_1 _2023_ (.A(net109),
    .B(_0290_),
    .C(_0307_),
    .D(_0313_),
    .X(_0315_));
 sky130_fd_sc_hd__a21oi_1 _2024_ (.A1(_0314_),
    .A2(_0315_),
    .B1(_0287_),
    .Y(_0095_));
 sky130_fd_sc_hd__nand4_1 _2025_ (.A(net106),
    .B(net107),
    .C(net108),
    .D(net109),
    .Y(_0316_));
 sky130_fd_sc_hd__o31ai_1 _2026_ (.A1(_0291_),
    .A2(_0303_),
    .A3(_0316_),
    .B1(net110),
    .Y(_0317_));
 sky130_fd_sc_hd__or4_1 _2027_ (.A(net110),
    .B(_0289_),
    .C(_0303_),
    .D(_0316_),
    .X(_0318_));
 sky130_fd_sc_hd__a21oi_1 _2028_ (.A1(_0317_),
    .A2(_0318_),
    .B1(_0287_),
    .Y(_0096_));
 sky130_fd_sc_hd__and4_1 _2029_ (.A(net106),
    .B(net107),
    .C(net108),
    .D(net109),
    .X(_0319_));
 sky130_fd_sc_hd__nand2_1 _2030_ (.A(net110),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__o31ai_1 _2031_ (.A1(_0291_),
    .A2(_0307_),
    .A3(_0320_),
    .B1(net111),
    .Y(_0321_));
 sky130_fd_sc_hd__or4_1 _2032_ (.A(net111),
    .B(_0289_),
    .C(_0307_),
    .D(_0320_),
    .X(_0322_));
 sky130_fd_sc_hd__a21oi_1 _2033_ (.A1(_0321_),
    .A2(_0322_),
    .B1(_0287_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand3_1 _2034_ (.A(net110),
    .B(net111),
    .C(_0319_),
    .Y(_0323_));
 sky130_fd_sc_hd__o31ai_1 _2035_ (.A1(_0291_),
    .A2(_0303_),
    .A3(_0323_),
    .B1(net112),
    .Y(_0324_));
 sky130_fd_sc_hd__or4_1 _2036_ (.A(net112),
    .B(_0289_),
    .C(_0303_),
    .D(_0323_),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_4 _2037_ (.A(_1287_),
    .X(_0326_));
 sky130_fd_sc_hd__a21oi_1 _2038_ (.A1(_0324_),
    .A2(_0325_),
    .B1(_0326_),
    .Y(_0098_));
 sky130_fd_sc_hd__nand3_1 _2039_ (.A(net91),
    .B(net102),
    .C(_0283_),
    .Y(_0327_));
 sky130_fd_sc_hd__o31ai_1 _2040_ (.A1(_1266_),
    .A2(_1352_),
    .A3(_0327_),
    .B1(net113),
    .Y(_0328_));
 sky130_fd_sc_hd__or4_1 _2041_ (.A(net113),
    .B(_1354_),
    .C(_1351_),
    .D(_0327_),
    .X(_0329_));
 sky130_fd_sc_hd__a21oi_1 _2042_ (.A1(_0328_),
    .A2(_0329_),
    .B1(_0326_),
    .Y(_0099_));
 sky130_fd_sc_hd__and3_1 _2043_ (.A(net110),
    .B(net111),
    .C(net112),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _2044_ (.A(_0319_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__o31ai_1 _2045_ (.A1(_0290_),
    .A2(_0307_),
    .A3(_0331_),
    .B1(net114),
    .Y(_0332_));
 sky130_fd_sc_hd__or4_1 _2046_ (.A(net114),
    .B(_0289_),
    .C(_0307_),
    .D(_0331_),
    .X(_0333_));
 sky130_fd_sc_hd__a21oi_1 _2047_ (.A1(_0332_),
    .A2(_0333_),
    .B1(_0326_),
    .Y(_0100_));
 sky130_fd_sc_hd__nand3_1 _2048_ (.A(net114),
    .B(_0319_),
    .C(_0330_),
    .Y(_0334_));
 sky130_fd_sc_hd__o31ai_1 _2049_ (.A1(_0290_),
    .A2(_0303_),
    .A3(_0334_),
    .B1(net115),
    .Y(_0335_));
 sky130_fd_sc_hd__or4_1 _2050_ (.A(net115),
    .B(_0289_),
    .C(_0303_),
    .D(_0334_),
    .X(_0336_));
 sky130_fd_sc_hd__a21oi_1 _2051_ (.A1(_0335_),
    .A2(_0336_),
    .B1(_0326_),
    .Y(_0101_));
 sky130_fd_sc_hd__nand3b_1 _2052_ (.A_N(\prev_event_inc[6] ),
    .B(net11),
    .C(_1220_),
    .Y(_0337_));
 sky130_fd_sc_hd__xor2_1 _2053_ (.A(net116),
    .B(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__nor2_1 _2054_ (.A(_1523_),
    .B(_0338_),
    .Y(_0102_));
 sky130_fd_sc_hd__mux2i_1 _2055_ (.A0(_1545_),
    .A1(net117),
    .S(_0337_),
    .Y(_0339_));
 sky130_fd_sc_hd__nor2_1 _2056_ (.A(_1523_),
    .B(_0339_),
    .Y(_0103_));
 sky130_fd_sc_hd__nand4b_1 _2057_ (.A_N(\prev_event_inc[6] ),
    .B(_1544_),
    .C(_1220_),
    .D(net11),
    .Y(_0340_));
 sky130_fd_sc_hd__xor2_1 _2058_ (.A(net118),
    .B(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_1 _2059_ (.A(_1523_),
    .B(_0341_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _2060_ (.A(net116),
    .B(net117),
    .Y(_0342_));
 sky130_fd_sc_hd__nand4b_1 _2061_ (.A_N(\prev_event_inc[6] ),
    .B(net118),
    .C(_1219_),
    .D(net11),
    .Y(_0343_));
 sky130_fd_sc_hd__o21ai_0 _2062_ (.A1(_0342_),
    .A2(_0343_),
    .B1(net119),
    .Y(_0344_));
 sky130_fd_sc_hd__or3_1 _2063_ (.A(net119),
    .B(_0342_),
    .C(_0343_),
    .X(_0345_));
 sky130_fd_sc_hd__a21oi_1 _2064_ (.A1(_0344_),
    .A2(_0345_),
    .B1(_0326_),
    .Y(_0105_));
 sky130_fd_sc_hd__and4b_1 _2065_ (.A_N(\prev_event_inc[6] ),
    .B(net118),
    .C(net4),
    .D(net11),
    .X(_0346_));
 sky130_fd_sc_hd__buf_2 _2066_ (.A(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__nand3_1 _2067_ (.A(net119),
    .B(_1544_),
    .C(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__xor2_1 _2068_ (.A(net120),
    .B(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__nor2_1 _2069_ (.A(_1523_),
    .B(_0349_),
    .Y(_0106_));
 sky130_fd_sc_hd__and2_1 _2070_ (.A(net116),
    .B(net117),
    .X(_0350_));
 sky130_fd_sc_hd__nand4_1 _2071_ (.A(net119),
    .B(net120),
    .C(_0350_),
    .D(_0347_),
    .Y(_0351_));
 sky130_fd_sc_hd__xor2_1 _2072_ (.A(net121),
    .B(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(_1523_),
    .B(_0352_),
    .Y(_0107_));
 sky130_fd_sc_hd__and3_2 _2074_ (.A(net119),
    .B(net120),
    .C(net121),
    .X(_0353_));
 sky130_fd_sc_hd__nand3_2 _2075_ (.A(_1544_),
    .B(_0347_),
    .C(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__xor2_1 _2076_ (.A(net122),
    .B(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__nor2_1 _2077_ (.A(_1523_),
    .B(_0355_),
    .Y(_0108_));
 sky130_fd_sc_hd__nand4_1 _2078_ (.A(net119),
    .B(net120),
    .C(net121),
    .D(net122),
    .Y(_0356_));
 sky130_fd_sc_hd__nor3_1 _2079_ (.A(_0342_),
    .B(_0343_),
    .C(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__xnor2_1 _2080_ (.A(net123),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nor2_1 _2081_ (.A(_1523_),
    .B(_0358_),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_1 _2082_ (.A(net113),
    .Y(_0359_));
 sky130_fd_sc_hd__o31ai_1 _2083_ (.A1(_0359_),
    .A2(_1399_),
    .A3(_0327_),
    .B1(net124),
    .Y(_0360_));
 sky130_fd_sc_hd__or4_1 _2084_ (.A(_0359_),
    .B(net124),
    .C(_1398_),
    .D(_0327_),
    .X(_0361_));
 sky130_fd_sc_hd__a21oi_1 _2085_ (.A1(_0360_),
    .A2(_0361_),
    .B1(_0326_),
    .Y(_0110_));
 sky130_fd_sc_hd__mux2i_1 _2086_ (.A0(net125),
    .A1(_1541_),
    .S(_1221_),
    .Y(_0362_));
 sky130_fd_sc_hd__nor2_1 _2087_ (.A(_1523_),
    .B(_0362_),
    .Y(_0111_));
 sky130_fd_sc_hd__and4_2 _2088_ (.A(net119),
    .B(net120),
    .C(net121),
    .D(net122),
    .X(_0363_));
 sky130_fd_sc_hd__nand4_1 _2089_ (.A(net123),
    .B(_1544_),
    .C(_0347_),
    .D(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__xor2_1 _2090_ (.A(net126),
    .B(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__nor2_1 _2091_ (.A(_1523_),
    .B(_0365_),
    .Y(_0112_));
 sky130_fd_sc_hd__clkbuf_4 _2092_ (.A(_1217_),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _2093_ (.A(net123),
    .B(net126),
    .Y(_0367_));
 sky130_fd_sc_hd__nor4_1 _2094_ (.A(_0342_),
    .B(_0343_),
    .C(_0356_),
    .D(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__xnor2_1 _2095_ (.A(net127),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _2096_ (.A(_0366_),
    .B(_0369_),
    .Y(_0113_));
 sky130_fd_sc_hd__and3_1 _2097_ (.A(net123),
    .B(net126),
    .C(net127),
    .X(_0370_));
 sky130_fd_sc_hd__nand4_1 _2098_ (.A(_1544_),
    .B(_0347_),
    .C(_0363_),
    .D(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__xor2_1 _2099_ (.A(net128),
    .B(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__nor2_1 _2100_ (.A(_0366_),
    .B(_0372_),
    .Y(_0114_));
 sky130_fd_sc_hd__and4_2 _2101_ (.A(net123),
    .B(net126),
    .C(net127),
    .D(net128),
    .X(_0373_));
 sky130_fd_sc_hd__nand4_4 _2102_ (.A(_0350_),
    .B(_0347_),
    .C(_0363_),
    .D(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__xor2_1 _2103_ (.A(net129),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__nor2_1 _2104_ (.A(_0366_),
    .B(_0375_),
    .Y(_0115_));
 sky130_fd_sc_hd__nand3_1 _2105_ (.A(_1544_),
    .B(_0347_),
    .C(_0363_),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2_1 _2106_ (.A(net129),
    .B(_0373_),
    .Y(_0377_));
 sky130_fd_sc_hd__o21ai_0 _2107_ (.A1(_0376_),
    .A2(_0377_),
    .B1(net130),
    .Y(_0378_));
 sky130_fd_sc_hd__or3_1 _2108_ (.A(net130),
    .B(_0376_),
    .C(_0377_),
    .X(_0379_));
 sky130_fd_sc_hd__a21oi_1 _2109_ (.A1(_0378_),
    .A2(_0379_),
    .B1(_0326_),
    .Y(_0116_));
 sky130_fd_sc_hd__nand2_1 _2110_ (.A(net129),
    .B(net130),
    .Y(_0380_));
 sky130_fd_sc_hd__o21ai_0 _2111_ (.A1(_0374_),
    .A2(_0380_),
    .B1(net131),
    .Y(_0381_));
 sky130_fd_sc_hd__or3_1 _2112_ (.A(net131),
    .B(_0374_),
    .C(_0380_),
    .X(_0382_));
 sky130_fd_sc_hd__a21oi_1 _2113_ (.A1(_0381_),
    .A2(_0382_),
    .B1(_0326_),
    .Y(_0117_));
 sky130_fd_sc_hd__and4_1 _2114_ (.A(net122),
    .B(net129),
    .C(net130),
    .D(net131),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _2115_ (.A(_0373_),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__o21ai_0 _2116_ (.A1(_0354_),
    .A2(_0384_),
    .B1(net132),
    .Y(_0385_));
 sky130_fd_sc_hd__or3_1 _2117_ (.A(net132),
    .B(_0354_),
    .C(_0384_),
    .X(_0386_));
 sky130_fd_sc_hd__a21oi_1 _2118_ (.A1(_0385_),
    .A2(_0386_),
    .B1(_0326_),
    .Y(_0118_));
 sky130_fd_sc_hd__and3_1 _2119_ (.A(net129),
    .B(net130),
    .C(net131),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _2120_ (.A(net132),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__o21ai_0 _2121_ (.A1(_0374_),
    .A2(_0388_),
    .B1(net133),
    .Y(_0389_));
 sky130_fd_sc_hd__or3_1 _2122_ (.A(net133),
    .B(_0374_),
    .C(_0388_),
    .X(_0390_));
 sky130_fd_sc_hd__a21oi_1 _2123_ (.A1(_0389_),
    .A2(_0390_),
    .B1(_0326_),
    .Y(_0119_));
 sky130_fd_sc_hd__nand2_1 _2124_ (.A(net132),
    .B(net133),
    .Y(_0391_));
 sky130_fd_sc_hd__o31ai_1 _2125_ (.A1(_0354_),
    .A2(_0384_),
    .A3(_0391_),
    .B1(net134),
    .Y(_0392_));
 sky130_fd_sc_hd__or4_1 _2126_ (.A(net134),
    .B(_0354_),
    .C(_0384_),
    .D(_0391_),
    .X(_0393_));
 sky130_fd_sc_hd__buf_4 _2127_ (.A(_1254_),
    .X(_0394_));
 sky130_fd_sc_hd__a21oi_1 _2128_ (.A1(_0392_),
    .A2(_0393_),
    .B1(_0394_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand4_1 _2129_ (.A(net132),
    .B(net133),
    .C(net134),
    .D(_0387_),
    .Y(_0395_));
 sky130_fd_sc_hd__o21ai_0 _2130_ (.A1(_0374_),
    .A2(_0395_),
    .B1(net135),
    .Y(_0396_));
 sky130_fd_sc_hd__or3_1 _2131_ (.A(net135),
    .B(_0374_),
    .C(_0395_),
    .X(_0397_));
 sky130_fd_sc_hd__a21oi_1 _2132_ (.A1(_0396_),
    .A2(_0397_),
    .B1(_0394_),
    .Y(_0121_));
 sky130_fd_sc_hd__and4_1 _2133_ (.A(net91),
    .B(net102),
    .C(net113),
    .D(net124),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _2134_ (.A(_0283_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__o31ai_1 _2135_ (.A1(_1266_),
    .A2(_1352_),
    .A3(_0399_),
    .B1(net136),
    .Y(_0400_));
 sky130_fd_sc_hd__or4_1 _2136_ (.A(net136),
    .B(_1354_),
    .C(_1351_),
    .D(_0399_),
    .X(_0401_));
 sky130_fd_sc_hd__a21oi_1 _2137_ (.A1(_0400_),
    .A2(_0401_),
    .B1(_0394_),
    .Y(_0122_));
 sky130_fd_sc_hd__nor2b_1 _2138_ (.A(_1216_),
    .B_N(net137),
    .Y(_0402_));
 sky130_fd_sc_hd__nor2_1 _2139_ (.A(_1478_),
    .B(net137),
    .Y(_0403_));
 sky130_fd_sc_hd__and4_1 _2140_ (.A(net132),
    .B(net133),
    .C(net134),
    .D(net135),
    .X(_0404_));
 sky130_fd_sc_hd__nor3b_1 _2141_ (.A(_0354_),
    .B(_0384_),
    .C_N(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__mux2_1 _2142_ (.A0(_0402_),
    .A1(_0403_),
    .S(_0405_),
    .X(_0123_));
 sky130_fd_sc_hd__nand3_1 _2143_ (.A(net137),
    .B(_0387_),
    .C(_0404_),
    .Y(_0406_));
 sky130_fd_sc_hd__o21ai_0 _2144_ (.A1(_0374_),
    .A2(_0406_),
    .B1(net138),
    .Y(_0407_));
 sky130_fd_sc_hd__or3_1 _2145_ (.A(net138),
    .B(_0374_),
    .C(_0406_),
    .X(_0408_));
 sky130_fd_sc_hd__a21oi_1 _2146_ (.A1(_0407_),
    .A2(_0408_),
    .B1(_0394_),
    .Y(_0124_));
 sky130_fd_sc_hd__nand4_2 _2147_ (.A(net138),
    .B(_0353_),
    .C(_0373_),
    .D(_0383_),
    .Y(_0409_));
 sky130_fd_sc_hd__nand4_1 _2148_ (.A(net137),
    .B(_1544_),
    .C(_0347_),
    .D(_0404_),
    .Y(_0410_));
 sky130_fd_sc_hd__buf_2 _2149_ (.A(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__o21ai_0 _2150_ (.A1(_0409_),
    .A2(_0411_),
    .B1(net139),
    .Y(_0412_));
 sky130_fd_sc_hd__or3_1 _2151_ (.A(net139),
    .B(_0409_),
    .C(_0411_),
    .X(_0413_));
 sky130_fd_sc_hd__a21oi_1 _2152_ (.A1(_0412_),
    .A2(_0413_),
    .B1(_0394_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_1 _2153_ (.A(net139),
    .Y(_0414_));
 sky130_fd_sc_hd__nand4_1 _2154_ (.A(net137),
    .B(_0350_),
    .C(_0347_),
    .D(_0404_),
    .Y(_0415_));
 sky130_fd_sc_hd__clkbuf_2 _2155_ (.A(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__o31ai_1 _2156_ (.A1(_0414_),
    .A2(_0409_),
    .A3(_0416_),
    .B1(net140),
    .Y(_0417_));
 sky130_fd_sc_hd__or4_1 _2157_ (.A(_0414_),
    .B(net140),
    .C(_0409_),
    .D(_0416_),
    .X(_0418_));
 sky130_fd_sc_hd__a21oi_1 _2158_ (.A1(_0417_),
    .A2(_0418_),
    .B1(_0394_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_1 _2159_ (.A(net139),
    .B(net140),
    .Y(_0419_));
 sky130_fd_sc_hd__o31ai_1 _2160_ (.A1(_0409_),
    .A2(_0411_),
    .A3(_0419_),
    .B1(net141),
    .Y(_0420_));
 sky130_fd_sc_hd__or4_1 _2161_ (.A(net141),
    .B(_0409_),
    .C(_0411_),
    .D(_0419_),
    .X(_0421_));
 sky130_fd_sc_hd__a21oi_1 _2162_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0394_),
    .Y(_0127_));
 sky130_fd_sc_hd__and4_1 _2163_ (.A(net138),
    .B(net139),
    .C(net140),
    .D(net141),
    .X(_0422_));
 sky130_fd_sc_hd__nand4_4 _2164_ (.A(_0353_),
    .B(_0373_),
    .C(_0383_),
    .D(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__buf_2 _2165_ (.A(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__o21ai_0 _2166_ (.A1(_0416_),
    .A2(_0424_),
    .B1(net142),
    .Y(_0425_));
 sky130_fd_sc_hd__or3_1 _2167_ (.A(net142),
    .B(_0416_),
    .C(_0424_),
    .X(_0426_));
 sky130_fd_sc_hd__a21oi_1 _2168_ (.A1(_0425_),
    .A2(_0426_),
    .B1(_0394_),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_1 _2169_ (.A(net142),
    .Y(_0427_));
 sky130_fd_sc_hd__o31ai_1 _2170_ (.A1(_0427_),
    .A2(_0411_),
    .A3(_0424_),
    .B1(net143),
    .Y(_0428_));
 sky130_fd_sc_hd__or4_1 _2171_ (.A(_0427_),
    .B(net143),
    .C(_0411_),
    .D(_0423_),
    .X(_0429_));
 sky130_fd_sc_hd__a21oi_1 _2172_ (.A1(_0428_),
    .A2(_0429_),
    .B1(_0394_),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2_1 _2173_ (.A(net142),
    .B(net143),
    .Y(_0430_));
 sky130_fd_sc_hd__o31ai_1 _2174_ (.A1(_0416_),
    .A2(_0424_),
    .A3(_0430_),
    .B1(net144),
    .Y(_0431_));
 sky130_fd_sc_hd__or4_1 _2175_ (.A(net144),
    .B(_0416_),
    .C(_0423_),
    .D(_0430_),
    .X(_0432_));
 sky130_fd_sc_hd__a21oi_1 _2176_ (.A1(_0431_),
    .A2(_0432_),
    .B1(_0394_),
    .Y(_0130_));
 sky130_fd_sc_hd__nand3_1 _2177_ (.A(net142),
    .B(net143),
    .C(net144),
    .Y(_0433_));
 sky130_fd_sc_hd__o31ai_1 _2178_ (.A1(_0411_),
    .A2(_0424_),
    .A3(_0433_),
    .B1(net145),
    .Y(_0434_));
 sky130_fd_sc_hd__or4_1 _2179_ (.A(net145),
    .B(_0411_),
    .C(_0423_),
    .D(_0433_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_4 _2180_ (.A(_1254_),
    .X(_0436_));
 sky130_fd_sc_hd__a21oi_1 _2181_ (.A1(_0434_),
    .A2(_0435_),
    .B1(_0436_),
    .Y(_0131_));
 sky130_fd_sc_hd__nand4_1 _2182_ (.A(net142),
    .B(net143),
    .C(net144),
    .D(net145),
    .Y(_0437_));
 sky130_fd_sc_hd__o31ai_1 _2183_ (.A1(_0416_),
    .A2(_0424_),
    .A3(_0437_),
    .B1(net146),
    .Y(_0438_));
 sky130_fd_sc_hd__or4_1 _2184_ (.A(net146),
    .B(_0416_),
    .C(_0423_),
    .D(_0437_),
    .X(_0439_));
 sky130_fd_sc_hd__a21oi_1 _2185_ (.A1(_0438_),
    .A2(_0439_),
    .B1(_0436_),
    .Y(_0132_));
 sky130_fd_sc_hd__nand3_1 _2186_ (.A(net136),
    .B(_0283_),
    .C(_0398_),
    .Y(_0440_));
 sky130_fd_sc_hd__o21ai_0 _2187_ (.A1(_1399_),
    .A2(_0440_),
    .B1(net147),
    .Y(_0441_));
 sky130_fd_sc_hd__or3_1 _2188_ (.A(net147),
    .B(_1398_),
    .C(_0440_),
    .X(_0442_));
 sky130_fd_sc_hd__a21oi_1 _2189_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0436_),
    .Y(_0133_));
 sky130_fd_sc_hd__and4_1 _2190_ (.A(net142),
    .B(net143),
    .C(net144),
    .D(net145),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _2191_ (.A(net146),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__o31ai_1 _2192_ (.A1(_0411_),
    .A2(_0424_),
    .A3(_0444_),
    .B1(net148),
    .Y(_0445_));
 sky130_fd_sc_hd__or4_1 _2193_ (.A(net148),
    .B(_0410_),
    .C(_0423_),
    .D(_0444_),
    .X(_0446_));
 sky130_fd_sc_hd__a21oi_1 _2194_ (.A1(_0445_),
    .A2(_0446_),
    .B1(_0436_),
    .Y(_0134_));
 sky130_fd_sc_hd__nand3_1 _2195_ (.A(net146),
    .B(net148),
    .C(_0443_),
    .Y(_0447_));
 sky130_fd_sc_hd__o31ai_1 _2196_ (.A1(_0416_),
    .A2(_0424_),
    .A3(_0447_),
    .B1(net149),
    .Y(_0448_));
 sky130_fd_sc_hd__or4_1 _2197_ (.A(net149),
    .B(_0415_),
    .C(_0423_),
    .D(_0447_),
    .X(_0449_));
 sky130_fd_sc_hd__a21oi_1 _2198_ (.A1(_0448_),
    .A2(_0449_),
    .B1(_0436_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand4_1 _2199_ (.A(net146),
    .B(net148),
    .C(net149),
    .D(_0443_),
    .Y(_0450_));
 sky130_fd_sc_hd__o31ai_1 _2200_ (.A1(_0411_),
    .A2(_0424_),
    .A3(_0450_),
    .B1(net150),
    .Y(_0451_));
 sky130_fd_sc_hd__or4_1 _2201_ (.A(net150),
    .B(_0410_),
    .C(_0423_),
    .D(_0450_),
    .X(_0452_));
 sky130_fd_sc_hd__a21oi_1 _2202_ (.A1(_0451_),
    .A2(_0452_),
    .B1(_0436_),
    .Y(_0136_));
 sky130_fd_sc_hd__nor2b_1 _2203_ (.A(_1216_),
    .B_N(net151),
    .Y(_0453_));
 sky130_fd_sc_hd__nor2_1 _2204_ (.A(_1478_),
    .B(net151),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_1 _2205_ (.A(net150),
    .Y(_0455_));
 sky130_fd_sc_hd__nor4_1 _2206_ (.A(_0455_),
    .B(_0416_),
    .C(_0424_),
    .D(_0450_),
    .Y(_0456_));
 sky130_fd_sc_hd__mux2_1 _2207_ (.A0(_0453_),
    .A1(_0454_),
    .S(_0456_),
    .X(_0137_));
 sky130_fd_sc_hd__nand3b_4 _2208_ (.A_N(\prev_event_inc[7] ),
    .B(net12),
    .C(net4),
    .Y(_0457_));
 sky130_fd_sc_hd__xor2_1 _2209_ (.A(net152),
    .B(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__nor2_1 _2210_ (.A(_0366_),
    .B(_0458_),
    .Y(_0138_));
 sky130_fd_sc_hd__mux2i_1 _2211_ (.A0(_1543_),
    .A1(net153),
    .S(_0457_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor2_1 _2212_ (.A(_0366_),
    .B(_0459_),
    .Y(_0139_));
 sky130_fd_sc_hd__and4b_1 _2213_ (.A_N(\prev_event_inc[7] ),
    .B(_1542_),
    .C(net4),
    .D(net12),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_4 _2214_ (.A(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__xnor2_1 _2215_ (.A(net154),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__nor2_1 _2216_ (.A(_0366_),
    .B(_0462_),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_1 _2217_ (.A(net154),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_2 _2218_ (.A(net152),
    .B(net153),
    .Y(_0464_));
 sky130_fd_sc_hd__nor3_1 _2219_ (.A(_0463_),
    .B(_0457_),
    .C(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__xnor2_1 _2220_ (.A(net155),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__nor2_1 _2221_ (.A(_0366_),
    .B(_0466_),
    .Y(_0141_));
 sky130_fd_sc_hd__nand3_1 _2222_ (.A(net154),
    .B(net155),
    .C(_0461_),
    .Y(_0467_));
 sky130_fd_sc_hd__xor2_1 _2223_ (.A(net156),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__nor2_1 _2224_ (.A(_0366_),
    .B(_0468_),
    .Y(_0142_));
 sky130_fd_sc_hd__nand3_2 _2225_ (.A(net154),
    .B(net155),
    .C(net156),
    .Y(_0469_));
 sky130_fd_sc_hd__nor3_1 _2226_ (.A(_0457_),
    .B(_0464_),
    .C(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__xnor2_1 _2227_ (.A(net157),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__nor2_1 _2228_ (.A(_0366_),
    .B(_0471_),
    .Y(_0143_));
 sky130_fd_sc_hd__nand4_1 _2229_ (.A(net136),
    .B(net147),
    .C(_0283_),
    .D(_0398_),
    .Y(_0472_));
 sky130_fd_sc_hd__o31ai_1 _2230_ (.A1(_1266_),
    .A2(_1352_),
    .A3(_0472_),
    .B1(net158),
    .Y(_0473_));
 sky130_fd_sc_hd__or4_1 _2231_ (.A(net158),
    .B(_1354_),
    .C(_1351_),
    .D(_0472_),
    .X(_0474_));
 sky130_fd_sc_hd__a21oi_1 _2232_ (.A1(_0473_),
    .A2(_0474_),
    .B1(_0436_),
    .Y(_0144_));
 sky130_fd_sc_hd__and3_1 _2233_ (.A(net154),
    .B(net155),
    .C(net156),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_2 _2234_ (.A(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__nand3_1 _2235_ (.A(net157),
    .B(_0461_),
    .C(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__xor2_1 _2236_ (.A(net159),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__nor2_1 _2237_ (.A(_0366_),
    .B(_0478_),
    .Y(_0145_));
 sky130_fd_sc_hd__buf_4 _2238_ (.A(_1287_),
    .X(_0479_));
 sky130_fd_sc_hd__nand2_1 _2239_ (.A(net157),
    .B(net159),
    .Y(_0480_));
 sky130_fd_sc_hd__nor4_1 _2240_ (.A(_0457_),
    .B(_0464_),
    .C(_0469_),
    .D(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__xnor2_1 _2241_ (.A(net160),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__nor2_1 _2242_ (.A(_0479_),
    .B(_0482_),
    .Y(_0146_));
 sky130_fd_sc_hd__and3_1 _2243_ (.A(net157),
    .B(net159),
    .C(net160),
    .X(_0483_));
 sky130_fd_sc_hd__nand3_1 _2244_ (.A(_0461_),
    .B(_0476_),
    .C(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__xor2_1 _2245_ (.A(net161),
    .B(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__nor2_1 _2246_ (.A(_0479_),
    .B(_0485_),
    .Y(_0147_));
 sky130_fd_sc_hd__nand4_1 _2247_ (.A(net157),
    .B(net159),
    .C(net160),
    .D(net161),
    .Y(_0486_));
 sky130_fd_sc_hd__nor4_1 _2248_ (.A(_0457_),
    .B(_0464_),
    .C(_0469_),
    .D(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__xnor2_1 _2249_ (.A(net162),
    .B(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_1 _2250_ (.A(_0479_),
    .B(_0488_),
    .Y(_0148_));
 sky130_fd_sc_hd__and4_1 _2251_ (.A(net157),
    .B(net159),
    .C(net160),
    .D(net161),
    .X(_0489_));
 sky130_fd_sc_hd__nand4_1 _2252_ (.A(net162),
    .B(_0461_),
    .C(_0476_),
    .D(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__xor2_1 _2253_ (.A(net163),
    .B(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__nor2_1 _2254_ (.A(_0479_),
    .B(_0491_),
    .Y(_0149_));
 sky130_fd_sc_hd__or2_1 _2255_ (.A(_0457_),
    .B(_0464_),
    .X(_0492_));
 sky130_fd_sc_hd__nand3_2 _2256_ (.A(net162),
    .B(net163),
    .C(_0489_),
    .Y(_0493_));
 sky130_fd_sc_hd__o31ai_1 _2257_ (.A1(_0492_),
    .A2(_0469_),
    .A3(_0493_),
    .B1(net164),
    .Y(_0494_));
 sky130_fd_sc_hd__or4_1 _2258_ (.A(net164),
    .B(_0492_),
    .C(_0469_),
    .D(_0493_),
    .X(_0495_));
 sky130_fd_sc_hd__a21oi_1 _2259_ (.A1(_0494_),
    .A2(_0495_),
    .B1(_0436_),
    .Y(_0150_));
 sky130_fd_sc_hd__nand3_1 _2260_ (.A(net164),
    .B(_0461_),
    .C(_0476_),
    .Y(_0496_));
 sky130_fd_sc_hd__o21ai_0 _2261_ (.A1(_0493_),
    .A2(_0496_),
    .B1(net165),
    .Y(_0497_));
 sky130_fd_sc_hd__or3_1 _2262_ (.A(net165),
    .B(_0493_),
    .C(_0496_),
    .X(_0498_));
 sky130_fd_sc_hd__a21oi_1 _2263_ (.A1(_0497_),
    .A2(_0498_),
    .B1(_0436_),
    .Y(_0151_));
 sky130_fd_sc_hd__and2_0 _2264_ (.A(net164),
    .B(net165),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_1 _2265_ (.A(_0476_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__o31ai_1 _2266_ (.A1(_0492_),
    .A2(_0493_),
    .A3(_0500_),
    .B1(net166),
    .Y(_0501_));
 sky130_fd_sc_hd__or4_1 _2267_ (.A(net166),
    .B(_0492_),
    .C(_0493_),
    .D(_0500_),
    .X(_0502_));
 sky130_fd_sc_hd__a21oi_1 _2268_ (.A1(_0501_),
    .A2(_0502_),
    .B1(_0436_),
    .Y(_0152_));
 sky130_fd_sc_hd__nand2_1 _2269_ (.A(net166),
    .B(_0461_),
    .Y(_0503_));
 sky130_fd_sc_hd__o31ai_1 _2270_ (.A1(_0493_),
    .A2(_0500_),
    .A3(_0503_),
    .B1(net167),
    .Y(_0504_));
 sky130_fd_sc_hd__or4_1 _2271_ (.A(net167),
    .B(_0493_),
    .C(_0500_),
    .D(_0503_),
    .X(_0505_));
 sky130_fd_sc_hd__buf_2 _2272_ (.A(_1254_),
    .X(_0506_));
 sky130_fd_sc_hd__a21oi_1 _2273_ (.A1(_0504_),
    .A2(_0505_),
    .B1(_0506_),
    .Y(_0153_));
 sky130_fd_sc_hd__nand4_1 _2274_ (.A(net162),
    .B(_0476_),
    .C(_0489_),
    .D(_0499_),
    .Y(_0507_));
 sky130_fd_sc_hd__clkbuf_2 _2275_ (.A(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__nand3_1 _2276_ (.A(net163),
    .B(net166),
    .C(net167),
    .Y(_0509_));
 sky130_fd_sc_hd__o31ai_1 _2277_ (.A1(_0492_),
    .A2(_0508_),
    .A3(_0509_),
    .B1(net168),
    .Y(_0510_));
 sky130_fd_sc_hd__or4_1 _2278_ (.A(net168),
    .B(_0492_),
    .C(_0508_),
    .D(_0509_),
    .X(_0511_));
 sky130_fd_sc_hd__a21oi_1 _2279_ (.A1(_0510_),
    .A2(_0511_),
    .B1(_0506_),
    .Y(_0154_));
 sky130_fd_sc_hd__nor2b_1 _2280_ (.A(_1216_),
    .B_N(net169),
    .Y(_0512_));
 sky130_fd_sc_hd__nor2_1 _2281_ (.A(_1478_),
    .B(net169),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_1 _2282_ (.A(net158),
    .Y(_0514_));
 sky130_fd_sc_hd__nor3_1 _2283_ (.A(_0514_),
    .B(_1398_),
    .C(_0472_),
    .Y(_0515_));
 sky130_fd_sc_hd__mux2_1 _2284_ (.A0(_0512_),
    .A1(_0513_),
    .S(_0515_),
    .X(_0155_));
 sky130_fd_sc_hd__and3_1 _2285_ (.A(net163),
    .B(net166),
    .C(net167),
    .X(_0516_));
 sky130_fd_sc_hd__nand3_4 _2286_ (.A(net168),
    .B(_0461_),
    .C(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__buf_2 _2287_ (.A(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__o21ai_0 _2288_ (.A1(_0508_),
    .A2(_0518_),
    .B1(net170),
    .Y(_0519_));
 sky130_fd_sc_hd__or3_1 _2289_ (.A(net170),
    .B(_0508_),
    .C(_0518_),
    .X(_0520_));
 sky130_fd_sc_hd__a21oi_1 _2290_ (.A1(_0519_),
    .A2(_0520_),
    .B1(_0506_),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_1 _2291_ (.A(net170),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_1 _2292_ (.A(net168),
    .Y(_0522_));
 sky130_fd_sc_hd__or4_4 _2293_ (.A(_0522_),
    .B(_0457_),
    .C(_0464_),
    .D(_0509_),
    .X(_0523_));
 sky130_fd_sc_hd__buf_2 _2294_ (.A(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__o31ai_1 _2295_ (.A1(_0521_),
    .A2(_0508_),
    .A3(_0524_),
    .B1(net171),
    .Y(_0525_));
 sky130_fd_sc_hd__or4_1 _2296_ (.A(_0521_),
    .B(net171),
    .C(_0508_),
    .D(_0524_),
    .X(_0526_));
 sky130_fd_sc_hd__a21oi_1 _2297_ (.A1(_0525_),
    .A2(_0526_),
    .B1(_0506_),
    .Y(_0157_));
 sky130_fd_sc_hd__nand2_1 _2298_ (.A(net170),
    .B(net171),
    .Y(_0527_));
 sky130_fd_sc_hd__o31ai_1 _2299_ (.A1(_0508_),
    .A2(_0518_),
    .A3(_0527_),
    .B1(net172),
    .Y(_0528_));
 sky130_fd_sc_hd__or4_1 _2300_ (.A(net172),
    .B(_0508_),
    .C(_0518_),
    .D(_0527_),
    .X(_0529_));
 sky130_fd_sc_hd__a21oi_1 _2301_ (.A1(_0528_),
    .A2(_0529_),
    .B1(_0506_),
    .Y(_0158_));
 sky130_fd_sc_hd__nand3_1 _2302_ (.A(net170),
    .B(net171),
    .C(net172),
    .Y(_0530_));
 sky130_fd_sc_hd__o31ai_1 _2303_ (.A1(_0508_),
    .A2(_0524_),
    .A3(_0530_),
    .B1(net173),
    .Y(_0531_));
 sky130_fd_sc_hd__or4_1 _2304_ (.A(net173),
    .B(_0507_),
    .C(_0523_),
    .D(_0530_),
    .X(_0532_));
 sky130_fd_sc_hd__a21oi_1 _2305_ (.A1(_0531_),
    .A2(_0532_),
    .B1(_0506_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand4_1 _2306_ (.A(net170),
    .B(net171),
    .C(net172),
    .D(net173),
    .Y(_0533_));
 sky130_fd_sc_hd__o31ai_1 _2307_ (.A1(_0508_),
    .A2(_0518_),
    .A3(_0533_),
    .B1(net174),
    .Y(_0534_));
 sky130_fd_sc_hd__or4_1 _2308_ (.A(net174),
    .B(_0507_),
    .C(_0517_),
    .D(_0533_),
    .X(_0535_));
 sky130_fd_sc_hd__a21oi_1 _2309_ (.A1(_0534_),
    .A2(_0535_),
    .B1(_0506_),
    .Y(_0160_));
 sky130_fd_sc_hd__nand4_1 _2310_ (.A(net162),
    .B(net164),
    .C(net165),
    .D(net174),
    .Y(_0536_));
 sky130_fd_sc_hd__or4_1 _2311_ (.A(_0469_),
    .B(_0486_),
    .C(_0533_),
    .D(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_2 _2312_ (.A(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__buf_2 _2313_ (.A(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__o21ai_0 _2314_ (.A1(_0524_),
    .A2(_0539_),
    .B1(net175),
    .Y(_0540_));
 sky130_fd_sc_hd__or3_1 _2315_ (.A(net175),
    .B(_0524_),
    .C(_0538_),
    .X(_0541_));
 sky130_fd_sc_hd__a21oi_1 _2316_ (.A1(_0540_),
    .A2(_0541_),
    .B1(_0506_),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_1 _2317_ (.A(net175),
    .Y(_0542_));
 sky130_fd_sc_hd__o31ai_1 _2318_ (.A1(_0542_),
    .A2(_0518_),
    .A3(_0539_),
    .B1(net176),
    .Y(_0543_));
 sky130_fd_sc_hd__or4_1 _2319_ (.A(_0542_),
    .B(net176),
    .C(_0517_),
    .D(_0538_),
    .X(_0544_));
 sky130_fd_sc_hd__a21oi_1 _2320_ (.A1(_0543_),
    .A2(_0544_),
    .B1(_0506_),
    .Y(_0162_));
 sky130_fd_sc_hd__nand2_1 _2321_ (.A(net175),
    .B(net176),
    .Y(_0545_));
 sky130_fd_sc_hd__o31ai_1 _2322_ (.A1(_0524_),
    .A2(_0539_),
    .A3(_0545_),
    .B1(net177),
    .Y(_0546_));
 sky130_fd_sc_hd__or4_1 _2323_ (.A(net177),
    .B(_0523_),
    .C(_0538_),
    .D(_0545_),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_1 _2324_ (.A1(_0546_),
    .A2(_0547_),
    .B1(_0506_),
    .Y(_0163_));
 sky130_fd_sc_hd__nand3_1 _2325_ (.A(net175),
    .B(net176),
    .C(net177),
    .Y(_0548_));
 sky130_fd_sc_hd__o31ai_1 _2326_ (.A1(_0518_),
    .A2(_0539_),
    .A3(_0548_),
    .B1(net178),
    .Y(_0549_));
 sky130_fd_sc_hd__or4_1 _2327_ (.A(net178),
    .B(_0517_),
    .C(_0538_),
    .D(_0548_),
    .X(_0550_));
 sky130_fd_sc_hd__clkbuf_4 _2328_ (.A(_1254_),
    .X(_0551_));
 sky130_fd_sc_hd__a21oi_1 _2329_ (.A1(_0549_),
    .A2(_0550_),
    .B1(_0551_),
    .Y(_0164_));
 sky130_fd_sc_hd__nor2b_1 _2330_ (.A(_1216_),
    .B_N(net179),
    .Y(_0552_));
 sky130_fd_sc_hd__nor2_1 _2331_ (.A(_1478_),
    .B(net179),
    .Y(_0553_));
 sky130_fd_sc_hd__and4_1 _2332_ (.A(net175),
    .B(net176),
    .C(net177),
    .D(net178),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_2 _2333_ (.A(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__nor3b_1 _2334_ (.A(_0524_),
    .B(_0538_),
    .C_N(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__mux2_1 _2335_ (.A0(_0552_),
    .A1(_0553_),
    .S(_0556_),
    .X(_0165_));
 sky130_fd_sc_hd__and4_1 _2336_ (.A(net136),
    .B(net147),
    .C(net158),
    .D(net169),
    .X(_0557_));
 sky130_fd_sc_hd__nand3_1 _2337_ (.A(_0283_),
    .B(_0398_),
    .C(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__o31ai_1 _2338_ (.A1(_1266_),
    .A2(_1352_),
    .A3(_0558_),
    .B1(net180),
    .Y(_0559_));
 sky130_fd_sc_hd__or4_1 _2339_ (.A(net180),
    .B(_1354_),
    .C(_1351_),
    .D(_0558_),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_1 _2340_ (.A1(_0559_),
    .A2(_0560_),
    .B1(_0551_),
    .Y(_0166_));
 sky130_fd_sc_hd__nand2_1 _2341_ (.A(net179),
    .B(_0555_),
    .Y(_0561_));
 sky130_fd_sc_hd__o31ai_1 _2342_ (.A1(_0518_),
    .A2(_0539_),
    .A3(_0561_),
    .B1(net181),
    .Y(_0562_));
 sky130_fd_sc_hd__or4_1 _2343_ (.A(net181),
    .B(_0517_),
    .C(_0538_),
    .D(_0561_),
    .X(_0563_));
 sky130_fd_sc_hd__a21oi_1 _2344_ (.A1(_0562_),
    .A2(_0563_),
    .B1(_0551_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand3_1 _2345_ (.A(net179),
    .B(net181),
    .C(_0555_),
    .Y(_0564_));
 sky130_fd_sc_hd__o31ai_1 _2346_ (.A1(_0524_),
    .A2(_0539_),
    .A3(_0564_),
    .B1(net182),
    .Y(_0565_));
 sky130_fd_sc_hd__or4_1 _2347_ (.A(net182),
    .B(_0523_),
    .C(_0538_),
    .D(_0564_),
    .X(_0566_));
 sky130_fd_sc_hd__a21oi_1 _2348_ (.A1(_0565_),
    .A2(_0566_),
    .B1(_0551_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand4_1 _2349_ (.A(net179),
    .B(net181),
    .C(net182),
    .D(_0555_),
    .Y(_0567_));
 sky130_fd_sc_hd__o31ai_1 _2350_ (.A1(_0518_),
    .A2(_0539_),
    .A3(_0567_),
    .B1(net183),
    .Y(_0568_));
 sky130_fd_sc_hd__or4_1 _2351_ (.A(net183),
    .B(_0517_),
    .C(_0538_),
    .D(_0567_),
    .X(_0569_));
 sky130_fd_sc_hd__a21oi_1 _2352_ (.A1(_0568_),
    .A2(_0569_),
    .B1(_0551_),
    .Y(_0169_));
 sky130_fd_sc_hd__and4_1 _2353_ (.A(net179),
    .B(net181),
    .C(net182),
    .D(net183),
    .X(_0570_));
 sky130_fd_sc_hd__nand2_1 _2354_ (.A(_0555_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__o31ai_1 _2355_ (.A1(_0524_),
    .A2(_0539_),
    .A3(_0571_),
    .B1(net184),
    .Y(_0572_));
 sky130_fd_sc_hd__or4_1 _2356_ (.A(net184),
    .B(_0523_),
    .C(_0538_),
    .D(_0571_),
    .X(_0573_));
 sky130_fd_sc_hd__a21oi_1 _2357_ (.A1(_0572_),
    .A2(_0573_),
    .B1(_0551_),
    .Y(_0170_));
 sky130_fd_sc_hd__nand3_1 _2358_ (.A(net184),
    .B(_0555_),
    .C(_0570_),
    .Y(_0574_));
 sky130_fd_sc_hd__o31ai_1 _2359_ (.A1(_0518_),
    .A2(_0539_),
    .A3(_0574_),
    .B1(net185),
    .Y(_0575_));
 sky130_fd_sc_hd__or4_1 _2360_ (.A(net185),
    .B(_0517_),
    .C(_0537_),
    .D(_0574_),
    .X(_0576_));
 sky130_fd_sc_hd__a21oi_1 _2361_ (.A1(_0575_),
    .A2(_0576_),
    .B1(_0551_),
    .Y(_0171_));
 sky130_fd_sc_hd__nand4_1 _2362_ (.A(net184),
    .B(net185),
    .C(_0555_),
    .D(_0570_),
    .Y(_0577_));
 sky130_fd_sc_hd__o31ai_1 _2363_ (.A1(_0524_),
    .A2(_0539_),
    .A3(_0577_),
    .B1(net186),
    .Y(_0578_));
 sky130_fd_sc_hd__or4_1 _2364_ (.A(net186),
    .B(_0523_),
    .C(_0537_),
    .D(_0577_),
    .X(_0579_));
 sky130_fd_sc_hd__a21oi_1 _2365_ (.A1(_0578_),
    .A2(_0579_),
    .B1(_0551_),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_1 _2366_ (.A(net180),
    .Y(_0580_));
 sky130_fd_sc_hd__o31ai_1 _2367_ (.A1(_0580_),
    .A2(_1399_),
    .A3(_0558_),
    .B1(net187),
    .Y(_0581_));
 sky130_fd_sc_hd__or4_1 _2368_ (.A(_0580_),
    .B(net187),
    .C(_1398_),
    .D(_0558_),
    .X(_0582_));
 sky130_fd_sc_hd__a21oi_1 _2369_ (.A1(_0581_),
    .A2(_0582_),
    .B1(_0551_),
    .Y(_0173_));
 sky130_fd_sc_hd__and2_0 _2370_ (.A(net180),
    .B(net187),
    .X(_0583_));
 sky130_fd_sc_hd__nand4_4 _2371_ (.A(_0283_),
    .B(_0398_),
    .C(_0557_),
    .D(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__o31ai_1 _2372_ (.A1(_1266_),
    .A2(_1352_),
    .A3(_0584_),
    .B1(net188),
    .Y(_0585_));
 sky130_fd_sc_hd__or4_1 _2373_ (.A(net188),
    .B(_1354_),
    .C(_1351_),
    .D(_0584_),
    .X(_0586_));
 sky130_fd_sc_hd__a21oi_1 _2374_ (.A1(_0585_),
    .A2(_0586_),
    .B1(_0551_),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_1 _2375_ (.A(net188),
    .Y(_0587_));
 sky130_fd_sc_hd__o31ai_1 _2376_ (.A1(_0587_),
    .A2(_1399_),
    .A3(_0584_),
    .B1(net189),
    .Y(_0588_));
 sky130_fd_sc_hd__or4_1 _2377_ (.A(_0587_),
    .B(net189),
    .C(_1398_),
    .D(_0584_),
    .X(_0589_));
 sky130_fd_sc_hd__buf_2 _2378_ (.A(_1254_),
    .X(_0590_));
 sky130_fd_sc_hd__a21oi_1 _2379_ (.A1(_0588_),
    .A2(_0589_),
    .B1(_0590_),
    .Y(_0175_));
 sky130_fd_sc_hd__nor2b_1 _2380_ (.A(_1216_),
    .B_N(net190),
    .Y(_0591_));
 sky130_fd_sc_hd__nor2_1 _2381_ (.A(_1478_),
    .B(net190),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _2382_ (.A(net188),
    .B(net189),
    .Y(_0593_));
 sky130_fd_sc_hd__nor4_1 _2383_ (.A(_1354_),
    .B(_1352_),
    .C(_0584_),
    .D(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__mux2_1 _2384_ (.A0(_0591_),
    .A1(_0592_),
    .S(_0594_),
    .X(_0176_));
 sky130_fd_sc_hd__nand3_1 _2385_ (.A(net188),
    .B(net189),
    .C(net190),
    .Y(_0595_));
 sky130_fd_sc_hd__o31ai_1 _2386_ (.A1(_1399_),
    .A2(_0584_),
    .A3(_0595_),
    .B1(net191),
    .Y(_0596_));
 sky130_fd_sc_hd__or4_1 _2387_ (.A(net191),
    .B(_1398_),
    .C(_0584_),
    .D(_0595_),
    .X(_0597_));
 sky130_fd_sc_hd__a21oi_1 _2388_ (.A1(_0596_),
    .A2(_0597_),
    .B1(_0590_),
    .Y(_0177_));
 sky130_fd_sc_hd__nand2_1 _2389_ (.A(_1540_),
    .B(_1221_),
    .Y(_0598_));
 sky130_fd_sc_hd__xor2_1 _2390_ (.A(net192),
    .B(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_1 _2391_ (.A(_0479_),
    .B(_0599_),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_1 _2392_ (.A(net193),
    .Y(_0600_));
 sky130_fd_sc_hd__nor2_1 _2393_ (.A(_1478_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__nor2_1 _2394_ (.A(_1478_),
    .B(net193),
    .Y(_0602_));
 sky130_fd_sc_hd__nand4_1 _2395_ (.A(net188),
    .B(net189),
    .C(net190),
    .D(net191),
    .Y(_0603_));
 sky130_fd_sc_hd__nor4_1 _2396_ (.A(_1354_),
    .B(_1351_),
    .C(_0584_),
    .D(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__mux2_1 _2397_ (.A0(_0601_),
    .A1(_0602_),
    .S(_0604_),
    .X(_0179_));
 sky130_fd_sc_hd__nor2b_1 _2398_ (.A(_1216_),
    .B_N(net194),
    .Y(_0605_));
 sky130_fd_sc_hd__nor2_1 _2399_ (.A(_1478_),
    .B(net194),
    .Y(_0606_));
 sky130_fd_sc_hd__nor4_1 _2400_ (.A(_0600_),
    .B(_1398_),
    .C(_0584_),
    .D(_0603_),
    .Y(_0607_));
 sky130_fd_sc_hd__mux2_1 _2401_ (.A0(_0605_),
    .A1(_0606_),
    .S(_0607_),
    .X(_0180_));
 sky130_fd_sc_hd__and3b_1 _2402_ (.A_N(\prev_event_inc[1] ),
    .B(net6),
    .C(_1220_),
    .X(_0608_));
 sky130_fd_sc_hd__xnor2_1 _2403_ (.A(net195),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor2_1 _2404_ (.A(_0479_),
    .B(_0609_),
    .Y(_0181_));
 sky130_fd_sc_hd__mux2i_1 _2405_ (.A0(net196),
    .A1(_1539_),
    .S(_0608_),
    .Y(_0610_));
 sky130_fd_sc_hd__nor2_1 _2406_ (.A(_0479_),
    .B(_0610_),
    .Y(_0182_));
 sky130_fd_sc_hd__nand2_1 _2407_ (.A(_1538_),
    .B(_0608_),
    .Y(_0611_));
 sky130_fd_sc_hd__xor2_1 _2408_ (.A(net197),
    .B(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__nor2_1 _2409_ (.A(_0479_),
    .B(_0612_),
    .Y(_0183_));
 sky130_fd_sc_hd__and4b_1 _2410_ (.A_N(\prev_event_inc[1] ),
    .B(net197),
    .C(_1219_),
    .D(net6),
    .X(_0613_));
 sky130_fd_sc_hd__clkbuf_4 _2411_ (.A(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__nand3_1 _2412_ (.A(net195),
    .B(net196),
    .C(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__xor2_1 _2413_ (.A(net198),
    .B(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__nor2_1 _2414_ (.A(_0479_),
    .B(_0616_),
    .Y(_0184_));
 sky130_fd_sc_hd__nand3_1 _2415_ (.A(_1538_),
    .B(net198),
    .C(_0614_),
    .Y(_0617_));
 sky130_fd_sc_hd__xor2_1 _2416_ (.A(net199),
    .B(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__nor2_1 _2417_ (.A(_0479_),
    .B(_0618_),
    .Y(_0185_));
 sky130_fd_sc_hd__buf_4 _2418_ (.A(_1287_),
    .X(_0619_));
 sky130_fd_sc_hd__and3_1 _2419_ (.A(net195),
    .B(net196),
    .C(net199),
    .X(_0620_));
 sky130_fd_sc_hd__nand3_1 _2420_ (.A(net198),
    .B(_0614_),
    .C(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__xor2_1 _2421_ (.A(net200),
    .B(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__nor2_1 _2422_ (.A(_0619_),
    .B(_0622_),
    .Y(_0186_));
 sky130_fd_sc_hd__and3_1 _2423_ (.A(_1538_),
    .B(net198),
    .C(net199),
    .X(_0623_));
 sky130_fd_sc_hd__clkbuf_2 _2424_ (.A(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__nand3_1 _2425_ (.A(net200),
    .B(_0614_),
    .C(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__xor2_1 _2426_ (.A(net201),
    .B(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__nor2_1 _2427_ (.A(_0619_),
    .B(_0626_),
    .Y(_0187_));
 sky130_fd_sc_hd__and4_1 _2428_ (.A(net195),
    .B(net196),
    .C(net198),
    .D(net199),
    .X(_0627_));
 sky130_fd_sc_hd__nand4_1 _2429_ (.A(net200),
    .B(net201),
    .C(_0614_),
    .D(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__xor2_1 _2430_ (.A(net202),
    .B(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__nor2_1 _2431_ (.A(_0619_),
    .B(_0629_),
    .Y(_0188_));
 sky130_fd_sc_hd__xor2_1 _2432_ (.A(net203),
    .B(_1315_),
    .X(_0630_));
 sky130_fd_sc_hd__nor2_1 _2433_ (.A(_0619_),
    .B(_0630_),
    .Y(_0189_));
 sky130_fd_sc_hd__and3_1 _2434_ (.A(net200),
    .B(net201),
    .C(net202),
    .X(_0631_));
 sky130_fd_sc_hd__nand3_1 _2435_ (.A(_0614_),
    .B(_0624_),
    .C(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__xor2_1 _2436_ (.A(net204),
    .B(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__nor2_1 _2437_ (.A(_0619_),
    .B(_0633_),
    .Y(_0190_));
 sky130_fd_sc_hd__and4b_1 _2438_ (.A_N(\prev_event_inc[1] ),
    .B(net199),
    .C(_1219_),
    .D(net6),
    .X(_0634_));
 sky130_fd_sc_hd__and4_1 _2439_ (.A(net195),
    .B(net197),
    .C(net196),
    .D(net198),
    .X(_0635_));
 sky130_fd_sc_hd__and4_2 _2440_ (.A(net200),
    .B(net201),
    .C(net202),
    .D(net204),
    .X(_0636_));
 sky130_fd_sc_hd__nand3_1 _2441_ (.A(_0634_),
    .B(_0635_),
    .C(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__xnor2_1 _2442_ (.A(net205),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__nor2b_1 _2443_ (.A(_1217_),
    .B_N(_0638_),
    .Y(_0191_));
 sky130_fd_sc_hd__nand4_1 _2444_ (.A(net205),
    .B(_0614_),
    .C(_0624_),
    .D(_0636_),
    .Y(_0639_));
 sky130_fd_sc_hd__xor2_1 _2445_ (.A(net206),
    .B(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__nor2_1 _2446_ (.A(_0619_),
    .B(_0640_),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_1 _2447_ (.A(net207),
    .Y(_0641_));
 sky130_fd_sc_hd__and2_1 _2448_ (.A(net205),
    .B(net206),
    .X(_0642_));
 sky130_fd_sc_hd__nand4_4 _2449_ (.A(_0614_),
    .B(_0627_),
    .C(_0636_),
    .D(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__xnor2_1 _2450_ (.A(_0641_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__nor2_1 _2451_ (.A(_0619_),
    .B(_0644_),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2_2 _2452_ (.A(_0614_),
    .B(_0624_),
    .Y(_0645_));
 sky130_fd_sc_hd__nand2_1 _2453_ (.A(_0636_),
    .B(_0642_),
    .Y(_0646_));
 sky130_fd_sc_hd__o31ai_1 _2454_ (.A1(_0641_),
    .A2(_0645_),
    .A3(_0646_),
    .B1(net208),
    .Y(_0647_));
 sky130_fd_sc_hd__or4_1 _2455_ (.A(_0641_),
    .B(net208),
    .C(_0645_),
    .D(_0646_),
    .X(_0648_));
 sky130_fd_sc_hd__a21oi_1 _2456_ (.A1(_0647_),
    .A2(_0648_),
    .B1(_0590_),
    .Y(_0194_));
 sky130_fd_sc_hd__nand2_1 _2457_ (.A(net207),
    .B(net208),
    .Y(_0649_));
 sky130_fd_sc_hd__o21ai_0 _2458_ (.A1(_0643_),
    .A2(_0649_),
    .B1(net209),
    .Y(_0650_));
 sky130_fd_sc_hd__or3_1 _2459_ (.A(net209),
    .B(_0643_),
    .C(_0649_),
    .X(_0651_));
 sky130_fd_sc_hd__a21oi_1 _2460_ (.A1(_0650_),
    .A2(_0651_),
    .B1(_0590_),
    .Y(_0195_));
 sky130_fd_sc_hd__nand3_1 _2461_ (.A(net207),
    .B(net208),
    .C(net209),
    .Y(_0652_));
 sky130_fd_sc_hd__o31ai_1 _2462_ (.A1(_0645_),
    .A2(_0646_),
    .A3(_0652_),
    .B1(net210),
    .Y(_0653_));
 sky130_fd_sc_hd__or4_1 _2463_ (.A(net210),
    .B(_0645_),
    .C(_0646_),
    .D(_0652_),
    .X(_0654_));
 sky130_fd_sc_hd__a21oi_1 _2464_ (.A1(_0653_),
    .A2(_0654_),
    .B1(_0590_),
    .Y(_0196_));
 sky130_fd_sc_hd__nand4_1 _2465_ (.A(net207),
    .B(net208),
    .C(net209),
    .D(net210),
    .Y(_0655_));
 sky130_fd_sc_hd__o21ai_0 _2466_ (.A1(_0643_),
    .A2(_0655_),
    .B1(net211),
    .Y(_0656_));
 sky130_fd_sc_hd__or3_1 _2467_ (.A(net211),
    .B(_0643_),
    .C(_0655_),
    .X(_0657_));
 sky130_fd_sc_hd__a21oi_1 _2468_ (.A1(_0656_),
    .A2(_0657_),
    .B1(_0590_),
    .Y(_0197_));
 sky130_fd_sc_hd__and4_1 _2469_ (.A(net207),
    .B(net208),
    .C(net209),
    .D(net210),
    .X(_0658_));
 sky130_fd_sc_hd__nand2_1 _2470_ (.A(net211),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__o31ai_1 _2471_ (.A1(_0645_),
    .A2(_0646_),
    .A3(_0659_),
    .B1(net212),
    .Y(_0660_));
 sky130_fd_sc_hd__or4_1 _2472_ (.A(net212),
    .B(_0645_),
    .C(_0646_),
    .D(_0659_),
    .X(_0661_));
 sky130_fd_sc_hd__a21oi_1 _2473_ (.A1(_0660_),
    .A2(_0661_),
    .B1(_0590_),
    .Y(_0198_));
 sky130_fd_sc_hd__and2_0 _2474_ (.A(net211),
    .B(net212),
    .X(_0662_));
 sky130_fd_sc_hd__nand2_1 _2475_ (.A(_0658_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__o21ai_0 _2476_ (.A1(_0643_),
    .A2(_0663_),
    .B1(net213),
    .Y(_0664_));
 sky130_fd_sc_hd__or3_1 _2477_ (.A(net213),
    .B(_0643_),
    .C(_0663_),
    .X(_0665_));
 sky130_fd_sc_hd__a21oi_1 _2478_ (.A1(_0664_),
    .A2(_0665_),
    .B1(_0590_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand3_1 _2479_ (.A(_1540_),
    .B(net203),
    .C(_1314_),
    .Y(_0666_));
 sky130_fd_sc_hd__xor2_1 _2480_ (.A(net214),
    .B(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__nor2_1 _2481_ (.A(_0619_),
    .B(_0667_),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_1 _2482_ (.A(net213),
    .Y(_0668_));
 sky130_fd_sc_hd__nand4_4 _2483_ (.A(_0636_),
    .B(_0642_),
    .C(_0658_),
    .D(_0662_),
    .Y(_0669_));
 sky130_fd_sc_hd__buf_2 _2484_ (.A(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__buf_2 _2485_ (.A(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__o31ai_1 _2486_ (.A1(_0668_),
    .A2(_0645_),
    .A3(_0671_),
    .B1(net215),
    .Y(_0672_));
 sky130_fd_sc_hd__or4_1 _2487_ (.A(_0668_),
    .B(net215),
    .C(_0645_),
    .D(_0670_),
    .X(_0673_));
 sky130_fd_sc_hd__a21oi_1 _2488_ (.A1(_0672_),
    .A2(_0673_),
    .B1(_0590_),
    .Y(_0201_));
 sky130_fd_sc_hd__nand2_1 _2489_ (.A(net213),
    .B(net215),
    .Y(_0674_));
 sky130_fd_sc_hd__o31ai_1 _2490_ (.A1(_0643_),
    .A2(_0663_),
    .A3(_0674_),
    .B1(net216),
    .Y(_0675_));
 sky130_fd_sc_hd__or4_1 _2491_ (.A(net216),
    .B(_0643_),
    .C(_0663_),
    .D(_0674_),
    .X(_0676_));
 sky130_fd_sc_hd__a21oi_1 _2492_ (.A1(_0675_),
    .A2(_0676_),
    .B1(_0590_),
    .Y(_0202_));
 sky130_fd_sc_hd__nand3_1 _2493_ (.A(net213),
    .B(net215),
    .C(net216),
    .Y(_0677_));
 sky130_fd_sc_hd__o31ai_1 _2494_ (.A1(_0645_),
    .A2(_0671_),
    .A3(_0677_),
    .B1(net217),
    .Y(_0678_));
 sky130_fd_sc_hd__or4_1 _2495_ (.A(net217),
    .B(_0645_),
    .C(_0670_),
    .D(_0677_),
    .X(_0679_));
 sky130_fd_sc_hd__buf_2 _2496_ (.A(_1254_),
    .X(_0680_));
 sky130_fd_sc_hd__a21oi_1 _2497_ (.A1(_0678_),
    .A2(_0679_),
    .B1(_0680_),
    .Y(_0203_));
 sky130_fd_sc_hd__and4_2 _2498_ (.A(net213),
    .B(net215),
    .C(net216),
    .D(net217),
    .X(_0681_));
 sky130_fd_sc_hd__nand3_4 _2499_ (.A(_0634_),
    .B(_0635_),
    .C(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__o21ai_0 _2500_ (.A1(_0671_),
    .A2(_0682_),
    .B1(net218),
    .Y(_0683_));
 sky130_fd_sc_hd__or3_1 _2501_ (.A(net218),
    .B(_0670_),
    .C(_0682_),
    .X(_0684_));
 sky130_fd_sc_hd__a21oi_1 _2502_ (.A1(_0683_),
    .A2(_0684_),
    .B1(_0680_),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_1 _2503_ (.A(net218),
    .Y(_0685_));
 sky130_fd_sc_hd__nand3_4 _2504_ (.A(_0614_),
    .B(_0624_),
    .C(_0681_),
    .Y(_0686_));
 sky130_fd_sc_hd__o31ai_1 _2505_ (.A1(_0685_),
    .A2(_0671_),
    .A3(_0686_),
    .B1(net219),
    .Y(_0687_));
 sky130_fd_sc_hd__or4_1 _2506_ (.A(_0685_),
    .B(net219),
    .C(_0670_),
    .D(_0686_),
    .X(_0688_));
 sky130_fd_sc_hd__a21oi_1 _2507_ (.A1(_0687_),
    .A2(_0688_),
    .B1(_0680_),
    .Y(_0205_));
 sky130_fd_sc_hd__nand2_1 _2508_ (.A(net218),
    .B(net219),
    .Y(_0689_));
 sky130_fd_sc_hd__o31ai_1 _2509_ (.A1(_0671_),
    .A2(_0682_),
    .A3(_0689_),
    .B1(net220),
    .Y(_0690_));
 sky130_fd_sc_hd__or4_1 _2510_ (.A(net220),
    .B(_0670_),
    .C(_0682_),
    .D(_0689_),
    .X(_0691_));
 sky130_fd_sc_hd__a21oi_1 _2511_ (.A1(_0690_),
    .A2(_0691_),
    .B1(_0680_),
    .Y(_0206_));
 sky130_fd_sc_hd__nand3_1 _2512_ (.A(net218),
    .B(net219),
    .C(net220),
    .Y(_0692_));
 sky130_fd_sc_hd__o31ai_1 _2513_ (.A1(_0671_),
    .A2(_0686_),
    .A3(_0692_),
    .B1(net221),
    .Y(_0693_));
 sky130_fd_sc_hd__or4_1 _2514_ (.A(net221),
    .B(_0670_),
    .C(_0686_),
    .D(_0692_),
    .X(_0694_));
 sky130_fd_sc_hd__a21oi_1 _2515_ (.A1(_0693_),
    .A2(_0694_),
    .B1(_0680_),
    .Y(_0207_));
 sky130_fd_sc_hd__buf_2 _2516_ (.A(net222),
    .X(_0695_));
 sky130_fd_sc_hd__nor2b_1 _2517_ (.A(_1216_),
    .B_N(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__buf_6 _2518_ (.A(_1215_),
    .X(_0697_));
 sky130_fd_sc_hd__nor2_1 _2519_ (.A(_0697_),
    .B(_0695_),
    .Y(_0698_));
 sky130_fd_sc_hd__and4_1 _2520_ (.A(net218),
    .B(net219),
    .C(net220),
    .D(net221),
    .X(_0699_));
 sky130_fd_sc_hd__clkbuf_2 _2521_ (.A(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__nor3b_1 _2522_ (.A(_0670_),
    .B(_0682_),
    .C_N(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(_0696_),
    .A1(_0698_),
    .S(_0701_),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_1 _2524_ (.A(_0695_),
    .B(_0700_),
    .Y(_0702_));
 sky130_fd_sc_hd__o31ai_1 _2525_ (.A1(_0671_),
    .A2(_0686_),
    .A3(_0702_),
    .B1(net223),
    .Y(_0703_));
 sky130_fd_sc_hd__or4_1 _2526_ (.A(net223),
    .B(_0669_),
    .C(_0686_),
    .D(_0702_),
    .X(_0704_));
 sky130_fd_sc_hd__a21oi_1 _2527_ (.A1(_0703_),
    .A2(_0704_),
    .B1(_0680_),
    .Y(_0209_));
 sky130_fd_sc_hd__nand3_1 _2528_ (.A(_0695_),
    .B(net223),
    .C(_0700_),
    .Y(_0705_));
 sky130_fd_sc_hd__o31ai_1 _2529_ (.A1(_0671_),
    .A2(_0682_),
    .A3(_0705_),
    .B1(net224),
    .Y(_0706_));
 sky130_fd_sc_hd__or4_1 _2530_ (.A(net224),
    .B(_0669_),
    .C(_0682_),
    .D(_0705_),
    .X(_0707_));
 sky130_fd_sc_hd__a21oi_1 _2531_ (.A1(_0706_),
    .A2(_0707_),
    .B1(_0680_),
    .Y(_0210_));
 sky130_fd_sc_hd__nand2_1 _2532_ (.A(net203),
    .B(net214),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2_1 _2533_ (.A(net14),
    .B(net125),
    .Y(_0709_));
 sky130_fd_sc_hd__nor3_1 _2534_ (.A(_1262_),
    .B(_0708_),
    .C(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__xnor2_1 _2535_ (.A(net225),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__nor2_1 _2536_ (.A(_0619_),
    .B(_0711_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand4_1 _2537_ (.A(_0695_),
    .B(net223),
    .C(net224),
    .D(_0700_),
    .Y(_0712_));
 sky130_fd_sc_hd__o31ai_1 _2538_ (.A1(_0671_),
    .A2(_0686_),
    .A3(_0712_),
    .B1(net226),
    .Y(_0713_));
 sky130_fd_sc_hd__or4_1 _2539_ (.A(net226),
    .B(_0669_),
    .C(_0686_),
    .D(_0712_),
    .X(_0714_));
 sky130_fd_sc_hd__a21oi_1 _2540_ (.A1(_0713_),
    .A2(_0714_),
    .B1(_0680_),
    .Y(_0212_));
 sky130_fd_sc_hd__and2_0 _2541_ (.A(net224),
    .B(net226),
    .X(_0715_));
 sky130_fd_sc_hd__nand4_1 _2542_ (.A(_0695_),
    .B(net223),
    .C(_0700_),
    .D(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__o31ai_1 _2543_ (.A1(_0671_),
    .A2(_0682_),
    .A3(_0716_),
    .B1(net227),
    .Y(_0717_));
 sky130_fd_sc_hd__or4_1 _2544_ (.A(net227),
    .B(_0669_),
    .C(_0682_),
    .D(_0716_),
    .X(_0718_));
 sky130_fd_sc_hd__a21oi_1 _2545_ (.A1(_0717_),
    .A2(_0718_),
    .B1(_0680_),
    .Y(_0213_));
 sky130_fd_sc_hd__and3_1 _2546_ (.A(net223),
    .B(net224),
    .C(net226),
    .X(_0719_));
 sky130_fd_sc_hd__nand4_1 _2547_ (.A(_0695_),
    .B(net227),
    .C(_0700_),
    .D(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__o31ai_1 _2548_ (.A1(_0670_),
    .A2(_0686_),
    .A3(_0720_),
    .B1(net228),
    .Y(_0721_));
 sky130_fd_sc_hd__or4_1 _2549_ (.A(net228),
    .B(_0669_),
    .C(_0686_),
    .D(_0720_),
    .X(_0722_));
 sky130_fd_sc_hd__a21oi_1 _2550_ (.A1(_0721_),
    .A2(_0722_),
    .B1(_0680_),
    .Y(_0214_));
 sky130_fd_sc_hd__nor2b_1 _2551_ (.A(_1215_),
    .B_N(net229),
    .Y(_0723_));
 sky130_fd_sc_hd__nor2_1 _2552_ (.A(_0697_),
    .B(net229),
    .Y(_0724_));
 sky130_fd_sc_hd__inv_1 _2553_ (.A(net228),
    .Y(_0725_));
 sky130_fd_sc_hd__nor4_1 _2554_ (.A(_0725_),
    .B(_0670_),
    .C(_0682_),
    .D(_0720_),
    .Y(_0726_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0726_),
    .X(_0215_));
 sky130_fd_sc_hd__nand3b_1 _2556_ (.A_N(\prev_event_inc[2] ),
    .B(_1219_),
    .C(net7),
    .Y(_0727_));
 sky130_fd_sc_hd__buf_2 _2557_ (.A(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__nand2_1 _2558_ (.A(net230),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__inv_1 _2559_ (.A(net230),
    .Y(_0730_));
 sky130_fd_sc_hd__and3b_1 _2560_ (.A_N(\prev_event_inc[2] ),
    .B(_1219_),
    .C(net7),
    .X(_0731_));
 sky130_fd_sc_hd__nand2_1 _2561_ (.A(_0730_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__clkbuf_4 _2562_ (.A(_1254_),
    .X(_0733_));
 sky130_fd_sc_hd__a21oi_1 _2563_ (.A1(_0729_),
    .A2(_0732_),
    .B1(_0733_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand2_1 _2564_ (.A(_1553_),
    .B(_0731_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _2565_ (.A(net231),
    .B(_0728_),
    .Y(_0735_));
 sky130_fd_sc_hd__a21oi_1 _2566_ (.A1(_0734_),
    .A2(_0735_),
    .B1(_0733_),
    .Y(_0217_));
 sky130_fd_sc_hd__and4b_2 _2567_ (.A_N(\prev_event_inc[2] ),
    .B(_1219_),
    .C(_1552_),
    .D(net7),
    .X(_0736_));
 sky130_fd_sc_hd__xnor2_1 _2568_ (.A(net232),
    .B(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__nor2_1 _2569_ (.A(_0619_),
    .B(_0737_),
    .Y(_0218_));
 sky130_fd_sc_hd__buf_4 _2570_ (.A(_1287_),
    .X(_0738_));
 sky130_fd_sc_hd__inv_1 _2571_ (.A(net233),
    .Y(_0739_));
 sky130_fd_sc_hd__inv_1 _2572_ (.A(net232),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _2573_ (.A(net231),
    .B(net230),
    .Y(_0741_));
 sky130_fd_sc_hd__or3_1 _2574_ (.A(_0740_),
    .B(_0728_),
    .C(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__xnor2_1 _2575_ (.A(_0739_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__nor2_1 _2576_ (.A(_0738_),
    .B(_0743_),
    .Y(_0219_));
 sky130_fd_sc_hd__nand3_2 _2577_ (.A(net233),
    .B(net232),
    .C(_1552_),
    .Y(_0744_));
 sky130_fd_sc_hd__o21ai_0 _2578_ (.A1(_0728_),
    .A2(_0744_),
    .B1(net234),
    .Y(_0745_));
 sky130_fd_sc_hd__or3_1 _2579_ (.A(net234),
    .B(_0728_),
    .C(_0744_),
    .X(_0746_));
 sky130_fd_sc_hd__a21oi_1 _2580_ (.A1(_0745_),
    .A2(_0746_),
    .B1(_0733_),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_1 _2581_ (.A(net234),
    .Y(_0747_));
 sky130_fd_sc_hd__nand4_2 _2582_ (.A(net233),
    .B(net232),
    .C(net231),
    .D(net230),
    .Y(_0748_));
 sky130_fd_sc_hd__nor3_1 _2583_ (.A(_0747_),
    .B(_0728_),
    .C(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__xnor2_1 _2584_ (.A(net235),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__nor2_1 _2585_ (.A(_0738_),
    .B(_0750_),
    .Y(_0221_));
 sky130_fd_sc_hd__and3_1 _2586_ (.A(net203),
    .B(net214),
    .C(net225),
    .X(_0751_));
 sky130_fd_sc_hd__nand3_1 _2587_ (.A(_1540_),
    .B(_1314_),
    .C(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__xor2_1 _2588_ (.A(net236),
    .B(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__nor2_1 _2589_ (.A(_0738_),
    .B(_0753_),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_1 _2590_ (.A(net235),
    .Y(_0754_));
 sky130_fd_sc_hd__nor4_1 _2591_ (.A(_0754_),
    .B(_0747_),
    .C(_0728_),
    .D(_0744_),
    .Y(_0755_));
 sky130_fd_sc_hd__xnor2_1 _2592_ (.A(net237),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__nor2_1 _2593_ (.A(_0738_),
    .B(_0756_),
    .Y(_0223_));
 sky130_fd_sc_hd__nand3_1 _2594_ (.A(net237),
    .B(net235),
    .C(net234),
    .Y(_0757_));
 sky130_fd_sc_hd__nor3_1 _2595_ (.A(_0728_),
    .B(_0748_),
    .C(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__xnor2_1 _2596_ (.A(net238),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__nor2_1 _2597_ (.A(_0738_),
    .B(_0759_),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_1 _2598_ (.A(net238),
    .Y(_0760_));
 sky130_fd_sc_hd__nor4_1 _2599_ (.A(_0760_),
    .B(_0728_),
    .C(_0744_),
    .D(_0757_),
    .Y(_0761_));
 sky130_fd_sc_hd__xnor2_1 _2600_ (.A(net239),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__nor2_1 _2601_ (.A(_0738_),
    .B(_0762_),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_1 _2602_ (.A(net240),
    .Y(_0763_));
 sky130_fd_sc_hd__inv_1 _2603_ (.A(net239),
    .Y(_0764_));
 sky130_fd_sc_hd__and4_1 _2604_ (.A(net238),
    .B(net237),
    .C(net235),
    .D(net234),
    .X(_0765_));
 sky130_fd_sc_hd__or4b_1 _2605_ (.A(_0764_),
    .B(_0727_),
    .C(_0748_),
    .D_N(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__clkbuf_2 _2606_ (.A(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__xnor2_1 _2607_ (.A(_0763_),
    .B(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__nor2_1 _2608_ (.A(_0738_),
    .B(_0768_),
    .Y(_0226_));
 sky130_fd_sc_hd__or4b_2 _2609_ (.A(_0764_),
    .B(_0728_),
    .C(_0744_),
    .D_N(_0765_),
    .X(_0769_));
 sky130_fd_sc_hd__o21ai_0 _2610_ (.A1(_0763_),
    .A2(_0769_),
    .B1(net241),
    .Y(_0770_));
 sky130_fd_sc_hd__or3_1 _2611_ (.A(net241),
    .B(_0763_),
    .C(_0769_),
    .X(_0771_));
 sky130_fd_sc_hd__a21oi_1 _2612_ (.A1(_0770_),
    .A2(_0771_),
    .B1(_0733_),
    .Y(_0227_));
 sky130_fd_sc_hd__nand2_1 _2613_ (.A(net241),
    .B(net240),
    .Y(_0772_));
 sky130_fd_sc_hd__o21ai_0 _2614_ (.A1(_0767_),
    .A2(_0772_),
    .B1(net242),
    .Y(_0773_));
 sky130_fd_sc_hd__or3_1 _2615_ (.A(net242),
    .B(_0767_),
    .C(_0772_),
    .X(_0774_));
 sky130_fd_sc_hd__a21oi_1 _2616_ (.A1(_0773_),
    .A2(_0774_),
    .B1(_0733_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand3_1 _2617_ (.A(net242),
    .B(net241),
    .C(net240),
    .Y(_0775_));
 sky130_fd_sc_hd__o21ai_0 _2618_ (.A1(_0769_),
    .A2(_0775_),
    .B1(net243),
    .Y(_0776_));
 sky130_fd_sc_hd__or3_1 _2619_ (.A(net243),
    .B(_0769_),
    .C(_0775_),
    .X(_0777_));
 sky130_fd_sc_hd__a21oi_1 _2620_ (.A1(_0776_),
    .A2(_0777_),
    .B1(_0733_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand4_1 _2621_ (.A(net243),
    .B(net242),
    .C(net241),
    .D(net240),
    .Y(_0778_));
 sky130_fd_sc_hd__o21ai_0 _2622_ (.A1(_0767_),
    .A2(_0778_),
    .B1(net244),
    .Y(_0779_));
 sky130_fd_sc_hd__or3_1 _2623_ (.A(net244),
    .B(_0767_),
    .C(_0778_),
    .X(_0780_));
 sky130_fd_sc_hd__a21oi_1 _2624_ (.A1(_0779_),
    .A2(_0780_),
    .B1(_0733_),
    .Y(_0230_));
 sky130_fd_sc_hd__and4_1 _2625_ (.A(net243),
    .B(net242),
    .C(net241),
    .D(net240),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_1 _2626_ (.A(net244),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__o21ai_0 _2627_ (.A1(_0769_),
    .A2(_0782_),
    .B1(net245),
    .Y(_0783_));
 sky130_fd_sc_hd__or3_1 _2628_ (.A(net245),
    .B(_0769_),
    .C(_0782_),
    .X(_0784_));
 sky130_fd_sc_hd__a21oi_1 _2629_ (.A1(_0783_),
    .A2(_0784_),
    .B1(_0733_),
    .Y(_0231_));
 sky130_fd_sc_hd__and2_0 _2630_ (.A(net245),
    .B(net244),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_1 _2631_ (.A(_0781_),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__o21ai_0 _2632_ (.A1(_0767_),
    .A2(_0786_),
    .B1(net246),
    .Y(_0787_));
 sky130_fd_sc_hd__or3_1 _2633_ (.A(net246),
    .B(_0767_),
    .C(_0786_),
    .X(_0788_));
 sky130_fd_sc_hd__a21oi_1 _2634_ (.A1(_0787_),
    .A2(_0788_),
    .B1(_0733_),
    .Y(_0232_));
 sky130_fd_sc_hd__nor3_1 _2635_ (.A(_1262_),
    .B(_1263_),
    .C(_0709_),
    .Y(_0789_));
 sky130_fd_sc_hd__xnor2_1 _2636_ (.A(net247),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__nor2_1 _2637_ (.A(_0738_),
    .B(_0790_),
    .Y(_0233_));
 sky130_fd_sc_hd__and3_1 _2638_ (.A(net246),
    .B(net233),
    .C(net232),
    .X(_0791_));
 sky130_fd_sc_hd__nand2_1 _2639_ (.A(_0736_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand4_2 _2640_ (.A(net239),
    .B(_0765_),
    .C(_0781_),
    .D(_0785_),
    .Y(_0793_));
 sky130_fd_sc_hd__buf_2 _2641_ (.A(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__buf_2 _2642_ (.A(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__o21ai_0 _2643_ (.A1(_0792_),
    .A2(_0795_),
    .B1(net248),
    .Y(_0796_));
 sky130_fd_sc_hd__or3_1 _2644_ (.A(net248),
    .B(_0792_),
    .C(_0794_),
    .X(_0797_));
 sky130_fd_sc_hd__a21oi_1 _2645_ (.A1(_0796_),
    .A2(_0797_),
    .B1(_0733_),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_1 _2646_ (.A(net248),
    .Y(_0798_));
 sky130_fd_sc_hd__nand4_2 _2647_ (.A(net231),
    .B(net230),
    .C(_0731_),
    .D(_0791_),
    .Y(_0799_));
 sky130_fd_sc_hd__o31ai_1 _2648_ (.A1(_0798_),
    .A2(_0795_),
    .A3(_0799_),
    .B1(net249),
    .Y(_0800_));
 sky130_fd_sc_hd__or4_1 _2649_ (.A(net249),
    .B(_0798_),
    .C(_0794_),
    .D(_0799_),
    .X(_0801_));
 sky130_fd_sc_hd__buf_2 _2650_ (.A(_1254_),
    .X(_0802_));
 sky130_fd_sc_hd__a21oi_1 _2651_ (.A1(_0800_),
    .A2(_0801_),
    .B1(_0802_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _2652_ (.A(net249),
    .B(net248),
    .Y(_0803_));
 sky130_fd_sc_hd__o31ai_1 _2653_ (.A1(_0792_),
    .A2(_0795_),
    .A3(_0803_),
    .B1(net250),
    .Y(_0804_));
 sky130_fd_sc_hd__buf_2 _2654_ (.A(_0793_),
    .X(_0805_));
 sky130_fd_sc_hd__or4_1 _2655_ (.A(net250),
    .B(_0792_),
    .C(_0805_),
    .D(_0803_),
    .X(_0806_));
 sky130_fd_sc_hd__a21oi_1 _2656_ (.A1(_0804_),
    .A2(_0806_),
    .B1(_0802_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand3_1 _2657_ (.A(net250),
    .B(net249),
    .C(net248),
    .Y(_0807_));
 sky130_fd_sc_hd__o31ai_1 _2658_ (.A1(_0795_),
    .A2(_0799_),
    .A3(_0807_),
    .B1(net251),
    .Y(_0808_));
 sky130_fd_sc_hd__or4_1 _2659_ (.A(net251),
    .B(_0805_),
    .C(_0799_),
    .D(_0807_),
    .X(_0809_));
 sky130_fd_sc_hd__a21oi_1 _2660_ (.A1(_0808_),
    .A2(_0809_),
    .B1(_0802_),
    .Y(_0237_));
 sky130_fd_sc_hd__nand4_1 _2661_ (.A(net251),
    .B(net250),
    .C(net249),
    .D(net248),
    .Y(_0810_));
 sky130_fd_sc_hd__o31ai_1 _2662_ (.A1(_0792_),
    .A2(_0795_),
    .A3(_0810_),
    .B1(net252),
    .Y(_0811_));
 sky130_fd_sc_hd__or4_1 _2663_ (.A(net252),
    .B(_0792_),
    .C(_0805_),
    .D(_0810_),
    .X(_0812_));
 sky130_fd_sc_hd__a21oi_1 _2664_ (.A1(_0811_),
    .A2(_0812_),
    .B1(_0802_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _2665_ (.A(net252),
    .B(net246),
    .Y(_0813_));
 sky130_fd_sc_hd__or4_2 _2666_ (.A(_0727_),
    .B(_0748_),
    .C(_0810_),
    .D(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__o21ai_0 _2667_ (.A1(_0795_),
    .A2(_0814_),
    .B1(net253),
    .Y(_0815_));
 sky130_fd_sc_hd__or3_1 _2668_ (.A(net253),
    .B(_0794_),
    .C(_0814_),
    .X(_0816_));
 sky130_fd_sc_hd__a21oi_1 _2669_ (.A1(_0815_),
    .A2(_0816_),
    .B1(_0802_),
    .Y(_0239_));
 sky130_fd_sc_hd__inv_1 _2670_ (.A(net253),
    .Y(_0817_));
 sky130_fd_sc_hd__and4_1 _2671_ (.A(net251),
    .B(net250),
    .C(net249),
    .D(net248),
    .X(_0818_));
 sky130_fd_sc_hd__nand4_4 _2672_ (.A(net252),
    .B(_0736_),
    .C(_0791_),
    .D(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__o31ai_1 _2673_ (.A1(_0817_),
    .A2(_0795_),
    .A3(_0819_),
    .B1(net254),
    .Y(_0820_));
 sky130_fd_sc_hd__or4_1 _2674_ (.A(net254),
    .B(_0817_),
    .C(_0805_),
    .D(_0819_),
    .X(_0821_));
 sky130_fd_sc_hd__a21oi_1 _2675_ (.A1(_0820_),
    .A2(_0821_),
    .B1(_0802_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand4_1 _2676_ (.A(net252),
    .B(net246),
    .C(net233),
    .D(net232),
    .Y(_0822_));
 sky130_fd_sc_hd__or4_4 _2677_ (.A(_0727_),
    .B(_0741_),
    .C(_0810_),
    .D(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_1 _2678_ (.A(net254),
    .B(net253),
    .Y(_0824_));
 sky130_fd_sc_hd__o31ai_1 _2679_ (.A1(_0795_),
    .A2(_0823_),
    .A3(_0824_),
    .B1(net255),
    .Y(_0825_));
 sky130_fd_sc_hd__or4_1 _2680_ (.A(net255),
    .B(_0805_),
    .C(_0823_),
    .D(_0824_),
    .X(_0826_));
 sky130_fd_sc_hd__a21oi_1 _2681_ (.A1(_0825_),
    .A2(_0826_),
    .B1(_0802_),
    .Y(_0241_));
 sky130_fd_sc_hd__nand3_1 _2682_ (.A(net255),
    .B(net254),
    .C(net253),
    .Y(_0827_));
 sky130_fd_sc_hd__o31ai_1 _2683_ (.A1(_0795_),
    .A2(_0819_),
    .A3(_0827_),
    .B1(net256),
    .Y(_0828_));
 sky130_fd_sc_hd__or4_1 _2684_ (.A(net256),
    .B(_0805_),
    .C(_0819_),
    .D(_0827_),
    .X(_0829_));
 sky130_fd_sc_hd__a21oi_1 _2685_ (.A1(_0828_),
    .A2(_0829_),
    .B1(_0802_),
    .Y(_0242_));
 sky130_fd_sc_hd__clkbuf_2 _2686_ (.A(net257),
    .X(_0830_));
 sky130_fd_sc_hd__inv_1 _2687_ (.A(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__nor2_1 _2688_ (.A(_1478_),
    .B(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__nor2_1 _2689_ (.A(_0697_),
    .B(_0830_),
    .Y(_0833_));
 sky130_fd_sc_hd__inv_1 _2690_ (.A(net256),
    .Y(_0834_));
 sky130_fd_sc_hd__nor4_1 _2691_ (.A(_0834_),
    .B(_0794_),
    .C(_0814_),
    .D(_0827_),
    .Y(_0835_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(_0832_),
    .A1(_0833_),
    .S(_0835_),
    .X(_0243_));
 sky130_fd_sc_hd__nand4_1 _2693_ (.A(_1540_),
    .B(net247),
    .C(_1314_),
    .D(_1311_),
    .Y(_0836_));
 sky130_fd_sc_hd__xor2_1 _2694_ (.A(net258),
    .B(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__nor2_1 _2695_ (.A(_0738_),
    .B(_0837_),
    .Y(_0244_));
 sky130_fd_sc_hd__and4_1 _2696_ (.A(net255),
    .B(net254),
    .C(net253),
    .D(net256),
    .X(_0838_));
 sky130_fd_sc_hd__clkbuf_2 _2697_ (.A(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__nand2_1 _2698_ (.A(_0830_),
    .B(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__o31ai_1 _2699_ (.A1(_0795_),
    .A2(_0819_),
    .A3(_0840_),
    .B1(net259),
    .Y(_0841_));
 sky130_fd_sc_hd__or4_1 _2700_ (.A(net259),
    .B(_0805_),
    .C(_0819_),
    .D(_0840_),
    .X(_0842_));
 sky130_fd_sc_hd__a21oi_1 _2701_ (.A1(_0841_),
    .A2(_0842_),
    .B1(_0802_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand3_1 _2702_ (.A(_0830_),
    .B(net259),
    .C(_0839_),
    .Y(_0843_));
 sky130_fd_sc_hd__o31ai_1 _2703_ (.A1(_0794_),
    .A2(_0823_),
    .A3(_0843_),
    .B1(net260),
    .Y(_0844_));
 sky130_fd_sc_hd__or4_1 _2704_ (.A(net260),
    .B(_0805_),
    .C(_0823_),
    .D(_0843_),
    .X(_0845_));
 sky130_fd_sc_hd__a21oi_1 _2705_ (.A1(_0844_),
    .A2(_0845_),
    .B1(_0802_),
    .Y(_0246_));
 sky130_fd_sc_hd__nand4_1 _2706_ (.A(_0830_),
    .B(net259),
    .C(net260),
    .D(_0839_),
    .Y(_0846_));
 sky130_fd_sc_hd__o31ai_1 _2707_ (.A1(_0794_),
    .A2(_0819_),
    .A3(_0846_),
    .B1(net261),
    .Y(_0847_));
 sky130_fd_sc_hd__or4_1 _2708_ (.A(net261),
    .B(_0805_),
    .C(_0819_),
    .D(_0846_),
    .X(_0848_));
 sky130_fd_sc_hd__a21oi_1 _2709_ (.A1(_0847_),
    .A2(_0848_),
    .B1(_1217_),
    .Y(_0247_));
 sky130_fd_sc_hd__and4_1 _2710_ (.A(_0830_),
    .B(net259),
    .C(net260),
    .D(net261),
    .X(_0849_));
 sky130_fd_sc_hd__nand2_1 _2711_ (.A(_0839_),
    .B(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__o31ai_1 _2712_ (.A1(_0794_),
    .A2(_0823_),
    .A3(_0850_),
    .B1(net262),
    .Y(_0851_));
 sky130_fd_sc_hd__or4_1 _2713_ (.A(net262),
    .B(_0805_),
    .C(_0823_),
    .D(_0850_),
    .X(_0852_));
 sky130_fd_sc_hd__a21oi_1 _2714_ (.A1(_0851_),
    .A2(_0852_),
    .B1(_1217_),
    .Y(_0248_));
 sky130_fd_sc_hd__and4_1 _2715_ (.A(net259),
    .B(net260),
    .C(net261),
    .D(net262),
    .X(_0853_));
 sky130_fd_sc_hd__nand3_1 _2716_ (.A(_0830_),
    .B(_0839_),
    .C(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__o31ai_1 _2717_ (.A1(_0794_),
    .A2(_0819_),
    .A3(_0854_),
    .B1(net263),
    .Y(_0855_));
 sky130_fd_sc_hd__or4_1 _2718_ (.A(net263),
    .B(_0793_),
    .C(_0819_),
    .D(_0854_),
    .X(_0856_));
 sky130_fd_sc_hd__a21oi_1 _2719_ (.A1(_0855_),
    .A2(_0856_),
    .B1(_1217_),
    .Y(_0249_));
 sky130_fd_sc_hd__nand4_1 _2720_ (.A(_0830_),
    .B(net263),
    .C(_0839_),
    .D(_0853_),
    .Y(_0857_));
 sky130_fd_sc_hd__o31ai_1 _2721_ (.A1(_0794_),
    .A2(_0814_),
    .A3(_0857_),
    .B1(net264),
    .Y(_0858_));
 sky130_fd_sc_hd__or4_1 _2722_ (.A(net264),
    .B(_0793_),
    .C(_0814_),
    .D(_0857_),
    .X(_0859_));
 sky130_fd_sc_hd__a21oi_1 _2723_ (.A1(_0858_),
    .A2(_0859_),
    .B1(_1217_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand3b_1 _2724_ (.A_N(\prev_event_inc[3] ),
    .B(net8),
    .C(_1220_),
    .Y(_0860_));
 sky130_fd_sc_hd__xor2_1 _2725_ (.A(net265),
    .B(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__nor2_1 _2726_ (.A(_0738_),
    .B(_0861_),
    .Y(_0251_));
 sky130_fd_sc_hd__mux2i_1 _2727_ (.A0(_1551_),
    .A1(net266),
    .S(_0860_),
    .Y(_0862_));
 sky130_fd_sc_hd__nor2_1 _2728_ (.A(_1255_),
    .B(_0862_),
    .Y(_0252_));
 sky130_fd_sc_hd__nand4b_1 _2729_ (.A_N(\prev_event_inc[3] ),
    .B(_1550_),
    .C(_1220_),
    .D(net8),
    .Y(_0863_));
 sky130_fd_sc_hd__xor2_1 _2730_ (.A(net267),
    .B(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__nor2_1 _2731_ (.A(_1255_),
    .B(_0864_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand3_1 _2732_ (.A(net265),
    .B(net266),
    .C(_1228_),
    .Y(_0865_));
 sky130_fd_sc_hd__xor2_1 _2733_ (.A(net268),
    .B(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__nor2_1 _2734_ (.A(_1255_),
    .B(_0866_),
    .Y(_0254_));
 sky130_fd_sc_hd__nor4_1 _2735_ (.A(_1262_),
    .B(_1263_),
    .C(_1264_),
    .D(_0709_),
    .Y(_0867_));
 sky130_fd_sc_hd__xnor2_1 _2736_ (.A(net269),
    .B(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__nor2_1 _2737_ (.A(_1255_),
    .B(_0868_),
    .Y(_0255_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(net5),
    .A1(\prev_event_inc[0] ),
    .S(_0697_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _2739_ (.A0(net6),
    .A1(\prev_event_inc[1] ),
    .S(_0697_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2740_ (.A0(net7),
    .A1(\prev_event_inc[2] ),
    .S(_0697_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _2741_ (.A0(net8),
    .A1(\prev_event_inc[3] ),
    .S(_0697_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _2742_ (.A0(net9),
    .A1(\prev_event_inc[4] ),
    .S(_0697_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _2743_ (.A0(net10),
    .A1(\prev_event_inc[5] ),
    .S(_0697_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(net11),
    .A1(\prev_event_inc[6] ),
    .S(_0697_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(net12),
    .A1(\prev_event_inc[7] ),
    .S(_1216_),
    .X(_0263_));
 sky130_fd_sc_hd__buf_2 _2746_ (.A(counter_sel[4]),
    .X(_0869_));
 sky130_fd_sc_hd__clkbuf_4 _2747_ (.A(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__buf_2 _2748_ (.A(counter_sel[2]),
    .X(_0871_));
 sky130_fd_sc_hd__buf_2 _2749_ (.A(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__buf_2 _2750_ (.A(counter_sel[1]),
    .X(_0873_));
 sky130_fd_sc_hd__clkbuf_2 _2751_ (.A(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__buf_2 _2752_ (.A(net1),
    .X(_0875_));
 sky130_fd_sc_hd__nand3b_1 _2753_ (.A_N(_0874_),
    .B(_0875_),
    .C(net14),
    .Y(_0876_));
 sky130_fd_sc_hd__buf_2 _2754_ (.A(_0871_),
    .X(_0877_));
 sky130_fd_sc_hd__a21oi_1 _2755_ (.A1(net195),
    .A2(_0874_),
    .B1(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__clkbuf_4 _2756_ (.A(counter_sel[3]),
    .X(_0879_));
 sky130_fd_sc_hd__buf_2 _2757_ (.A(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__a221o_1 _2758_ (.A1(_0730_),
    .A2(_0872_),
    .B1(_0876_),
    .B2(_0878_),
    .C1(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__buf_2 _2759_ (.A(_0879_),
    .X(_0882_));
 sky130_fd_sc_hd__buf_2 _2760_ (.A(_0869_),
    .X(_0883_));
 sky130_fd_sc_hd__a21oi_1 _2761_ (.A1(net265),
    .A2(_0882_),
    .B1(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__clkbuf_4 _2762_ (.A(counter_sel[5]),
    .X(_0885_));
 sky130_fd_sc_hd__clkbuf_4 _2763_ (.A(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__a221o_1 _2764_ (.A1(_1346_),
    .A2(_0870_),
    .B1(_0881_),
    .B2(_0884_),
    .C1(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__buf_2 _2765_ (.A(_0885_),
    .X(_0888_));
 sky130_fd_sc_hd__nand2_1 _2766_ (.A(net81),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_1 _2767_ (.A(net2),
    .B(net3),
    .Y(_0890_));
 sky130_fd_sc_hd__clkbuf_4 _2768_ (.A(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__buf_2 _2769_ (.A(net2),
    .X(_0892_));
 sky130_fd_sc_hd__nand2b_1 _2770_ (.A_N(net116),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__buf_2 _2771_ (.A(net3),
    .X(_0894_));
 sky130_fd_sc_hd__buf_4 _2772_ (.A(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__mux2i_1 _2773_ (.A0(_0893_),
    .A1(net152),
    .S(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__a31oi_1 _2774_ (.A1(_0887_),
    .A2(_0889_),
    .A3(_0891_),
    .B1(_0896_),
    .Y(net270));
 sky130_fd_sc_hd__buf_2 _2775_ (.A(_0890_),
    .X(_0897_));
 sky130_fd_sc_hd__inv_1 _2776_ (.A(net241),
    .Y(_0898_));
 sky130_fd_sc_hd__clkbuf_2 _2777_ (.A(_0873_),
    .X(_0899_));
 sky130_fd_sc_hd__nand3b_1 _2778_ (.A_N(_0899_),
    .B(_0875_),
    .C(net25),
    .Y(_0900_));
 sky130_fd_sc_hd__a21oi_1 _2779_ (.A1(net206),
    .A2(_0874_),
    .B1(_0877_),
    .Y(_0901_));
 sky130_fd_sc_hd__a221o_1 _2780_ (.A1(_0898_),
    .A2(_0872_),
    .B1(_0900_),
    .B2(_0901_),
    .C1(_0880_),
    .X(_0902_));
 sky130_fd_sc_hd__a21oi_1 _2781_ (.A1(_0882_),
    .A2(net21),
    .B1(_0883_),
    .Y(_0903_));
 sky130_fd_sc_hd__a221o_1 _2782_ (.A1(_0870_),
    .A2(_1387_),
    .B1(_0902_),
    .B2(_0903_),
    .C1(_0886_),
    .X(_0904_));
 sky130_fd_sc_hd__clkbuf_2 _2783_ (.A(_0885_),
    .X(_0905_));
 sky130_fd_sc_hd__nand2_1 _2784_ (.A(_0905_),
    .B(net92),
    .Y(_0906_));
 sky130_fd_sc_hd__nand2b_1 _2785_ (.A_N(net128),
    .B(_0892_),
    .Y(_0907_));
 sky130_fd_sc_hd__mux2i_1 _2786_ (.A0(_0907_),
    .A1(net163),
    .S(_0895_),
    .Y(_0908_));
 sky130_fd_sc_hd__a31oi_1 _2787_ (.A1(_0897_),
    .A2(_0904_),
    .A3(_0906_),
    .B1(_0908_),
    .Y(net271));
 sky130_fd_sc_hd__inv_1 _2788_ (.A(net242),
    .Y(_0909_));
 sky130_fd_sc_hd__nand3b_1 _2789_ (.A_N(_0899_),
    .B(_0875_),
    .C(net36),
    .Y(_0910_));
 sky130_fd_sc_hd__a21oi_1 _2790_ (.A1(net207),
    .A2(_0874_),
    .B1(_0877_),
    .Y(_0911_));
 sky130_fd_sc_hd__a221o_1 _2791_ (.A1(_0909_),
    .A2(_0872_),
    .B1(_0910_),
    .B2(_0911_),
    .C1(_0880_),
    .X(_0912_));
 sky130_fd_sc_hd__a21oi_1 _2792_ (.A1(_0882_),
    .A2(net22),
    .B1(_0883_),
    .Y(_0913_));
 sky130_fd_sc_hd__a221o_1 _2793_ (.A1(_0870_),
    .A2(_1391_),
    .B1(_0912_),
    .B2(_0913_),
    .C1(_0886_),
    .X(_0914_));
 sky130_fd_sc_hd__nand2_1 _2794_ (.A(_0905_),
    .B(net93),
    .Y(_0915_));
 sky130_fd_sc_hd__buf_2 _2795_ (.A(net2),
    .X(_0916_));
 sky130_fd_sc_hd__nand2b_1 _2796_ (.A_N(net129),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__mux2i_1 _2797_ (.A0(_0917_),
    .A1(net164),
    .S(_0895_),
    .Y(_0918_));
 sky130_fd_sc_hd__a31oi_1 _2798_ (.A1(_0897_),
    .A2(_0914_),
    .A3(_0915_),
    .B1(_0918_),
    .Y(net272));
 sky130_fd_sc_hd__inv_1 _2799_ (.A(net59),
    .Y(_0919_));
 sky130_fd_sc_hd__inv_1 _2800_ (.A(net243),
    .Y(_0920_));
 sky130_fd_sc_hd__nand3b_1 _2801_ (.A_N(_0899_),
    .B(_0875_),
    .C(net47),
    .Y(_0921_));
 sky130_fd_sc_hd__a21oi_1 _2802_ (.A1(net208),
    .A2(_0874_),
    .B1(_0877_),
    .Y(_0922_));
 sky130_fd_sc_hd__a221o_1 _2803_ (.A1(_0920_),
    .A2(_0872_),
    .B1(_0921_),
    .B2(_0922_),
    .C1(_0880_),
    .X(_0923_));
 sky130_fd_sc_hd__a21oi_1 _2804_ (.A1(_0882_),
    .A2(net23),
    .B1(_0883_),
    .Y(_0924_));
 sky130_fd_sc_hd__a221o_1 _2805_ (.A1(_0870_),
    .A2(_0919_),
    .B1(_0923_),
    .B2(_0924_),
    .C1(_0886_),
    .X(_0925_));
 sky130_fd_sc_hd__nand2_1 _2806_ (.A(_0905_),
    .B(net94),
    .Y(_0926_));
 sky130_fd_sc_hd__nand2b_1 _2807_ (.A_N(net130),
    .B(_0916_),
    .Y(_0927_));
 sky130_fd_sc_hd__mux2i_1 _2808_ (.A0(_0927_),
    .A1(net165),
    .S(_0895_),
    .Y(_0928_));
 sky130_fd_sc_hd__a31oi_1 _2809_ (.A1(_0897_),
    .A2(_0925_),
    .A3(_0926_),
    .B1(_0928_),
    .Y(net273));
 sky130_fd_sc_hd__inv_1 _2810_ (.A(net60),
    .Y(_0929_));
 sky130_fd_sc_hd__inv_1 _2811_ (.A(net244),
    .Y(_0930_));
 sky130_fd_sc_hd__nand3b_1 _2812_ (.A_N(_0899_),
    .B(_0875_),
    .C(net58),
    .Y(_0931_));
 sky130_fd_sc_hd__a21oi_1 _2813_ (.A1(net209),
    .A2(_0874_),
    .B1(_0877_),
    .Y(_0932_));
 sky130_fd_sc_hd__a221o_1 _2814_ (.A1(_0930_),
    .A2(_0872_),
    .B1(_0931_),
    .B2(_0932_),
    .C1(_0880_),
    .X(_0933_));
 sky130_fd_sc_hd__a21oi_1 _2815_ (.A1(_0882_),
    .A2(net24),
    .B1(_0883_),
    .Y(_0934_));
 sky130_fd_sc_hd__a221o_1 _2816_ (.A1(_0870_),
    .A2(_0929_),
    .B1(_0933_),
    .B2(_0934_),
    .C1(_0886_),
    .X(_0935_));
 sky130_fd_sc_hd__nand2_1 _2817_ (.A(_0905_),
    .B(net95),
    .Y(_0936_));
 sky130_fd_sc_hd__nand2b_1 _2818_ (.A_N(net131),
    .B(_0916_),
    .Y(_0937_));
 sky130_fd_sc_hd__mux2i_1 _2819_ (.A0(_0937_),
    .A1(net166),
    .S(_0895_),
    .Y(_0938_));
 sky130_fd_sc_hd__a31oi_1 _2820_ (.A1(_0897_),
    .A2(_0935_),
    .A3(_0936_),
    .B1(_0938_),
    .Y(net274));
 sky130_fd_sc_hd__inv_1 _2821_ (.A(net245),
    .Y(_0939_));
 sky130_fd_sc_hd__nand3b_1 _2822_ (.A_N(_0899_),
    .B(_0875_),
    .C(net69),
    .Y(_0940_));
 sky130_fd_sc_hd__clkbuf_2 _2823_ (.A(_0873_),
    .X(_0941_));
 sky130_fd_sc_hd__a21oi_1 _2824_ (.A1(net210),
    .A2(_0941_),
    .B1(_0877_),
    .Y(_0942_));
 sky130_fd_sc_hd__a221o_1 _2825_ (.A1(_0939_),
    .A2(_0872_),
    .B1(_0940_),
    .B2(_0942_),
    .C1(_0880_),
    .X(_0943_));
 sky130_fd_sc_hd__a21oi_1 _2826_ (.A1(_0882_),
    .A2(net26),
    .B1(_0883_),
    .Y(_0944_));
 sky130_fd_sc_hd__a221o_1 _2827_ (.A1(_0870_),
    .A2(_1414_),
    .B1(_0943_),
    .B2(_0944_),
    .C1(_0886_),
    .X(_0945_));
 sky130_fd_sc_hd__nand2_1 _2828_ (.A(_0905_),
    .B(net96),
    .Y(_0946_));
 sky130_fd_sc_hd__nand2b_1 _2829_ (.A_N(net132),
    .B(_0916_),
    .Y(_0947_));
 sky130_fd_sc_hd__mux2i_1 _2830_ (.A0(_0947_),
    .A1(net167),
    .S(_0895_),
    .Y(_0948_));
 sky130_fd_sc_hd__a31oi_1 _2831_ (.A1(_0897_),
    .A2(_0945_),
    .A3(_0946_),
    .B1(_0948_),
    .Y(net275));
 sky130_fd_sc_hd__inv_1 _2832_ (.A(net62),
    .Y(_0949_));
 sky130_fd_sc_hd__inv_1 _2833_ (.A(net246),
    .Y(_0950_));
 sky130_fd_sc_hd__nand3b_1 _2834_ (.A_N(_0874_),
    .B(_0875_),
    .C(net80),
    .Y(_0951_));
 sky130_fd_sc_hd__a21oi_1 _2835_ (.A1(net211),
    .A2(_0874_),
    .B1(_0872_),
    .Y(_0952_));
 sky130_fd_sc_hd__a221o_1 _2836_ (.A1(_0950_),
    .A2(_0872_),
    .B1(_0951_),
    .B2(_0952_),
    .C1(_0880_),
    .X(_0953_));
 sky130_fd_sc_hd__a21oi_1 _2837_ (.A1(_0882_),
    .A2(net27),
    .B1(_0883_),
    .Y(_0954_));
 sky130_fd_sc_hd__a221oi_2 _2838_ (.A1(_0870_),
    .A2(_0949_),
    .B1(_0953_),
    .B2(_0954_),
    .C1(_0886_),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _2839_ (.A(_0886_),
    .B(net97),
    .Y(_0956_));
 sky130_fd_sc_hd__nand2_1 _2840_ (.A(_0890_),
    .B(_0956_),
    .Y(_0957_));
 sky130_fd_sc_hd__nor3b_1 _2841_ (.A(net133),
    .B(_0894_),
    .C_N(_0892_),
    .Y(_0958_));
 sky130_fd_sc_hd__a21oi_1 _2842_ (.A1(_0522_),
    .A2(_0895_),
    .B1(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__o21a_1 _2843_ (.A1(_0955_),
    .A2(_0957_),
    .B1(_0959_),
    .X(net276));
 sky130_fd_sc_hd__inv_1 _2844_ (.A(net63),
    .Y(_0960_));
 sky130_fd_sc_hd__buf_2 _2845_ (.A(_0871_),
    .X(_0961_));
 sky130_fd_sc_hd__clkbuf_2 _2846_ (.A(_0873_),
    .X(_0962_));
 sky130_fd_sc_hd__nand3b_1 _2847_ (.A_N(_0962_),
    .B(_0875_),
    .C(net91),
    .Y(_0963_));
 sky130_fd_sc_hd__clkbuf_2 _2848_ (.A(_0871_),
    .X(_0964_));
 sky130_fd_sc_hd__a21oi_1 _2849_ (.A1(net212),
    .A2(_0941_),
    .B1(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__buf_2 _2850_ (.A(_0879_),
    .X(_0966_));
 sky130_fd_sc_hd__a221o_1 _2851_ (.A1(_0798_),
    .A2(_0961_),
    .B1(_0963_),
    .B2(_0965_),
    .C1(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__buf_2 _2852_ (.A(_0869_),
    .X(_0968_));
 sky130_fd_sc_hd__a21oi_1 _2853_ (.A1(_0882_),
    .A2(net28),
    .B1(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__buf_2 _2854_ (.A(_0885_),
    .X(_0970_));
 sky130_fd_sc_hd__a221o_1 _2855_ (.A1(_0870_),
    .A2(_0960_),
    .B1(_0967_),
    .B2(_0969_),
    .C1(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__nand2_1 _2856_ (.A(_0905_),
    .B(net98),
    .Y(_0972_));
 sky130_fd_sc_hd__buf_4 _2857_ (.A(_0894_),
    .X(_0973_));
 sky130_fd_sc_hd__nor3b_1 _2858_ (.A(net134),
    .B(_0894_),
    .C_N(_0892_),
    .Y(_0974_));
 sky130_fd_sc_hd__a21o_1 _2859_ (.A1(_0521_),
    .A2(_0973_),
    .B1(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__a31oi_1 _2860_ (.A1(_0897_),
    .A2(_0971_),
    .A3(_0972_),
    .B1(_0975_),
    .Y(net277));
 sky130_fd_sc_hd__inv_1 _2861_ (.A(net64),
    .Y(_0976_));
 sky130_fd_sc_hd__inv_1 _2862_ (.A(net249),
    .Y(_0977_));
 sky130_fd_sc_hd__nand3b_1 _2863_ (.A_N(_0962_),
    .B(_0875_),
    .C(net102),
    .Y(_0978_));
 sky130_fd_sc_hd__a21oi_1 _2864_ (.A1(net213),
    .A2(_0941_),
    .B1(_0964_),
    .Y(_0979_));
 sky130_fd_sc_hd__a221o_1 _2865_ (.A1(_0977_),
    .A2(_0961_),
    .B1(_0978_),
    .B2(_0979_),
    .C1(_0966_),
    .X(_0980_));
 sky130_fd_sc_hd__a21oi_1 _2866_ (.A1(_0882_),
    .A2(net29),
    .B1(_0968_),
    .Y(_0981_));
 sky130_fd_sc_hd__a221o_1 _2867_ (.A1(_0870_),
    .A2(_0976_),
    .B1(_0980_),
    .B2(_0981_),
    .C1(_0970_),
    .X(_0982_));
 sky130_fd_sc_hd__nand2_1 _2868_ (.A(_0905_),
    .B(net99),
    .Y(_0983_));
 sky130_fd_sc_hd__nand2b_1 _2869_ (.A_N(net135),
    .B(_0916_),
    .Y(_0984_));
 sky130_fd_sc_hd__mux2i_1 _2870_ (.A0(_0984_),
    .A1(net171),
    .S(_0895_),
    .Y(_0985_));
 sky130_fd_sc_hd__a31oi_1 _2871_ (.A1(_0897_),
    .A2(_0982_),
    .A3(_0983_),
    .B1(_0985_),
    .Y(net278));
 sky130_fd_sc_hd__buf_2 _2872_ (.A(_0869_),
    .X(_0986_));
 sky130_fd_sc_hd__inv_1 _2873_ (.A(net65),
    .Y(_0987_));
 sky130_fd_sc_hd__inv_1 _2874_ (.A(net250),
    .Y(_0988_));
 sky130_fd_sc_hd__buf_2 _2875_ (.A(net1),
    .X(_0989_));
 sky130_fd_sc_hd__nand3b_1 _2876_ (.A_N(_0962_),
    .B(_0989_),
    .C(net113),
    .Y(_0990_));
 sky130_fd_sc_hd__a21oi_1 _2877_ (.A1(net215),
    .A2(_0941_),
    .B1(_0964_),
    .Y(_0991_));
 sky130_fd_sc_hd__a221o_1 _2878_ (.A1(_0988_),
    .A2(_0961_),
    .B1(_0990_),
    .B2(_0991_),
    .C1(_0966_),
    .X(_0992_));
 sky130_fd_sc_hd__buf_2 _2879_ (.A(_0879_),
    .X(_0993_));
 sky130_fd_sc_hd__a21oi_1 _2880_ (.A1(_0993_),
    .A2(net30),
    .B1(_0968_),
    .Y(_0994_));
 sky130_fd_sc_hd__a221o_1 _2881_ (.A1(_0986_),
    .A2(_0987_),
    .B1(_0992_),
    .B2(_0994_),
    .C1(_0970_),
    .X(_0995_));
 sky130_fd_sc_hd__nand2_1 _2882_ (.A(_0905_),
    .B(net100),
    .Y(_0996_));
 sky130_fd_sc_hd__nand2b_1 _2883_ (.A_N(net137),
    .B(_0916_),
    .Y(_0997_));
 sky130_fd_sc_hd__mux2i_1 _2884_ (.A0(_0997_),
    .A1(net172),
    .S(_0895_),
    .Y(_0998_));
 sky130_fd_sc_hd__a31oi_1 _2885_ (.A1(_0897_),
    .A2(_0995_),
    .A3(_0996_),
    .B1(_0998_),
    .Y(net279));
 sky130_fd_sc_hd__inv_1 _2886_ (.A(net66),
    .Y(_0999_));
 sky130_fd_sc_hd__inv_1 _2887_ (.A(net251),
    .Y(_1000_));
 sky130_fd_sc_hd__nand3b_1 _2888_ (.A_N(_0962_),
    .B(_0989_),
    .C(net124),
    .Y(_1001_));
 sky130_fd_sc_hd__a21oi_1 _2889_ (.A1(net216),
    .A2(_0941_),
    .B1(_0964_),
    .Y(_1002_));
 sky130_fd_sc_hd__a221o_1 _2890_ (.A1(_1000_),
    .A2(_0961_),
    .B1(_1001_),
    .B2(_1002_),
    .C1(_0966_),
    .X(_1003_));
 sky130_fd_sc_hd__a21oi_1 _2891_ (.A1(_0993_),
    .A2(net31),
    .B1(_0968_),
    .Y(_1004_));
 sky130_fd_sc_hd__a221o_1 _2892_ (.A1(_0986_),
    .A2(_0999_),
    .B1(_1003_),
    .B2(_1004_),
    .C1(_0970_),
    .X(_1005_));
 sky130_fd_sc_hd__nand2_1 _2893_ (.A(_0905_),
    .B(net101),
    .Y(_1006_));
 sky130_fd_sc_hd__nand2b_1 _2894_ (.A_N(net138),
    .B(_0916_),
    .Y(_1007_));
 sky130_fd_sc_hd__buf_4 _2895_ (.A(_0894_),
    .X(_1008_));
 sky130_fd_sc_hd__mux2i_1 _2896_ (.A0(_1007_),
    .A1(net173),
    .S(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__a31oi_1 _2897_ (.A1(_0897_),
    .A2(_1005_),
    .A3(_1006_),
    .B1(_1009_),
    .Y(net280));
 sky130_fd_sc_hd__inv_1 _2898_ (.A(net46),
    .Y(_1010_));
 sky130_fd_sc_hd__inv_1 _2899_ (.A(net231),
    .Y(_1011_));
 sky130_fd_sc_hd__nand3b_1 _2900_ (.A_N(_0962_),
    .B(_0989_),
    .C(net125),
    .Y(_1012_));
 sky130_fd_sc_hd__a21oi_1 _2901_ (.A1(net196),
    .A2(_0941_),
    .B1(_0964_),
    .Y(_1013_));
 sky130_fd_sc_hd__a221o_1 _2902_ (.A1(_1011_),
    .A2(_0961_),
    .B1(_1012_),
    .B2(_1013_),
    .C1(_0966_),
    .X(_1014_));
 sky130_fd_sc_hd__a21oi_1 _2903_ (.A1(_0993_),
    .A2(net266),
    .B1(_0968_),
    .Y(_1015_));
 sky130_fd_sc_hd__a221o_1 _2904_ (.A1(_0986_),
    .A2(_1010_),
    .B1(_1014_),
    .B2(_1015_),
    .C1(_0970_),
    .X(_1016_));
 sky130_fd_sc_hd__nand2_1 _2905_ (.A(_0905_),
    .B(net82),
    .Y(_1017_));
 sky130_fd_sc_hd__nand2b_1 _2906_ (.A_N(net117),
    .B(_0916_),
    .Y(_1018_));
 sky130_fd_sc_hd__mux2i_1 _2907_ (.A0(_1018_),
    .A1(net153),
    .S(_1008_),
    .Y(_1019_));
 sky130_fd_sc_hd__a31oi_1 _2908_ (.A1(_0897_),
    .A2(_1016_),
    .A3(_1017_),
    .B1(_1019_),
    .Y(net281));
 sky130_fd_sc_hd__buf_2 _2909_ (.A(_0890_),
    .X(_1020_));
 sky130_fd_sc_hd__inv_1 _2910_ (.A(net252),
    .Y(_1021_));
 sky130_fd_sc_hd__nand3b_1 _2911_ (.A_N(_0962_),
    .B(_0989_),
    .C(net136),
    .Y(_1022_));
 sky130_fd_sc_hd__a21oi_1 _2912_ (.A1(net217),
    .A2(_0941_),
    .B1(_0964_),
    .Y(_1023_));
 sky130_fd_sc_hd__a221o_1 _2913_ (.A1(_1021_),
    .A2(_0961_),
    .B1(_1022_),
    .B2(_1023_),
    .C1(_0966_),
    .X(_1024_));
 sky130_fd_sc_hd__a21oi_1 _2914_ (.A1(_0993_),
    .A2(net32),
    .B1(_0968_),
    .Y(_1025_));
 sky130_fd_sc_hd__a221o_1 _2915_ (.A1(_0986_),
    .A2(_1437_),
    .B1(_1024_),
    .B2(_1025_),
    .C1(_0970_),
    .X(_1026_));
 sky130_fd_sc_hd__clkbuf_2 _2916_ (.A(_0885_),
    .X(_1027_));
 sky130_fd_sc_hd__nand2_1 _2917_ (.A(_1027_),
    .B(net103),
    .Y(_1028_));
 sky130_fd_sc_hd__nand2_1 _2918_ (.A(_0892_),
    .B(_0414_),
    .Y(_1029_));
 sky130_fd_sc_hd__mux2i_1 _2919_ (.A0(_1029_),
    .A1(net174),
    .S(_1008_),
    .Y(_1030_));
 sky130_fd_sc_hd__a31oi_1 _2920_ (.A1(_1020_),
    .A2(_1026_),
    .A3(_1028_),
    .B1(_1030_),
    .Y(net282));
 sky130_fd_sc_hd__inv_1 _2921_ (.A(net68),
    .Y(_1031_));
 sky130_fd_sc_hd__nand3b_1 _2922_ (.A_N(_0962_),
    .B(_0989_),
    .C(net147),
    .Y(_1032_));
 sky130_fd_sc_hd__a21oi_1 _2923_ (.A1(net218),
    .A2(_0941_),
    .B1(_0964_),
    .Y(_1033_));
 sky130_fd_sc_hd__a221o_1 _2924_ (.A1(_0817_),
    .A2(_0961_),
    .B1(_1032_),
    .B2(_1033_),
    .C1(_0966_),
    .X(_1034_));
 sky130_fd_sc_hd__a21oi_1 _2925_ (.A1(_0993_),
    .A2(net33),
    .B1(_0968_),
    .Y(_1035_));
 sky130_fd_sc_hd__a221o_1 _2926_ (.A1(_0986_),
    .A2(_1031_),
    .B1(_1034_),
    .B2(_1035_),
    .C1(_0970_),
    .X(_1036_));
 sky130_fd_sc_hd__nand2_1 _2927_ (.A(_1027_),
    .B(net104),
    .Y(_1037_));
 sky130_fd_sc_hd__nor3b_1 _2928_ (.A(net140),
    .B(_0894_),
    .C_N(_0892_),
    .Y(_1038_));
 sky130_fd_sc_hd__a21o_1 _2929_ (.A1(_0542_),
    .A2(_0894_),
    .B1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__a31oi_1 _2930_ (.A1(_1020_),
    .A2(_1036_),
    .A3(_1037_),
    .B1(_1039_),
    .Y(net283));
 sky130_fd_sc_hd__inv_1 _2931_ (.A(net70),
    .Y(_1040_));
 sky130_fd_sc_hd__inv_1 _2932_ (.A(net254),
    .Y(_1041_));
 sky130_fd_sc_hd__nand3b_1 _2933_ (.A_N(_0962_),
    .B(_0989_),
    .C(net158),
    .Y(_1042_));
 sky130_fd_sc_hd__a21oi_1 _2934_ (.A1(net219),
    .A2(_0941_),
    .B1(_0964_),
    .Y(_1043_));
 sky130_fd_sc_hd__a221o_1 _2935_ (.A1(_1041_),
    .A2(_0961_),
    .B1(_1042_),
    .B2(_1043_),
    .C1(_0966_),
    .X(_1044_));
 sky130_fd_sc_hd__a21oi_1 _2936_ (.A1(_0993_),
    .A2(net34),
    .B1(_0968_),
    .Y(_1045_));
 sky130_fd_sc_hd__a221o_1 _2937_ (.A1(_0986_),
    .A2(_1040_),
    .B1(_1044_),
    .B2(_1045_),
    .C1(_0970_),
    .X(_1046_));
 sky130_fd_sc_hd__nand2_1 _2938_ (.A(_1027_),
    .B(net105),
    .Y(_1047_));
 sky130_fd_sc_hd__nand2b_1 _2939_ (.A_N(net141),
    .B(_0916_),
    .Y(_1048_));
 sky130_fd_sc_hd__mux2i_1 _2940_ (.A0(_1048_),
    .A1(net176),
    .S(_1008_),
    .Y(_1049_));
 sky130_fd_sc_hd__a31oi_1 _2941_ (.A1(_1020_),
    .A2(_1046_),
    .A3(_1047_),
    .B1(_1049_),
    .Y(net284));
 sky130_fd_sc_hd__inv_1 _2942_ (.A(net255),
    .Y(_1050_));
 sky130_fd_sc_hd__nand3b_1 _2943_ (.A_N(_0962_),
    .B(_0989_),
    .C(net169),
    .Y(_1051_));
 sky130_fd_sc_hd__a21oi_1 _2944_ (.A1(net220),
    .A2(_0941_),
    .B1(_0964_),
    .Y(_1052_));
 sky130_fd_sc_hd__a221o_1 _2945_ (.A1(_1050_),
    .A2(_0961_),
    .B1(_1051_),
    .B2(_1052_),
    .C1(_0966_),
    .X(_1053_));
 sky130_fd_sc_hd__a21oi_1 _2946_ (.A1(_0993_),
    .A2(net35),
    .B1(_0968_),
    .Y(_1054_));
 sky130_fd_sc_hd__a221o_1 _2947_ (.A1(_0986_),
    .A2(_1454_),
    .B1(_1053_),
    .B2(_1054_),
    .C1(_0970_),
    .X(_1055_));
 sky130_fd_sc_hd__nand2_1 _2948_ (.A(_1027_),
    .B(net106),
    .Y(_1056_));
 sky130_fd_sc_hd__nand2_1 _2949_ (.A(_0892_),
    .B(_0427_),
    .Y(_1057_));
 sky130_fd_sc_hd__mux2i_1 _2950_ (.A0(_1057_),
    .A1(net177),
    .S(_1008_),
    .Y(_1058_));
 sky130_fd_sc_hd__a31oi_1 _2951_ (.A1(_1020_),
    .A2(_1055_),
    .A3(_1056_),
    .B1(_1058_),
    .Y(net285));
 sky130_fd_sc_hd__inv_1 _2952_ (.A(net72),
    .Y(_1059_));
 sky130_fd_sc_hd__nand3b_1 _2953_ (.A_N(_0962_),
    .B(_0989_),
    .C(net180),
    .Y(_1060_));
 sky130_fd_sc_hd__clkbuf_2 _2954_ (.A(_0873_),
    .X(_1061_));
 sky130_fd_sc_hd__a21oi_1 _2955_ (.A1(net221),
    .A2(_1061_),
    .B1(_0964_),
    .Y(_1062_));
 sky130_fd_sc_hd__a221o_1 _2956_ (.A1(_0834_),
    .A2(_0961_),
    .B1(_1060_),
    .B2(_1062_),
    .C1(_0966_),
    .X(_1063_));
 sky130_fd_sc_hd__a21oi_1 _2957_ (.A1(_0993_),
    .A2(net37),
    .B1(_0968_),
    .Y(_1064_));
 sky130_fd_sc_hd__a221o_1 _2958_ (.A1(_0986_),
    .A2(_1059_),
    .B1(_1063_),
    .B2(_1064_),
    .C1(_0970_),
    .X(_1065_));
 sky130_fd_sc_hd__nand2_1 _2959_ (.A(_1027_),
    .B(net107),
    .Y(_1066_));
 sky130_fd_sc_hd__nand2b_1 _2960_ (.A_N(net143),
    .B(_0916_),
    .Y(_1067_));
 sky130_fd_sc_hd__mux2i_1 _2961_ (.A0(_1067_),
    .A1(net178),
    .S(_1008_),
    .Y(_1068_));
 sky130_fd_sc_hd__a31oi_1 _2962_ (.A1(_1020_),
    .A2(_1065_),
    .A3(_1066_),
    .B1(_1068_),
    .Y(net286));
 sky130_fd_sc_hd__inv_1 _2963_ (.A(net73),
    .Y(_1069_));
 sky130_fd_sc_hd__buf_2 _2964_ (.A(_0871_),
    .X(_1070_));
 sky130_fd_sc_hd__clkbuf_2 _2965_ (.A(_0873_),
    .X(_1071_));
 sky130_fd_sc_hd__nand3b_1 _2966_ (.A_N(_1071_),
    .B(_0989_),
    .C(net187),
    .Y(_1072_));
 sky130_fd_sc_hd__clkbuf_2 _2967_ (.A(_0871_),
    .X(_1073_));
 sky130_fd_sc_hd__a21oi_1 _2968_ (.A1(_0695_),
    .A2(_1061_),
    .B1(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__buf_2 _2969_ (.A(_0879_),
    .X(_1075_));
 sky130_fd_sc_hd__a221o_1 _2970_ (.A1(_0831_),
    .A2(_1070_),
    .B1(_1072_),
    .B2(_1074_),
    .C1(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__buf_2 _2971_ (.A(_0869_),
    .X(_1077_));
 sky130_fd_sc_hd__a21oi_1 _2972_ (.A1(_0993_),
    .A2(net38),
    .B1(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__buf_2 _2973_ (.A(_0885_),
    .X(_1079_));
 sky130_fd_sc_hd__a221o_1 _2974_ (.A1(_0986_),
    .A2(_1069_),
    .B1(_1076_),
    .B2(_1078_),
    .C1(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__nand2_1 _2975_ (.A(_1027_),
    .B(net108),
    .Y(_1081_));
 sky130_fd_sc_hd__clkbuf_4 _2976_ (.A(net2),
    .X(_1082_));
 sky130_fd_sc_hd__nand2b_1 _2977_ (.A_N(net144),
    .B(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__mux2i_1 _2978_ (.A0(_1083_),
    .A1(net179),
    .S(_1008_),
    .Y(_1084_));
 sky130_fd_sc_hd__a31oi_1 _2979_ (.A1(_1020_),
    .A2(_1080_),
    .A3(_1081_),
    .B1(_1084_),
    .Y(net287));
 sky130_fd_sc_hd__inv_1 _2980_ (.A(net74),
    .Y(_1085_));
 sky130_fd_sc_hd__inv_1 _2981_ (.A(net259),
    .Y(_1086_));
 sky130_fd_sc_hd__nand3b_1 _2982_ (.A_N(_1071_),
    .B(_0989_),
    .C(net188),
    .Y(_1087_));
 sky130_fd_sc_hd__a21oi_1 _2983_ (.A1(net223),
    .A2(_1061_),
    .B1(_1073_),
    .Y(_1088_));
 sky130_fd_sc_hd__a221o_1 _2984_ (.A1(_1086_),
    .A2(_1070_),
    .B1(_1087_),
    .B2(_1088_),
    .C1(_1075_),
    .X(_1089_));
 sky130_fd_sc_hd__a21oi_1 _2985_ (.A1(_0993_),
    .A2(net39),
    .B1(_1077_),
    .Y(_1090_));
 sky130_fd_sc_hd__a221o_1 _2986_ (.A1(_0986_),
    .A2(_1085_),
    .B1(_1089_),
    .B2(_1090_),
    .C1(_1079_),
    .X(_1091_));
 sky130_fd_sc_hd__nand2_1 _2987_ (.A(_1027_),
    .B(net109),
    .Y(_1092_));
 sky130_fd_sc_hd__nand2b_1 _2988_ (.A_N(net145),
    .B(_1082_),
    .Y(_1093_));
 sky130_fd_sc_hd__mux2i_1 _2989_ (.A0(_1093_),
    .A1(net181),
    .S(_1008_),
    .Y(_1094_));
 sky130_fd_sc_hd__a31oi_1 _2990_ (.A1(_1020_),
    .A2(_1091_),
    .A3(_1092_),
    .B1(_1094_),
    .Y(net288));
 sky130_fd_sc_hd__inv_1 _2991_ (.A(net75),
    .Y(_1095_));
 sky130_fd_sc_hd__inv_1 _2992_ (.A(net260),
    .Y(_1096_));
 sky130_fd_sc_hd__nand3b_1 _2993_ (.A_N(_0874_),
    .B(_0875_),
    .C(net189),
    .Y(_1097_));
 sky130_fd_sc_hd__a21oi_1 _2994_ (.A1(net224),
    .A2(_0874_),
    .B1(_0872_),
    .Y(_1098_));
 sky130_fd_sc_hd__a221o_2 _2995_ (.A1(_1096_),
    .A2(_0872_),
    .B1(_1097_),
    .B2(_1098_),
    .C1(_0880_),
    .X(_1099_));
 sky130_fd_sc_hd__a21oi_2 _2996_ (.A1(_0882_),
    .A2(net40),
    .B1(_0883_),
    .Y(_1100_));
 sky130_fd_sc_hd__a221oi_4 _2997_ (.A1(_0870_),
    .A2(_1095_),
    .B1(_1099_),
    .B2(_1100_),
    .C1(_0886_),
    .Y(_1101_));
 sky130_fd_sc_hd__nand2_1 _2998_ (.A(_0886_),
    .B(net110),
    .Y(_1102_));
 sky130_fd_sc_hd__nand2_1 _2999_ (.A(_0890_),
    .B(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__inv_1 _3000_ (.A(net182),
    .Y(_1104_));
 sky130_fd_sc_hd__nor3b_1 _3001_ (.A(net146),
    .B(_0894_),
    .C_N(_0892_),
    .Y(_1105_));
 sky130_fd_sc_hd__a21oi_1 _3002_ (.A1(_1104_),
    .A2(_0895_),
    .B1(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__o21a_1 _3003_ (.A1(_1101_),
    .A2(_1103_),
    .B1(_1106_),
    .X(net289));
 sky130_fd_sc_hd__buf_2 _3004_ (.A(_0869_),
    .X(_1107_));
 sky130_fd_sc_hd__inv_1 _3005_ (.A(net76),
    .Y(_1108_));
 sky130_fd_sc_hd__inv_1 _3006_ (.A(net261),
    .Y(_1109_));
 sky130_fd_sc_hd__buf_2 _3007_ (.A(net1),
    .X(_1110_));
 sky130_fd_sc_hd__nand3b_1 _3008_ (.A_N(_1071_),
    .B(_1110_),
    .C(net190),
    .Y(_1111_));
 sky130_fd_sc_hd__a21oi_1 _3009_ (.A1(net226),
    .A2(_1061_),
    .B1(_1073_),
    .Y(_1112_));
 sky130_fd_sc_hd__a221o_1 _3010_ (.A1(_1109_),
    .A2(_1070_),
    .B1(_1111_),
    .B2(_1112_),
    .C1(_1075_),
    .X(_1113_));
 sky130_fd_sc_hd__buf_2 _3011_ (.A(_0879_),
    .X(_1114_));
 sky130_fd_sc_hd__a21oi_1 _3012_ (.A1(_1114_),
    .A2(net41),
    .B1(_1077_),
    .Y(_1115_));
 sky130_fd_sc_hd__a221o_1 _3013_ (.A1(_1107_),
    .A2(_1108_),
    .B1(_1113_),
    .B2(_1115_),
    .C1(_1079_),
    .X(_1116_));
 sky130_fd_sc_hd__nand2_1 _3014_ (.A(_1027_),
    .B(net111),
    .Y(_1117_));
 sky130_fd_sc_hd__nand2b_1 _3015_ (.A_N(net148),
    .B(_1082_),
    .Y(_1118_));
 sky130_fd_sc_hd__mux2i_1 _3016_ (.A0(_1118_),
    .A1(net183),
    .S(_1008_),
    .Y(_1119_));
 sky130_fd_sc_hd__a31oi_1 _3017_ (.A1(_1020_),
    .A2(_1116_),
    .A3(_1117_),
    .B1(_1119_),
    .Y(net290));
 sky130_fd_sc_hd__inv_1 _3018_ (.A(net77),
    .Y(_1120_));
 sky130_fd_sc_hd__inv_1 _3019_ (.A(net262),
    .Y(_1121_));
 sky130_fd_sc_hd__nand3b_1 _3020_ (.A_N(_1071_),
    .B(_1110_),
    .C(net191),
    .Y(_1122_));
 sky130_fd_sc_hd__a21oi_1 _3021_ (.A1(net227),
    .A2(_1061_),
    .B1(_1073_),
    .Y(_1123_));
 sky130_fd_sc_hd__a221o_1 _3022_ (.A1(_1121_),
    .A2(_1070_),
    .B1(_1122_),
    .B2(_1123_),
    .C1(_1075_),
    .X(_1124_));
 sky130_fd_sc_hd__a21oi_1 _3023_ (.A1(_1114_),
    .A2(net42),
    .B1(_1077_),
    .Y(_1125_));
 sky130_fd_sc_hd__a221o_1 _3024_ (.A1(_1107_),
    .A2(_1120_),
    .B1(_1124_),
    .B2(_1125_),
    .C1(_1079_),
    .X(_1126_));
 sky130_fd_sc_hd__nand2_1 _3025_ (.A(_1027_),
    .B(net112),
    .Y(_1127_));
 sky130_fd_sc_hd__nand2b_1 _3026_ (.A_N(net149),
    .B(_1082_),
    .Y(_1128_));
 sky130_fd_sc_hd__mux2i_1 _3027_ (.A0(_1128_),
    .A1(net184),
    .S(_1008_),
    .Y(_1129_));
 sky130_fd_sc_hd__a31oi_1 _3028_ (.A1(_1020_),
    .A2(_1126_),
    .A3(_1127_),
    .B1(_1129_),
    .Y(net291));
 sky130_fd_sc_hd__nand3b_1 _3029_ (.A_N(_1071_),
    .B(_1110_),
    .C(net192),
    .Y(_1130_));
 sky130_fd_sc_hd__a21oi_1 _3030_ (.A1(net197),
    .A2(_1061_),
    .B1(_1073_),
    .Y(_1131_));
 sky130_fd_sc_hd__a221o_1 _3031_ (.A1(_0740_),
    .A2(_1070_),
    .B1(_1130_),
    .B2(_1131_),
    .C1(_1075_),
    .X(_1132_));
 sky130_fd_sc_hd__a21oi_1 _3032_ (.A1(_1114_),
    .A2(net267),
    .B1(_1077_),
    .Y(_1133_));
 sky130_fd_sc_hd__a221o_1 _3033_ (.A1(_1107_),
    .A2(_1356_),
    .B1(_1132_),
    .B2(_1133_),
    .C1(_1079_),
    .X(_1134_));
 sky130_fd_sc_hd__nand2_1 _3034_ (.A(_1027_),
    .B(net83),
    .Y(_1135_));
 sky130_fd_sc_hd__nor3b_1 _3035_ (.A(net118),
    .B(_0894_),
    .C_N(_0892_),
    .Y(_1136_));
 sky130_fd_sc_hd__a21o_1 _3036_ (.A1(_0463_),
    .A2(_0894_),
    .B1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__a31oi_2 _3037_ (.A1(_1020_),
    .A2(_1134_),
    .A3(_1135_),
    .B1(_1137_),
    .Y(net292));
 sky130_fd_sc_hd__inv_1 _3038_ (.A(net263),
    .Y(_1138_));
 sky130_fd_sc_hd__nand3b_1 _3039_ (.A_N(_1071_),
    .B(_1110_),
    .C(net193),
    .Y(_1139_));
 sky130_fd_sc_hd__a21oi_1 _3040_ (.A1(net228),
    .A2(_1061_),
    .B1(_1073_),
    .Y(_1140_));
 sky130_fd_sc_hd__a221o_1 _3041_ (.A1(_1138_),
    .A2(_1070_),
    .B1(_1139_),
    .B2(_1140_),
    .C1(_1075_),
    .X(_1141_));
 sky130_fd_sc_hd__a21oi_1 _3042_ (.A1(_1114_),
    .A2(net43),
    .B1(_1077_),
    .Y(_1142_));
 sky130_fd_sc_hd__a221o_1 _3043_ (.A1(_1107_),
    .A2(_1480_),
    .B1(_1141_),
    .B2(_1142_),
    .C1(_1079_),
    .X(_1143_));
 sky130_fd_sc_hd__nand2_1 _3044_ (.A(_0888_),
    .B(net114),
    .Y(_1144_));
 sky130_fd_sc_hd__nand2_1 _3045_ (.A(_0892_),
    .B(_0455_),
    .Y(_1145_));
 sky130_fd_sc_hd__mux2i_1 _3046_ (.A0(_1145_),
    .A1(net185),
    .S(_0973_),
    .Y(_1146_));
 sky130_fd_sc_hd__a31oi_1 _3047_ (.A1(_0891_),
    .A2(_1143_),
    .A3(_1144_),
    .B1(_1146_),
    .Y(net293));
 sky130_fd_sc_hd__inv_1 _3048_ (.A(net264),
    .Y(_1147_));
 sky130_fd_sc_hd__nand3b_1 _3049_ (.A_N(_1071_),
    .B(_1110_),
    .C(net194),
    .Y(_1148_));
 sky130_fd_sc_hd__a21oi_1 _3050_ (.A1(net229),
    .A2(_1061_),
    .B1(_1073_),
    .Y(_1149_));
 sky130_fd_sc_hd__a221o_1 _3051_ (.A1(_1147_),
    .A2(_1070_),
    .B1(_1148_),
    .B2(_1149_),
    .C1(_1075_),
    .X(_1150_));
 sky130_fd_sc_hd__a21oi_1 _3052_ (.A1(_1114_),
    .A2(net44),
    .B1(_1077_),
    .Y(_1151_));
 sky130_fd_sc_hd__a221o_1 _3053_ (.A1(_1107_),
    .A2(_1476_),
    .B1(_1150_),
    .B2(_1151_),
    .C1(_1079_),
    .X(_1152_));
 sky130_fd_sc_hd__nand2_1 _3054_ (.A(_0888_),
    .B(net115),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2b_1 _3055_ (.A_N(net151),
    .B(_1082_),
    .Y(_1154_));
 sky130_fd_sc_hd__mux2i_1 _3056_ (.A0(_1154_),
    .A1(net186),
    .S(_0973_),
    .Y(_1155_));
 sky130_fd_sc_hd__a31oi_1 _3057_ (.A1(_0891_),
    .A2(_1152_),
    .A3(_1153_),
    .B1(_1155_),
    .Y(net294));
 sky130_fd_sc_hd__nand3b_1 _3058_ (.A_N(_1071_),
    .B(_1110_),
    .C(net203),
    .Y(_1156_));
 sky130_fd_sc_hd__a21oi_1 _3059_ (.A1(net198),
    .A2(_1061_),
    .B1(_1073_),
    .Y(_1157_));
 sky130_fd_sc_hd__a221o_1 _3060_ (.A1(_0739_),
    .A2(_1070_),
    .B1(_1156_),
    .B2(_1157_),
    .C1(_1075_),
    .X(_1158_));
 sky130_fd_sc_hd__a21oi_1 _3061_ (.A1(_1114_),
    .A2(net268),
    .B1(_1077_),
    .Y(_1159_));
 sky130_fd_sc_hd__a221o_2 _3062_ (.A1(_1107_),
    .A2(_1362_),
    .B1(_1158_),
    .B2(_1159_),
    .C1(_1079_),
    .X(_1160_));
 sky130_fd_sc_hd__nand2_1 _3063_ (.A(_0888_),
    .B(net84),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2b_1 _3064_ (.A_N(net119),
    .B(_1082_),
    .Y(_1162_));
 sky130_fd_sc_hd__mux2i_1 _3065_ (.A0(_1162_),
    .A1(net155),
    .S(_0973_),
    .Y(_1163_));
 sky130_fd_sc_hd__a31oi_1 _3066_ (.A1(_0891_),
    .A2(_1160_),
    .A3(_1161_),
    .B1(_1163_),
    .Y(net295));
 sky130_fd_sc_hd__nand3b_1 _3067_ (.A_N(_1071_),
    .B(_1110_),
    .C(net214),
    .Y(_1164_));
 sky130_fd_sc_hd__a21oi_1 _3068_ (.A1(net199),
    .A2(_1061_),
    .B1(_1073_),
    .Y(_1165_));
 sky130_fd_sc_hd__a221o_1 _3069_ (.A1(_0747_),
    .A2(_1070_),
    .B1(_1164_),
    .B2(_1165_),
    .C1(_1075_),
    .X(_1166_));
 sky130_fd_sc_hd__a21oi_1 _3070_ (.A1(_1114_),
    .A2(net15),
    .B1(_1077_),
    .Y(_1167_));
 sky130_fd_sc_hd__a221o_2 _3071_ (.A1(_1107_),
    .A2(_1367_),
    .B1(_1166_),
    .B2(_1167_),
    .C1(_1079_),
    .X(_1168_));
 sky130_fd_sc_hd__nand2_1 _3072_ (.A(_0888_),
    .B(net85),
    .Y(_1169_));
 sky130_fd_sc_hd__nand2b_1 _3073_ (.A_N(net120),
    .B(_1082_),
    .Y(_1170_));
 sky130_fd_sc_hd__mux2i_1 _3074_ (.A0(_1170_),
    .A1(net156),
    .S(_0973_),
    .Y(_1171_));
 sky130_fd_sc_hd__a31oi_1 _3075_ (.A1(_0891_),
    .A2(_1168_),
    .A3(_1169_),
    .B1(_1171_),
    .Y(net296));
 sky130_fd_sc_hd__nand3b_1 _3076_ (.A_N(_1071_),
    .B(_1110_),
    .C(net225),
    .Y(_1172_));
 sky130_fd_sc_hd__a21oi_1 _3077_ (.A1(net200),
    .A2(_0899_),
    .B1(_1073_),
    .Y(_1173_));
 sky130_fd_sc_hd__a221o_1 _3078_ (.A1(_0754_),
    .A2(_1070_),
    .B1(_1172_),
    .B2(_1173_),
    .C1(_1075_),
    .X(_1174_));
 sky130_fd_sc_hd__a21oi_1 _3079_ (.A1(_1114_),
    .A2(net16),
    .B1(_1077_),
    .Y(_1175_));
 sky130_fd_sc_hd__a221o_2 _3080_ (.A1(_1107_),
    .A2(_1370_),
    .B1(_1174_),
    .B2(_1175_),
    .C1(_1079_),
    .X(_1176_));
 sky130_fd_sc_hd__nand2_1 _3081_ (.A(_0888_),
    .B(net86),
    .Y(_1177_));
 sky130_fd_sc_hd__nand2b_1 _3082_ (.A_N(net121),
    .B(_1082_),
    .Y(_1178_));
 sky130_fd_sc_hd__mux2i_1 _3083_ (.A0(_1178_),
    .A1(net157),
    .S(_0973_),
    .Y(_1179_));
 sky130_fd_sc_hd__a31oi_1 _3084_ (.A1(_0891_),
    .A2(_1176_),
    .A3(_1177_),
    .B1(_1179_),
    .Y(net297));
 sky130_fd_sc_hd__inv_1 _3085_ (.A(net237),
    .Y(_1180_));
 sky130_fd_sc_hd__nand3b_1 _3086_ (.A_N(_0873_),
    .B(_1110_),
    .C(net236),
    .Y(_1181_));
 sky130_fd_sc_hd__a21oi_1 _3087_ (.A1(net201),
    .A2(_0899_),
    .B1(_0871_),
    .Y(_1182_));
 sky130_fd_sc_hd__a221o_1 _3088_ (.A1(_1180_),
    .A2(_0877_),
    .B1(_1181_),
    .B2(_1182_),
    .C1(_0879_),
    .X(_1183_));
 sky130_fd_sc_hd__a21oi_1 _3089_ (.A1(_1114_),
    .A2(net17),
    .B1(_0869_),
    .Y(_1184_));
 sky130_fd_sc_hd__a221o_2 _3090_ (.A1(_1107_),
    .A2(_1373_),
    .B1(_1183_),
    .B2(_1184_),
    .C1(_0885_),
    .X(_1185_));
 sky130_fd_sc_hd__nand2_1 _3091_ (.A(_0888_),
    .B(net87),
    .Y(_1186_));
 sky130_fd_sc_hd__nand2b_1 _3092_ (.A_N(net122),
    .B(_1082_),
    .Y(_1187_));
 sky130_fd_sc_hd__mux2i_1 _3093_ (.A0(_1187_),
    .A1(net159),
    .S(_0973_),
    .Y(_1188_));
 sky130_fd_sc_hd__a31oi_1 _3094_ (.A1(_0891_),
    .A2(_1185_),
    .A3(_1186_),
    .B1(_1188_),
    .Y(net298));
 sky130_fd_sc_hd__inv_1 _3095_ (.A(net53),
    .Y(_1189_));
 sky130_fd_sc_hd__nand3b_1 _3096_ (.A_N(_0873_),
    .B(_1110_),
    .C(net247),
    .Y(_1190_));
 sky130_fd_sc_hd__a21oi_1 _3097_ (.A1(net202),
    .A2(_0899_),
    .B1(_0871_),
    .Y(_1191_));
 sky130_fd_sc_hd__a221o_1 _3098_ (.A1(_0760_),
    .A2(_0877_),
    .B1(_1190_),
    .B2(_1191_),
    .C1(_0879_),
    .X(_1192_));
 sky130_fd_sc_hd__a21oi_1 _3099_ (.A1(_1114_),
    .A2(net18),
    .B1(_0869_),
    .Y(_1193_));
 sky130_fd_sc_hd__a221o_2 _3100_ (.A1(_1107_),
    .A2(_1189_),
    .B1(_1192_),
    .B2(_1193_),
    .C1(_0885_),
    .X(_1194_));
 sky130_fd_sc_hd__nand2_1 _3101_ (.A(_0888_),
    .B(net88),
    .Y(_1195_));
 sky130_fd_sc_hd__nand2b_1 _3102_ (.A_N(net123),
    .B(_1082_),
    .Y(_1196_));
 sky130_fd_sc_hd__mux2i_1 _3103_ (.A0(_1196_),
    .A1(net160),
    .S(_0973_),
    .Y(_1197_));
 sky130_fd_sc_hd__a31oi_1 _3104_ (.A1(_0891_),
    .A2(_1194_),
    .A3(_1195_),
    .B1(_1197_),
    .Y(net299));
 sky130_fd_sc_hd__nand3b_1 _3105_ (.A_N(_0873_),
    .B(net1),
    .C(net258),
    .Y(_1198_));
 sky130_fd_sc_hd__a21oi_1 _3106_ (.A1(net204),
    .A2(_0899_),
    .B1(_0871_),
    .Y(_1199_));
 sky130_fd_sc_hd__a221o_1 _3107_ (.A1(_0764_),
    .A2(_0877_),
    .B1(_1198_),
    .B2(_1199_),
    .C1(_0879_),
    .X(_1200_));
 sky130_fd_sc_hd__a21oi_1 _3108_ (.A1(_0880_),
    .A2(net19),
    .B1(_0869_),
    .Y(_1201_));
 sky130_fd_sc_hd__a221o_2 _3109_ (.A1(_0883_),
    .A2(_1380_),
    .B1(_1200_),
    .B2(_1201_),
    .C1(_0885_),
    .X(_1202_));
 sky130_fd_sc_hd__nand2_1 _3110_ (.A(_0888_),
    .B(net89),
    .Y(_1203_));
 sky130_fd_sc_hd__nand2b_1 _3111_ (.A_N(net126),
    .B(net2),
    .Y(_1204_));
 sky130_fd_sc_hd__mux2i_1 _3112_ (.A0(_1204_),
    .A1(net161),
    .S(_0973_),
    .Y(_1205_));
 sky130_fd_sc_hd__a31oi_1 _3113_ (.A1(_0891_),
    .A2(_1202_),
    .A3(_1203_),
    .B1(_1205_),
    .Y(net300));
 sky130_fd_sc_hd__inv_1 _3114_ (.A(net55),
    .Y(_1206_));
 sky130_fd_sc_hd__nand3b_1 _3115_ (.A_N(_0873_),
    .B(net1),
    .C(net269),
    .Y(_1207_));
 sky130_fd_sc_hd__a21oi_1 _3116_ (.A1(net205),
    .A2(_0899_),
    .B1(_0871_),
    .Y(_1208_));
 sky130_fd_sc_hd__a221o_1 _3117_ (.A1(_0763_),
    .A2(_0877_),
    .B1(_1207_),
    .B2(_1208_),
    .C1(_0879_),
    .X(_1209_));
 sky130_fd_sc_hd__a21oi_1 _3118_ (.A1(_0880_),
    .A2(net20),
    .B1(_0869_),
    .Y(_1210_));
 sky130_fd_sc_hd__a221o_2 _3119_ (.A1(_0883_),
    .A2(_1206_),
    .B1(_1209_),
    .B2(_1210_),
    .C1(_0885_),
    .X(_1211_));
 sky130_fd_sc_hd__nand2_1 _3120_ (.A(_0888_),
    .B(net90),
    .Y(_1212_));
 sky130_fd_sc_hd__nand2b_1 _3121_ (.A_N(net127),
    .B(net2),
    .Y(_1213_));
 sky130_fd_sc_hd__mux2i_1 _3122_ (.A0(_1213_),
    .A1(net162),
    .S(_0973_),
    .Y(_1214_));
 sky130_fd_sc_hd__a31oi_1 _3123_ (.A1(_0891_),
    .A2(_1211_),
    .A3(_1212_),
    .B1(_1214_),
    .Y(net301));
 sky130_fd_sc_hd__ha_1 _3124_ (.A(net195),
    .B(net196),
    .COUT(_1538_),
    .SUM(_1539_));
 sky130_fd_sc_hd__ha_1 _3125_ (.A(net14),
    .B(net125),
    .COUT(_1540_),
    .SUM(_1541_));
 sky130_fd_sc_hd__ha_1 _3126_ (.A(net152),
    .B(net153),
    .COUT(_1542_),
    .SUM(_1543_));
 sky130_fd_sc_hd__ha_2 _3127_ (.A(net116),
    .B(net117),
    .COUT(_1544_),
    .SUM(_1545_));
 sky130_fd_sc_hd__ha_1 _3128_ (.A(net81),
    .B(net82),
    .COUT(_1546_),
    .SUM(_1547_));
 sky130_fd_sc_hd__ha_2 _3129_ (.A(net45),
    .B(net46),
    .COUT(_1548_),
    .SUM(_1549_));
 sky130_fd_sc_hd__ha_1 _3130_ (.A(net265),
    .B(net266),
    .COUT(_1550_),
    .SUM(_1551_));
 sky130_fd_sc_hd__ha_1 _3131_ (.A(net230),
    .B(net231),
    .COUT(_1552_),
    .SUM(_1553_));
 sky130_fd_sc_hd__dfrtp_4 \counters[0]$_DFFE_PN0P_  (.D(_0000_),
    .Q(net14),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[100]$_DFFE_PN0P_  (.D(_0001_),
    .Q(net15),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[101]$_DFFE_PN0P_  (.D(_0002_),
    .Q(net16),
    .RESET_B(net13),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[102]$_DFFE_PN0P_  (.D(_0003_),
    .Q(net17),
    .RESET_B(net13),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[103]$_DFFE_PN0P_  (.D(_0004_),
    .Q(net18),
    .RESET_B(net13),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[104]$_DFFE_PN0P_  (.D(_0005_),
    .Q(net19),
    .RESET_B(net13),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[105]$_DFFE_PN0P_  (.D(_0006_),
    .Q(net20),
    .RESET_B(net13),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[106]$_DFFE_PN0P_  (.D(_0007_),
    .Q(net21),
    .RESET_B(net13),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[107]$_DFFE_PN0P_  (.D(_0008_),
    .Q(net22),
    .RESET_B(net13),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[108]$_DFFE_PN0P_  (.D(_0009_),
    .Q(net23),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[109]$_DFFE_PN0P_  (.D(_0010_),
    .Q(net24),
    .RESET_B(net13),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[10]$_DFFE_PN0P_  (.D(_0011_),
    .Q(net25),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[110]$_DFFE_PN0P_  (.D(_0012_),
    .Q(net26),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[111]$_DFFE_PN0P_  (.D(_0013_),
    .Q(net27),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[112]$_DFFE_PN0P_  (.D(_0014_),
    .Q(net28),
    .RESET_B(net13),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[113]$_DFFE_PN0P_  (.D(_0015_),
    .Q(net29),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[114]$_DFFE_PN0P_  (.D(_0016_),
    .Q(net30),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[115]$_DFFE_PN0P_  (.D(_0017_),
    .Q(net31),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[116]$_DFFE_PN0P_  (.D(_0018_),
    .Q(net32),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[117]$_DFFE_PN0P_  (.D(_0019_),
    .Q(net33),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[118]$_DFFE_PN0P_  (.D(_0020_),
    .Q(net34),
    .RESET_B(net13),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[119]$_DFFE_PN0P_  (.D(_0021_),
    .Q(net35),
    .RESET_B(net13),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[11]$_DFFE_PN0P_  (.D(_0022_),
    .Q(net36),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[120]$_DFFE_PN0P_  (.D(_0023_),
    .Q(net37),
    .RESET_B(net13),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[121]$_DFFE_PN0P_  (.D(_0024_),
    .Q(net38),
    .RESET_B(net13),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[122]$_DFFE_PN0P_  (.D(_0025_),
    .Q(net39),
    .RESET_B(net13),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[123]$_DFFE_PN0P_  (.D(_0026_),
    .Q(net40),
    .RESET_B(net13),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[124]$_DFFE_PN0P_  (.D(_0027_),
    .Q(net41),
    .RESET_B(net13),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[125]$_DFFE_PN0P_  (.D(_0028_),
    .Q(net42),
    .RESET_B(net13),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[126]$_DFFE_PN0P_  (.D(_0029_),
    .Q(net43),
    .RESET_B(net13),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[127]$_DFFE_PN0P_  (.D(_0030_),
    .Q(net44),
    .RESET_B(net13),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[128]$_DFFE_PN0P_  (.D(_0031_),
    .Q(net45),
    .RESET_B(net13),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[129]$_DFFE_PN0P_  (.D(_0032_),
    .Q(net46),
    .RESET_B(net13),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[12]$_DFFE_PN0P_  (.D(_0033_),
    .Q(net47),
    .RESET_B(net13),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[130]$_DFFE_PN0P_  (.D(_0034_),
    .Q(net48),
    .RESET_B(net13),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[131]$_DFFE_PN0P_  (.D(_0035_),
    .Q(net49),
    .RESET_B(net13),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[132]$_DFFE_PN0P_  (.D(_0036_),
    .Q(net50),
    .RESET_B(net13),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[133]$_DFFE_PN0P_  (.D(_0037_),
    .Q(net51),
    .RESET_B(net13),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[134]$_DFFE_PN0P_  (.D(_0038_),
    .Q(net52),
    .RESET_B(net13),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[135]$_DFFE_PN0P_  (.D(_0039_),
    .Q(net53),
    .RESET_B(net13),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[136]$_DFFE_PN0P_  (.D(_0040_),
    .Q(net54),
    .RESET_B(net13),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[137]$_DFFE_PN0P_  (.D(_0041_),
    .Q(net55),
    .RESET_B(net13),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[138]$_DFFE_PN0P_  (.D(_0042_),
    .Q(net56),
    .RESET_B(net13),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[139]$_DFFE_PN0P_  (.D(_0043_),
    .Q(net57),
    .RESET_B(net13),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[13]$_DFFE_PN0P_  (.D(_0044_),
    .Q(net58),
    .RESET_B(net13),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[140]$_DFFE_PN0P_  (.D(_0045_),
    .Q(net59),
    .RESET_B(net13),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[141]$_DFFE_PN0P_  (.D(_0046_),
    .Q(net60),
    .RESET_B(net13),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[142]$_DFFE_PN0P_  (.D(_0047_),
    .Q(net61),
    .RESET_B(net13),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[143]$_DFFE_PN0P_  (.D(_0048_),
    .Q(net62),
    .RESET_B(net13),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[144]$_DFFE_PN0P_  (.D(_0049_),
    .Q(net63),
    .RESET_B(net13),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[145]$_DFFE_PN0P_  (.D(_0050_),
    .Q(net64),
    .RESET_B(net13),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[146]$_DFFE_PN0P_  (.D(_0051_),
    .Q(net65),
    .RESET_B(net13),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[147]$_DFFE_PN0P_  (.D(_0052_),
    .Q(net66),
    .RESET_B(net13),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[148]$_DFFE_PN0P_  (.D(_0053_),
    .Q(net67),
    .RESET_B(net13),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[149]$_DFFE_PN0P_  (.D(_0054_),
    .Q(net68),
    .RESET_B(net13),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[14]$_DFFE_PN0P_  (.D(_0055_),
    .Q(net69),
    .RESET_B(net13),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[150]$_DFFE_PN0P_  (.D(_0056_),
    .Q(net70),
    .RESET_B(net13),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[151]$_DFFE_PN0P_  (.D(_0057_),
    .Q(net71),
    .RESET_B(net13),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[152]$_DFFE_PN0P_  (.D(_0058_),
    .Q(net72),
    .RESET_B(net13),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[153]$_DFFE_PN0P_  (.D(_0059_),
    .Q(net73),
    .RESET_B(net13),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[154]$_DFFE_PN0P_  (.D(_0060_),
    .Q(net74),
    .RESET_B(net13),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[155]$_DFFE_PN0P_  (.D(_0061_),
    .Q(net75),
    .RESET_B(net13),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[156]$_DFFE_PN0P_  (.D(_0062_),
    .Q(net76),
    .RESET_B(net13),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[157]$_DFFE_PN0P_  (.D(_0063_),
    .Q(net77),
    .RESET_B(net13),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[158]$_DFFE_PN0P_  (.D(_0064_),
    .Q(net78),
    .RESET_B(net13),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[159]$_DFFE_PN0P_  (.D(_0065_),
    .Q(net79),
    .RESET_B(net13),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[15]$_DFFE_PN0P_  (.D(_0066_),
    .Q(net80),
    .RESET_B(net13),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[160]$_DFFE_PN0P_  (.D(_0067_),
    .Q(net81),
    .RESET_B(net13),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[161]$_DFFE_PN0P_  (.D(_0068_),
    .Q(net82),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[162]$_DFFE_PN0P_  (.D(_0069_),
    .Q(net83),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[163]$_DFFE_PN0P_  (.D(_0070_),
    .Q(net84),
    .RESET_B(net13),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[164]$_DFFE_PN0P_  (.D(_0071_),
    .Q(net85),
    .RESET_B(net13),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[165]$_DFFE_PN0P_  (.D(_0072_),
    .Q(net86),
    .RESET_B(net13),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[166]$_DFFE_PN0P_  (.D(_0073_),
    .Q(net87),
    .RESET_B(net13),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[167]$_DFFE_PN0P_  (.D(_0074_),
    .Q(net88),
    .RESET_B(net13),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[168]$_DFFE_PN0P_  (.D(_0075_),
    .Q(net89),
    .RESET_B(net13),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[169]$_DFFE_PN0P_  (.D(_0076_),
    .Q(net90),
    .RESET_B(net13),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[16]$_DFFE_PN0P_  (.D(_0077_),
    .Q(net91),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[170]$_DFFE_PN0P_  (.D(_0078_),
    .Q(net92),
    .RESET_B(net13),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[171]$_DFFE_PN0P_  (.D(_0079_),
    .Q(net93),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[172]$_DFFE_PN0P_  (.D(_0080_),
    .Q(net94),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[173]$_DFFE_PN0P_  (.D(_0081_),
    .Q(net95),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[174]$_DFFE_PN0P_  (.D(_0082_),
    .Q(net96),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[175]$_DFFE_PN0P_  (.D(_0083_),
    .Q(net97),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[176]$_DFFE_PN0P_  (.D(_0084_),
    .Q(net98),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[177]$_DFFE_PN0P_  (.D(_0085_),
    .Q(net99),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[178]$_DFFE_PN0P_  (.D(_0086_),
    .Q(net100),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[179]$_DFFE_PN0P_  (.D(_0087_),
    .Q(net101),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[17]$_DFFE_PN0P_  (.D(_0088_),
    .Q(net102),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[180]$_DFFE_PN0P_  (.D(_0089_),
    .Q(net103),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[181]$_DFFE_PN0P_  (.D(_0090_),
    .Q(net104),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[182]$_DFFE_PN0P_  (.D(_0091_),
    .Q(net105),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[183]$_DFFE_PN0P_  (.D(_0092_),
    .Q(net106),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[184]$_DFFE_PN0P_  (.D(_0093_),
    .Q(net107),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[185]$_DFFE_PN0P_  (.D(_0094_),
    .Q(net108),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[186]$_DFFE_PN0P_  (.D(_0095_),
    .Q(net109),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[187]$_DFFE_PN0P_  (.D(_0096_),
    .Q(net110),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[188]$_DFFE_PN0P_  (.D(_0097_),
    .Q(net111),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[189]$_DFFE_PN0P_  (.D(_0098_),
    .Q(net112),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[18]$_DFFE_PN0P_  (.D(_0099_),
    .Q(net113),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[190]$_DFFE_PN0P_  (.D(_0100_),
    .Q(net114),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[191]$_DFFE_PN0P_  (.D(_0101_),
    .Q(net115),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[192]$_DFFE_PN0P_  (.D(_0102_),
    .Q(net116),
    .RESET_B(net13),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[193]$_DFFE_PN0P_  (.D(_0103_),
    .Q(net117),
    .RESET_B(net13),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[194]$_DFFE_PN0P_  (.D(_0104_),
    .Q(net118),
    .RESET_B(net13),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[195]$_DFFE_PN0P_  (.D(_0105_),
    .Q(net119),
    .RESET_B(net13),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[196]$_DFFE_PN0P_  (.D(_0106_),
    .Q(net120),
    .RESET_B(net13),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[197]$_DFFE_PN0P_  (.D(_0107_),
    .Q(net121),
    .RESET_B(net13),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[198]$_DFFE_PN0P_  (.D(_0108_),
    .Q(net122),
    .RESET_B(net13),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[199]$_DFFE_PN0P_  (.D(_0109_),
    .Q(net123),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[19]$_DFFE_PN0P_  (.D(_0110_),
    .Q(net124),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[1]$_DFFE_PN0P_  (.D(_0111_),
    .Q(net125),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[200]$_DFFE_PN0P_  (.D(_0112_),
    .Q(net126),
    .RESET_B(net13),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[201]$_DFFE_PN0P_  (.D(_0113_),
    .Q(net127),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[202]$_DFFE_PN0P_  (.D(_0114_),
    .Q(net128),
    .RESET_B(net13),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[203]$_DFFE_PN0P_  (.D(_0115_),
    .Q(net129),
    .RESET_B(net13),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[204]$_DFFE_PN0P_  (.D(_0116_),
    .Q(net130),
    .RESET_B(net13),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[205]$_DFFE_PN0P_  (.D(_0117_),
    .Q(net131),
    .RESET_B(net13),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[206]$_DFFE_PN0P_  (.D(_0118_),
    .Q(net132),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[207]$_DFFE_PN0P_  (.D(_0119_),
    .Q(net133),
    .RESET_B(net13),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[208]$_DFFE_PN0P_  (.D(_0120_),
    .Q(net134),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[209]$_DFFE_PN0P_  (.D(_0121_),
    .Q(net135),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[20]$_DFFE_PN0P_  (.D(_0122_),
    .Q(net136),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[210]$_DFFE_PN0P_  (.D(_0123_),
    .Q(net137),
    .RESET_B(net13),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[211]$_DFFE_PN0P_  (.D(_0124_),
    .Q(net138),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[212]$_DFFE_PN0P_  (.D(_0125_),
    .Q(net139),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[213]$_DFFE_PN0P_  (.D(_0126_),
    .Q(net140),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[214]$_DFFE_PN0P_  (.D(_0127_),
    .Q(net141),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[215]$_DFFE_PN0P_  (.D(_0128_),
    .Q(net142),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[216]$_DFFE_PN0P_  (.D(_0129_),
    .Q(net143),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[217]$_DFFE_PN0P_  (.D(_0130_),
    .Q(net144),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[218]$_DFFE_PN0P_  (.D(_0131_),
    .Q(net145),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[219]$_DFFE_PN0P_  (.D(_0132_),
    .Q(net146),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[21]$_DFFE_PN0P_  (.D(_0133_),
    .Q(net147),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[220]$_DFFE_PN0P_  (.D(_0134_),
    .Q(net148),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[221]$_DFFE_PN0P_  (.D(_0135_),
    .Q(net149),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[222]$_DFFE_PN0P_  (.D(_0136_),
    .Q(net150),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[223]$_DFFE_PN0P_  (.D(_0137_),
    .Q(net151),
    .RESET_B(net13),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[224]$_DFFE_PN0P_  (.D(_0138_),
    .Q(net152),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[225]$_DFFE_PN0P_  (.D(_0139_),
    .Q(net153),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[226]$_DFFE_PN0P_  (.D(_0140_),
    .Q(net154),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[227]$_DFFE_PN0P_  (.D(_0141_),
    .Q(net155),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[228]$_DFFE_PN0P_  (.D(_0142_),
    .Q(net156),
    .RESET_B(net13),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[229]$_DFFE_PN0P_  (.D(_0143_),
    .Q(net157),
    .RESET_B(net13),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[22]$_DFFE_PN0P_  (.D(_0144_),
    .Q(net158),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[230]$_DFFE_PN0P_  (.D(_0145_),
    .Q(net159),
    .RESET_B(net13),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[231]$_DFFE_PN0P_  (.D(_0146_),
    .Q(net160),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[232]$_DFFE_PN0P_  (.D(_0147_),
    .Q(net161),
    .RESET_B(net13),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[233]$_DFFE_PN0P_  (.D(_0148_),
    .Q(net162),
    .RESET_B(net13),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[234]$_DFFE_PN0P_  (.D(_0149_),
    .Q(net163),
    .RESET_B(net13),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[235]$_DFFE_PN0P_  (.D(_0150_),
    .Q(net164),
    .RESET_B(net13),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[236]$_DFFE_PN0P_  (.D(_0151_),
    .Q(net165),
    .RESET_B(net13),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[237]$_DFFE_PN0P_  (.D(_0152_),
    .Q(net166),
    .RESET_B(net13),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[238]$_DFFE_PN0P_  (.D(_0153_),
    .Q(net167),
    .RESET_B(net13),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[239]$_DFFE_PN0P_  (.D(_0154_),
    .Q(net168),
    .RESET_B(net13),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[23]$_DFFE_PN0P_  (.D(_0155_),
    .Q(net169),
    .RESET_B(net13),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[240]$_DFFE_PN0P_  (.D(_0156_),
    .Q(net170),
    .RESET_B(net13),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[241]$_DFFE_PN0P_  (.D(_0157_),
    .Q(net171),
    .RESET_B(net13),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[242]$_DFFE_PN0P_  (.D(_0158_),
    .Q(net172),
    .RESET_B(net13),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[243]$_DFFE_PN0P_  (.D(_0159_),
    .Q(net173),
    .RESET_B(net13),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[244]$_DFFE_PN0P_  (.D(_0160_),
    .Q(net174),
    .RESET_B(net13),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[245]$_DFFE_PN0P_  (.D(_0161_),
    .Q(net175),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[246]$_DFFE_PN0P_  (.D(_0162_),
    .Q(net176),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[247]$_DFFE_PN0P_  (.D(_0163_),
    .Q(net177),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[248]$_DFFE_PN0P_  (.D(_0164_),
    .Q(net178),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[249]$_DFFE_PN0P_  (.D(_0165_),
    .Q(net179),
    .RESET_B(net13),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[24]$_DFFE_PN0P_  (.D(_0166_),
    .Q(net180),
    .RESET_B(net13),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[250]$_DFFE_PN0P_  (.D(_0167_),
    .Q(net181),
    .RESET_B(net13),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[251]$_DFFE_PN0P_  (.D(_0168_),
    .Q(net182),
    .RESET_B(net13),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[252]$_DFFE_PN0P_  (.D(_0169_),
    .Q(net183),
    .RESET_B(net13),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[253]$_DFFE_PN0P_  (.D(_0170_),
    .Q(net184),
    .RESET_B(net13),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[254]$_DFFE_PN0P_  (.D(_0171_),
    .Q(net185),
    .RESET_B(net13),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[255]$_DFFE_PN0P_  (.D(_0172_),
    .Q(net186),
    .RESET_B(net13),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[25]$_DFFE_PN0P_  (.D(_0173_),
    .Q(net187),
    .RESET_B(net13),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[26]$_DFFE_PN0P_  (.D(_0174_),
    .Q(net188),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[27]$_DFFE_PN0P_  (.D(_0175_),
    .Q(net189),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[28]$_DFFE_PN0P_  (.D(_0176_),
    .Q(net190),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[29]$_DFFE_PN0P_  (.D(_0177_),
    .Q(net191),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[2]$_DFFE_PN0P_  (.D(_0178_),
    .Q(net192),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[30]$_DFFE_PN0P_  (.D(_0179_),
    .Q(net193),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[31]$_DFFE_PN0P_  (.D(_0180_),
    .Q(net194),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[32]$_DFFE_PN0P_  (.D(_0181_),
    .Q(net195),
    .RESET_B(net13),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[33]$_DFFE_PN0P_  (.D(_0182_),
    .Q(net196),
    .RESET_B(net13),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[34]$_DFFE_PN0P_  (.D(_0183_),
    .Q(net197),
    .RESET_B(net13),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[35]$_DFFE_PN0P_  (.D(_0184_),
    .Q(net198),
    .RESET_B(net13),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[36]$_DFFE_PN0P_  (.D(_0185_),
    .Q(net199),
    .RESET_B(net13),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[37]$_DFFE_PN0P_  (.D(_0186_),
    .Q(net200),
    .RESET_B(net13),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[38]$_DFFE_PN0P_  (.D(_0187_),
    .Q(net201),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[39]$_DFFE_PN0P_  (.D(_0188_),
    .Q(net202),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[3]$_DFFE_PN0P_  (.D(_0189_),
    .Q(net203),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[40]$_DFFE_PN0P_  (.D(_0190_),
    .Q(net204),
    .RESET_B(net13),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[41]$_DFFE_PN0P_  (.D(_0191_),
    .Q(net205),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[42]$_DFFE_PN0P_  (.D(_0192_),
    .Q(net206),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[43]$_DFFE_PN0P_  (.D(_0193_),
    .Q(net207),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[44]$_DFFE_PN0P_  (.D(_0194_),
    .Q(net208),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[45]$_DFFE_PN0P_  (.D(_0195_),
    .Q(net209),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[46]$_DFFE_PN0P_  (.D(_0196_),
    .Q(net210),
    .RESET_B(net13),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[47]$_DFFE_PN0P_  (.D(_0197_),
    .Q(net211),
    .RESET_B(net13),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[48]$_DFFE_PN0P_  (.D(_0198_),
    .Q(net212),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[49]$_DFFE_PN0P_  (.D(_0199_),
    .Q(net213),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[4]$_DFFE_PN0P_  (.D(_0200_),
    .Q(net214),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[50]$_DFFE_PN0P_  (.D(_0201_),
    .Q(net215),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[51]$_DFFE_PN0P_  (.D(_0202_),
    .Q(net216),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[52]$_DFFE_PN0P_  (.D(_0203_),
    .Q(net217),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[53]$_DFFE_PN0P_  (.D(_0204_),
    .Q(net218),
    .RESET_B(net13),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[54]$_DFFE_PN0P_  (.D(_0205_),
    .Q(net219),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[55]$_DFFE_PN0P_  (.D(_0206_),
    .Q(net220),
    .RESET_B(net13),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[56]$_DFFE_PN0P_  (.D(_0207_),
    .Q(net221),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[57]$_DFFE_PN0P_  (.D(_0208_),
    .Q(net222),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[58]$_DFFE_PN0P_  (.D(_0209_),
    .Q(net223),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[59]$_DFFE_PN0P_  (.D(_0210_),
    .Q(net224),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[5]$_DFFE_PN0P_  (.D(_0211_),
    .Q(net225),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[60]$_DFFE_PN0P_  (.D(_0212_),
    .Q(net226),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[61]$_DFFE_PN0P_  (.D(_0213_),
    .Q(net227),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[62]$_DFFE_PN0P_  (.D(_0214_),
    .Q(net228),
    .RESET_B(net13),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[63]$_DFFE_PN0P_  (.D(_0215_),
    .Q(net229),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[64]$_DFFE_PN0P_  (.D(_0216_),
    .Q(net230),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[65]$_DFFE_PN0P_  (.D(_0217_),
    .Q(net231),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[66]$_DFFE_PN0P_  (.D(_0218_),
    .Q(net232),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[67]$_DFFE_PN0P_  (.D(_0219_),
    .Q(net233),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[68]$_DFFE_PN0P_  (.D(_0220_),
    .Q(net234),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[69]$_DFFE_PN0P_  (.D(_0221_),
    .Q(net235),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[6]$_DFFE_PN0P_  (.D(_0222_),
    .Q(net236),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[70]$_DFFE_PN0P_  (.D(_0223_),
    .Q(net237),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[71]$_DFFE_PN0P_  (.D(_0224_),
    .Q(net238),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[72]$_DFFE_PN0P_  (.D(_0225_),
    .Q(net239),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[73]$_DFFE_PN0P_  (.D(_0226_),
    .Q(net240),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[74]$_DFFE_PN0P_  (.D(_0227_),
    .Q(net241),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[75]$_DFFE_PN0P_  (.D(_0228_),
    .Q(net242),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[76]$_DFFE_PN0P_  (.D(_0229_),
    .Q(net243),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[77]$_DFFE_PN0P_  (.D(_0230_),
    .Q(net244),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[78]$_DFFE_PN0P_  (.D(_0231_),
    .Q(net245),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[79]$_DFFE_PN0P_  (.D(_0232_),
    .Q(net246),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[7]$_DFFE_PN0P_  (.D(_0233_),
    .Q(net247),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[80]$_DFFE_PN0P_  (.D(_0234_),
    .Q(net248),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[81]$_DFFE_PN0P_  (.D(_0235_),
    .Q(net249),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[82]$_DFFE_PN0P_  (.D(_0236_),
    .Q(net250),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[83]$_DFFE_PN0P_  (.D(_0237_),
    .Q(net251),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[84]$_DFFE_PN0P_  (.D(_0238_),
    .Q(net252),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[85]$_DFFE_PN0P_  (.D(_0239_),
    .Q(net253),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[86]$_DFFE_PN0P_  (.D(_0240_),
    .Q(net254),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[87]$_DFFE_PN0P_  (.D(_0241_),
    .Q(net255),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[88]$_DFFE_PN0P_  (.D(_0242_),
    .Q(net256),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[89]$_DFFE_PN0P_  (.D(_0243_),
    .Q(net257),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[8]$_DFFE_PN0P_  (.D(_0244_),
    .Q(net258),
    .RESET_B(net13),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[90]$_DFFE_PN0P_  (.D(_0245_),
    .Q(net259),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[91]$_DFFE_PN0P_  (.D(_0246_),
    .Q(net260),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[92]$_DFFE_PN0P_  (.D(_0247_),
    .Q(net261),
    .RESET_B(net13),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[93]$_DFFE_PN0P_  (.D(_0248_),
    .Q(net262),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[94]$_DFFE_PN0P_  (.D(_0249_),
    .Q(net263),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[95]$_DFFE_PN0P_  (.D(_0250_),
    .Q(net264),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[96]$_DFFE_PN0P_  (.D(_0251_),
    .Q(net265),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_2 \counters[97]$_DFFE_PN0P_  (.D(_0252_),
    .Q(net266),
    .RESET_B(net13),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[98]$_DFFE_PN0P_  (.D(_0253_),
    .Q(net267),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \counters[99]$_DFFE_PN0P_  (.D(_0254_),
    .Q(net268),
    .RESET_B(net13),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \counters[9]$_DFFE_PN0P_  (.D(_0255_),
    .Q(net269),
    .RESET_B(net13),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \prev_event_inc[0]$_DFFE_PN0N_  (.D(_0256_),
    .Q(\prev_event_inc[0] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \prev_event_inc[1]$_DFFE_PN0N_  (.D(_0257_),
    .Q(\prev_event_inc[1] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \prev_event_inc[2]$_DFFE_PN0N_  (.D(_0258_),
    .Q(\prev_event_inc[2] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \prev_event_inc[3]$_DFFE_PN0N_  (.D(_0259_),
    .Q(\prev_event_inc[3] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \prev_event_inc[4]$_DFFE_PN0N_  (.D(_0260_),
    .Q(\prev_event_inc[4] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \prev_event_inc[5]$_DFFE_PN0N_  (.D(_0261_),
    .Q(\prev_event_inc[5] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \prev_event_inc[6]$_DFFE_PN0N_  (.D(_0262_),
    .Q(\prev_event_inc[6] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \prev_event_inc[7]$_DFFE_PN0N_  (.D(_0263_),
    .Q(\prev_event_inc[7] ),
    .RESET_B(net13),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_383 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(counter_sel[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(counter_sel[6]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(counter_sel[7]),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input4 (.A(enable),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(net304),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(net302),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(net307),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(net306),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(net303),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(net305),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(net309),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(net308),
    .X(net12));
 sky130_fd_sc_hd__buf_16 input13 (.A(rst_n),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .X(all_counts[0]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(all_counts[100]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(all_counts[101]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(all_counts[102]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(all_counts[103]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(all_counts[104]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(all_counts[105]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(all_counts[106]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(all_counts[107]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(all_counts[108]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(all_counts[109]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(all_counts[10]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(all_counts[110]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(all_counts[111]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(all_counts[112]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(all_counts[113]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .X(all_counts[114]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .X(all_counts[115]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net32),
    .X(all_counts[116]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .X(all_counts[117]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net34),
    .X(all_counts[118]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net35),
    .X(all_counts[119]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(all_counts[11]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net37),
    .X(all_counts[120]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net38),
    .X(all_counts[121]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net39),
    .X(all_counts[122]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net40),
    .X(all_counts[123]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net41),
    .X(all_counts[124]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net42),
    .X(all_counts[125]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net43),
    .X(all_counts[126]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net44),
    .X(all_counts[127]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net45),
    .X(all_counts[128]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net46),
    .X(all_counts[129]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net47),
    .X(all_counts[12]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net48),
    .X(all_counts[130]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net49),
    .X(all_counts[131]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net50),
    .X(all_counts[132]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net51),
    .X(all_counts[133]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net52),
    .X(all_counts[134]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(all_counts[135]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(all_counts[136]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(all_counts[137]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(all_counts[138]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(all_counts[139]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(all_counts[13]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(all_counts[140]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(all_counts[141]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(all_counts[142]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(all_counts[143]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(all_counts[144]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .X(all_counts[145]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .X(all_counts[146]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(all_counts[147]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(all_counts[148]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(all_counts[149]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(all_counts[14]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(all_counts[150]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(all_counts[151]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(all_counts[152]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(all_counts[153]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(all_counts[154]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(all_counts[155]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(all_counts[156]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(all_counts[157]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(all_counts[158]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(all_counts[159]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(all_counts[15]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(all_counts[160]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(all_counts[161]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(all_counts[162]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(all_counts[163]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .X(all_counts[164]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .X(all_counts[165]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(all_counts[166]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(all_counts[167]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(all_counts[168]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .X(all_counts[169]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .X(all_counts[16]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(all_counts[170]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .X(all_counts[171]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .X(all_counts[172]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(all_counts[173]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .X(all_counts[174]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .X(all_counts[175]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .X(all_counts[176]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net99),
    .X(all_counts[177]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net100),
    .X(all_counts[178]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net101),
    .X(all_counts[179]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net102),
    .X(all_counts[17]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net103),
    .X(all_counts[180]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net104),
    .X(all_counts[181]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net105),
    .X(all_counts[182]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net106),
    .X(all_counts[183]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net107),
    .X(all_counts[184]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net108),
    .X(all_counts[185]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net109),
    .X(all_counts[186]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net110),
    .X(all_counts[187]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net111),
    .X(all_counts[188]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net112),
    .X(all_counts[189]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net113),
    .X(all_counts[18]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net114),
    .X(all_counts[190]));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net115),
    .X(all_counts[191]));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net116),
    .X(all_counts[192]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net117),
    .X(all_counts[193]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net118),
    .X(all_counts[194]));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net119),
    .X(all_counts[195]));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net120),
    .X(all_counts[196]));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net121),
    .X(all_counts[197]));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net122),
    .X(all_counts[198]));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net123),
    .X(all_counts[199]));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net124),
    .X(all_counts[19]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net125),
    .X(all_counts[1]));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net126),
    .X(all_counts[200]));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net127),
    .X(all_counts[201]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net128),
    .X(all_counts[202]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net129),
    .X(all_counts[203]));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net130),
    .X(all_counts[204]));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net131),
    .X(all_counts[205]));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net132),
    .X(all_counts[206]));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net133),
    .X(all_counts[207]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net134),
    .X(all_counts[208]));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net135),
    .X(all_counts[209]));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net136),
    .X(all_counts[20]));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net137),
    .X(all_counts[210]));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net138),
    .X(all_counts[211]));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net139),
    .X(all_counts[212]));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net140),
    .X(all_counts[213]));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net141),
    .X(all_counts[214]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net142),
    .X(all_counts[215]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net143),
    .X(all_counts[216]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net144),
    .X(all_counts[217]));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net145),
    .X(all_counts[218]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net146),
    .X(all_counts[219]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net147),
    .X(all_counts[21]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net148),
    .X(all_counts[220]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net149),
    .X(all_counts[221]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net150),
    .X(all_counts[222]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net151),
    .X(all_counts[223]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net152),
    .X(all_counts[224]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net153),
    .X(all_counts[225]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net154),
    .X(all_counts[226]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net155),
    .X(all_counts[227]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net156),
    .X(all_counts[228]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net157),
    .X(all_counts[229]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net158),
    .X(all_counts[22]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net159),
    .X(all_counts[230]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net160),
    .X(all_counts[231]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net161),
    .X(all_counts[232]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net162),
    .X(all_counts[233]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net163),
    .X(all_counts[234]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net164),
    .X(all_counts[235]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net165),
    .X(all_counts[236]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net166),
    .X(all_counts[237]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net167),
    .X(all_counts[238]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net168),
    .X(all_counts[239]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net169),
    .X(all_counts[23]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net170),
    .X(all_counts[240]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net171),
    .X(all_counts[241]));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net172),
    .X(all_counts[242]));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net173),
    .X(all_counts[243]));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net174),
    .X(all_counts[244]));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net175),
    .X(all_counts[245]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net176),
    .X(all_counts[246]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net177),
    .X(all_counts[247]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net178),
    .X(all_counts[248]));
 sky130_fd_sc_hd__clkbuf_1 output179 (.A(net179),
    .X(all_counts[249]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net180),
    .X(all_counts[24]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net181),
    .X(all_counts[250]));
 sky130_fd_sc_hd__clkbuf_1 output182 (.A(net182),
    .X(all_counts[251]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net183),
    .X(all_counts[252]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net184),
    .X(all_counts[253]));
 sky130_fd_sc_hd__clkbuf_1 output185 (.A(net185),
    .X(all_counts[254]));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net186),
    .X(all_counts[255]));
 sky130_fd_sc_hd__clkbuf_1 output187 (.A(net187),
    .X(all_counts[25]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net188),
    .X(all_counts[26]));
 sky130_fd_sc_hd__clkbuf_1 output189 (.A(net189),
    .X(all_counts[27]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net190),
    .X(all_counts[28]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net191),
    .X(all_counts[29]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(net192),
    .X(all_counts[2]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net193),
    .X(all_counts[30]));
 sky130_fd_sc_hd__clkbuf_1 output194 (.A(net194),
    .X(all_counts[31]));
 sky130_fd_sc_hd__clkbuf_1 output195 (.A(net195),
    .X(all_counts[32]));
 sky130_fd_sc_hd__clkbuf_1 output196 (.A(net196),
    .X(all_counts[33]));
 sky130_fd_sc_hd__clkbuf_1 output197 (.A(net197),
    .X(all_counts[34]));
 sky130_fd_sc_hd__clkbuf_1 output198 (.A(net198),
    .X(all_counts[35]));
 sky130_fd_sc_hd__clkbuf_1 output199 (.A(net199),
    .X(all_counts[36]));
 sky130_fd_sc_hd__clkbuf_1 output200 (.A(net200),
    .X(all_counts[37]));
 sky130_fd_sc_hd__clkbuf_1 output201 (.A(net201),
    .X(all_counts[38]));
 sky130_fd_sc_hd__clkbuf_1 output202 (.A(net202),
    .X(all_counts[39]));
 sky130_fd_sc_hd__clkbuf_1 output203 (.A(net203),
    .X(all_counts[3]));
 sky130_fd_sc_hd__clkbuf_1 output204 (.A(net204),
    .X(all_counts[40]));
 sky130_fd_sc_hd__clkbuf_1 output205 (.A(net205),
    .X(all_counts[41]));
 sky130_fd_sc_hd__clkbuf_1 output206 (.A(net206),
    .X(all_counts[42]));
 sky130_fd_sc_hd__clkbuf_1 output207 (.A(net207),
    .X(all_counts[43]));
 sky130_fd_sc_hd__clkbuf_1 output208 (.A(net208),
    .X(all_counts[44]));
 sky130_fd_sc_hd__clkbuf_1 output209 (.A(net209),
    .X(all_counts[45]));
 sky130_fd_sc_hd__clkbuf_1 output210 (.A(net210),
    .X(all_counts[46]));
 sky130_fd_sc_hd__clkbuf_1 output211 (.A(net211),
    .X(all_counts[47]));
 sky130_fd_sc_hd__clkbuf_1 output212 (.A(net212),
    .X(all_counts[48]));
 sky130_fd_sc_hd__clkbuf_1 output213 (.A(net213),
    .X(all_counts[49]));
 sky130_fd_sc_hd__clkbuf_1 output214 (.A(net214),
    .X(all_counts[4]));
 sky130_fd_sc_hd__clkbuf_1 output215 (.A(net215),
    .X(all_counts[50]));
 sky130_fd_sc_hd__clkbuf_1 output216 (.A(net216),
    .X(all_counts[51]));
 sky130_fd_sc_hd__clkbuf_1 output217 (.A(net217),
    .X(all_counts[52]));
 sky130_fd_sc_hd__clkbuf_1 output218 (.A(net218),
    .X(all_counts[53]));
 sky130_fd_sc_hd__clkbuf_1 output219 (.A(net219),
    .X(all_counts[54]));
 sky130_fd_sc_hd__clkbuf_1 output220 (.A(net220),
    .X(all_counts[55]));
 sky130_fd_sc_hd__clkbuf_1 output221 (.A(net221),
    .X(all_counts[56]));
 sky130_fd_sc_hd__clkbuf_1 output222 (.A(net222),
    .X(all_counts[57]));
 sky130_fd_sc_hd__clkbuf_1 output223 (.A(net223),
    .X(all_counts[58]));
 sky130_fd_sc_hd__clkbuf_1 output224 (.A(net224),
    .X(all_counts[59]));
 sky130_fd_sc_hd__clkbuf_1 output225 (.A(net225),
    .X(all_counts[5]));
 sky130_fd_sc_hd__clkbuf_1 output226 (.A(net226),
    .X(all_counts[60]));
 sky130_fd_sc_hd__clkbuf_1 output227 (.A(net227),
    .X(all_counts[61]));
 sky130_fd_sc_hd__clkbuf_1 output228 (.A(net228),
    .X(all_counts[62]));
 sky130_fd_sc_hd__clkbuf_1 output229 (.A(net229),
    .X(all_counts[63]));
 sky130_fd_sc_hd__clkbuf_1 output230 (.A(net230),
    .X(all_counts[64]));
 sky130_fd_sc_hd__clkbuf_1 output231 (.A(net231),
    .X(all_counts[65]));
 sky130_fd_sc_hd__clkbuf_1 output232 (.A(net232),
    .X(all_counts[66]));
 sky130_fd_sc_hd__clkbuf_1 output233 (.A(net233),
    .X(all_counts[67]));
 sky130_fd_sc_hd__clkbuf_1 output234 (.A(net234),
    .X(all_counts[68]));
 sky130_fd_sc_hd__clkbuf_1 output235 (.A(net235),
    .X(all_counts[69]));
 sky130_fd_sc_hd__clkbuf_1 output236 (.A(net236),
    .X(all_counts[6]));
 sky130_fd_sc_hd__clkbuf_1 output237 (.A(net237),
    .X(all_counts[70]));
 sky130_fd_sc_hd__clkbuf_1 output238 (.A(net238),
    .X(all_counts[71]));
 sky130_fd_sc_hd__clkbuf_1 output239 (.A(net239),
    .X(all_counts[72]));
 sky130_fd_sc_hd__clkbuf_1 output240 (.A(net240),
    .X(all_counts[73]));
 sky130_fd_sc_hd__clkbuf_1 output241 (.A(net241),
    .X(all_counts[74]));
 sky130_fd_sc_hd__clkbuf_1 output242 (.A(net242),
    .X(all_counts[75]));
 sky130_fd_sc_hd__clkbuf_1 output243 (.A(net243),
    .X(all_counts[76]));
 sky130_fd_sc_hd__clkbuf_1 output244 (.A(net244),
    .X(all_counts[77]));
 sky130_fd_sc_hd__clkbuf_1 output245 (.A(net245),
    .X(all_counts[78]));
 sky130_fd_sc_hd__clkbuf_1 output246 (.A(net246),
    .X(all_counts[79]));
 sky130_fd_sc_hd__clkbuf_1 output247 (.A(net247),
    .X(all_counts[7]));
 sky130_fd_sc_hd__clkbuf_1 output248 (.A(net248),
    .X(all_counts[80]));
 sky130_fd_sc_hd__clkbuf_1 output249 (.A(net249),
    .X(all_counts[81]));
 sky130_fd_sc_hd__clkbuf_1 output250 (.A(net250),
    .X(all_counts[82]));
 sky130_fd_sc_hd__clkbuf_1 output251 (.A(net251),
    .X(all_counts[83]));
 sky130_fd_sc_hd__clkbuf_1 output252 (.A(net252),
    .X(all_counts[84]));
 sky130_fd_sc_hd__clkbuf_1 output253 (.A(net253),
    .X(all_counts[85]));
 sky130_fd_sc_hd__clkbuf_1 output254 (.A(net254),
    .X(all_counts[86]));
 sky130_fd_sc_hd__clkbuf_1 output255 (.A(net255),
    .X(all_counts[87]));
 sky130_fd_sc_hd__clkbuf_1 output256 (.A(net256),
    .X(all_counts[88]));
 sky130_fd_sc_hd__clkbuf_1 output257 (.A(net257),
    .X(all_counts[89]));
 sky130_fd_sc_hd__clkbuf_1 output258 (.A(net258),
    .X(all_counts[8]));
 sky130_fd_sc_hd__clkbuf_1 output259 (.A(net259),
    .X(all_counts[90]));
 sky130_fd_sc_hd__clkbuf_1 output260 (.A(net260),
    .X(all_counts[91]));
 sky130_fd_sc_hd__clkbuf_1 output261 (.A(net261),
    .X(all_counts[92]));
 sky130_fd_sc_hd__clkbuf_1 output262 (.A(net262),
    .X(all_counts[93]));
 sky130_fd_sc_hd__clkbuf_1 output263 (.A(net263),
    .X(all_counts[94]));
 sky130_fd_sc_hd__clkbuf_1 output264 (.A(net264),
    .X(all_counts[95]));
 sky130_fd_sc_hd__clkbuf_1 output265 (.A(net265),
    .X(all_counts[96]));
 sky130_fd_sc_hd__clkbuf_1 output266 (.A(net266),
    .X(all_counts[97]));
 sky130_fd_sc_hd__clkbuf_1 output267 (.A(net267),
    .X(all_counts[98]));
 sky130_fd_sc_hd__clkbuf_1 output268 (.A(net268),
    .X(all_counts[99]));
 sky130_fd_sc_hd__clkbuf_1 output269 (.A(net269),
    .X(all_counts[9]));
 sky130_fd_sc_hd__clkbuf_1 output270 (.A(net270),
    .X(count_value[0]));
 sky130_fd_sc_hd__clkbuf_1 output271 (.A(net271),
    .X(count_value[10]));
 sky130_fd_sc_hd__clkbuf_1 output272 (.A(net272),
    .X(count_value[11]));
 sky130_fd_sc_hd__clkbuf_1 output273 (.A(net273),
    .X(count_value[12]));
 sky130_fd_sc_hd__clkbuf_1 output274 (.A(net274),
    .X(count_value[13]));
 sky130_fd_sc_hd__clkbuf_1 output275 (.A(net275),
    .X(count_value[14]));
 sky130_fd_sc_hd__clkbuf_1 output276 (.A(net276),
    .X(count_value[15]));
 sky130_fd_sc_hd__clkbuf_1 output277 (.A(net277),
    .X(count_value[16]));
 sky130_fd_sc_hd__clkbuf_1 output278 (.A(net278),
    .X(count_value[17]));
 sky130_fd_sc_hd__clkbuf_1 output279 (.A(net279),
    .X(count_value[18]));
 sky130_fd_sc_hd__clkbuf_1 output280 (.A(net280),
    .X(count_value[19]));
 sky130_fd_sc_hd__clkbuf_1 output281 (.A(net281),
    .X(count_value[1]));
 sky130_fd_sc_hd__clkbuf_1 output282 (.A(net282),
    .X(count_value[20]));
 sky130_fd_sc_hd__clkbuf_1 output283 (.A(net283),
    .X(count_value[21]));
 sky130_fd_sc_hd__clkbuf_1 output284 (.A(net284),
    .X(count_value[22]));
 sky130_fd_sc_hd__clkbuf_1 output285 (.A(net285),
    .X(count_value[23]));
 sky130_fd_sc_hd__clkbuf_1 output286 (.A(net286),
    .X(count_value[24]));
 sky130_fd_sc_hd__clkbuf_1 output287 (.A(net287),
    .X(count_value[25]));
 sky130_fd_sc_hd__clkbuf_1 output288 (.A(net288),
    .X(count_value[26]));
 sky130_fd_sc_hd__clkbuf_1 output289 (.A(net289),
    .X(count_value[27]));
 sky130_fd_sc_hd__clkbuf_1 output290 (.A(net290),
    .X(count_value[28]));
 sky130_fd_sc_hd__clkbuf_1 output291 (.A(net291),
    .X(count_value[29]));
 sky130_fd_sc_hd__clkbuf_1 output292 (.A(net292),
    .X(count_value[2]));
 sky130_fd_sc_hd__clkbuf_1 output293 (.A(net293),
    .X(count_value[30]));
 sky130_fd_sc_hd__clkbuf_1 output294 (.A(net294),
    .X(count_value[31]));
 sky130_fd_sc_hd__clkbuf_1 output295 (.A(net295),
    .X(count_value[3]));
 sky130_fd_sc_hd__clkbuf_1 output296 (.A(net296),
    .X(count_value[4]));
 sky130_fd_sc_hd__clkbuf_1 output297 (.A(net297),
    .X(count_value[5]));
 sky130_fd_sc_hd__clkbuf_1 output298 (.A(net298),
    .X(count_value[6]));
 sky130_fd_sc_hd__clkbuf_1 output299 (.A(net299),
    .X(count_value[7]));
 sky130_fd_sc_hd__clkbuf_1 output300 (.A(net300),
    .X(count_value[8]));
 sky130_fd_sc_hd__clkbuf_1 output301 (.A(net301),
    .X(count_value[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload1 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinv_2 clkload5 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload6 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload7 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkinv_2 clkload8 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload9 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload11 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload12 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload13 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__inv_8 clkload14 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload15 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload16 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload17 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload18 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload19 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__bufinv_16 clkload20 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload21 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_2 clkload22 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload23 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload24 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload25 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinv_2 clkload26 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(event_inc[1]),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(event_inc[4]),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(event_inc[0]),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(event_inc[5]),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(event_inc[3]),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(event_inc[2]),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(event_inc[7]),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(event_inc[6]),
    .X(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net191));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_7 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_371 ();
endmodule
