module parameterized_loadable_counter (clk,
    enable,
    load,
    rst_n,
    count,
    data_in);
 input clk;
 input enable;
 input load;
 input rst_n;
 output [7:0] count;
 input [7:0] data_in;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net20;

 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _34_ (.A1(net10),
    .A2(net12),
    .Z(_08_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _35_ (.I(net11),
    .ZN(_09_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _36_ (.I0(net2),
    .I1(_08_),
    .S(_09_),
    .Z(_00_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _37_ (.I0(net13),
    .I1(_33_),
    .S(net10),
    .Z(_10_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _38_ (.I0(net3),
    .I1(_10_),
    .S(_09_),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _39_ (.A1(net10),
    .A2(_32_),
    .ZN(_11_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _40_ (.A1(net14),
    .A2(_11_),
    .ZN(_12_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _41_ (.I0(net4),
    .I1(_12_),
    .S(_09_),
    .Z(_02_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _42_ (.A1(net10),
    .A2(net12),
    .A3(net14),
    .A4(net13),
    .Z(_13_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _43_ (.A1(net15),
    .A2(_13_),
    .Z(_14_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _44_ (.I0(net5),
    .I1(_14_),
    .S(_09_),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _45_ (.A1(net10),
    .A2(_32_),
    .A3(net14),
    .A4(net15),
    .Z(_15_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _46_ (.A1(net16),
    .A2(_15_),
    .Z(_16_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _47_ (.I0(net6),
    .I1(_16_),
    .S(_09_),
    .Z(_04_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _48_ (.A1(net11),
    .A2(net7),
    .Z(_17_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _49_ (.A1(net15),
    .A2(net16),
    .Z(_18_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _50_ (.I(net17),
    .ZN(_19_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _51_ (.A1(_13_),
    .A2(_18_),
    .B(net11),
    .C(_19_),
    .ZN(_20_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _52_ (.A1(_09_),
    .A2(_19_),
    .A3(_13_),
    .A4(_18_),
    .Z(_21_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _53_ (.A1(_17_),
    .A2(_20_),
    .A3(_21_),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _54_ (.A1(net11),
    .A2(net8),
    .ZN(_22_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _55_ (.A1(net10),
    .A2(_32_),
    .A3(net14),
    .ZN(_23_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _56_ (.A1(net15),
    .A2(net16),
    .A3(net17),
    .ZN(_24_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _57_ (.A1(_23_),
    .A2(_24_),
    .B(_09_),
    .C(net18),
    .ZN(_25_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _58_ (.A1(net11),
    .A2(net18),
    .A3(_23_),
    .A4(_24_),
    .Z(_26_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _59_ (.A1(_22_),
    .A2(_25_),
    .A3(_26_),
    .ZN(_06_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _60_ (.A1(net15),
    .A2(net16),
    .A3(net17),
    .A4(net18),
    .Z(_27_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _61_ (.I(net19),
    .ZN(_28_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _62_ (.A1(_13_),
    .A2(_27_),
    .B(net11),
    .C(_28_),
    .ZN(_29_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _63_ (.A1(_09_),
    .A2(_28_),
    .A3(_13_),
    .A4(_27_),
    .Z(_30_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _64_ (.A1(net11),
    .A2(net9),
    .Z(_31_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _65_ (.A1(_29_),
    .A2(_30_),
    .A3(_31_),
    .Z(_07_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _66_ (.A(net12),
    .B(net13),
    .CO(_32_),
    .S(_33_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[0]$_DFFE_PN0P_  (.D(_00_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net12));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[1]$_DFFE_PN0P_  (.D(_01_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[2]$_DFFE_PN0P_  (.D(_02_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[3]$_DFFE_PN0P_  (.D(_03_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[4]$_DFFE_PN0P_  (.D(_04_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[5]$_DFFE_PN0P_  (.D(_05_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[6]$_DFFE_PN0P_  (.D(_06_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[7]$_DFFE_PN0P_  (.D(_07_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 hold1 (.I(net20),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_67 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(data_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(data_in[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(data_in[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(data_in[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(data_in[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(data_in[5]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(data_in[6]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(data_in[7]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input9 (.I(enable),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input10 (.I(load),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output11 (.I(net12),
    .Z(count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(count[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(count[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(count[7]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_244 ();
endmodule
