module final_spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire \bit_counter[0] ;
 wire \bit_counter[1] ;
 wire \bit_counter[2] ;
 wire \bit_counter[3] ;
 wire \miso_capture[0] ;
 wire \miso_capture[1] ;
 wire \miso_capture[2] ;
 wire \miso_capture[3] ;
 wire \miso_capture[4] ;
 wire \miso_capture[5] ;
 wire \miso_capture[6] ;
 wire \miso_capture[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \tx_shift[0] ;
 wire \tx_shift[1] ;
 wire \tx_shift[2] ;
 wire \tx_shift[3] ;
 wire \tx_shift[4] ;
 wire \tx_shift[5] ;
 wire \tx_shift[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net26;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _131_ (.I(\bit_counter[2] ),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _132_ (.I(_126_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _133_ (.A1(\bit_counter[3] ),
    .A2(_108_),
    .A3(_109_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _134_ (.I(_113_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _135_ (.I(\state[0] ),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _136_ (.A1(\state[1] ),
    .A2(_110_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _137_ (.I(_111_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _138_ (.I(\bit_counter[3] ),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _139_ (.A1(\bit_counter[2] ),
    .A2(\bit_counter[1] ),
    .A3(\bit_counter[0] ),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _140_ (.A1(\bit_counter[3] ),
    .A2(_128_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _141_ (.A1(net22),
    .A2(\bit_counter[3] ),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _142_ (.I(\state[1] ),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _143_ (.A1(_110_),
    .A2(_034_),
    .B(_035_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _144_ (.I(_036_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _145_ (.A1(_035_),
    .A2(\state[0] ),
    .A3(_034_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _146_ (.I(\bit_counter[0] ),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _147_ (.I0(_037_),
    .I1(_038_),
    .S(_039_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _148_ (.A1(\bit_counter[1] ),
    .A2(_037_),
    .B1(_038_),
    .B2(_127_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _149_ (.I(_040_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _150_ (.A1(_109_),
    .A2(_038_),
    .B(_037_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _151_ (.A1(_108_),
    .A2(_126_),
    .A3(_038_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _152_ (.A1(_108_),
    .A2(_041_),
    .B(_042_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _153_ (.I(_130_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _154_ (.A1(\state[1] ),
    .A2(net22),
    .A3(_043_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _155_ (.A1(_035_),
    .A2(_110_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _156_ (.A1(_112_),
    .A2(_044_),
    .B(_045_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _157_ (.I(_127_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _158_ (.A1(_115_),
    .A2(_046_),
    .A3(_130_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _159_ (.A1(\bit_counter[2] ),
    .A2(_126_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _160_ (.A1(_121_),
    .A2(_118_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _161_ (.A1(_039_),
    .A2(_048_),
    .A3(_049_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _162_ (.A1(_124_),
    .A2(_129_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _163_ (.A1(_115_),
    .A2(_125_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _164_ (.A1(_124_),
    .A2(_129_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _165_ (.A1(_115_),
    .A2(_125_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _166_ (.A1(_051_),
    .A2(_052_),
    .B1(_053_),
    .B2(_054_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _167_ (.A1(_047_),
    .A2(_050_),
    .A3(_055_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _168_ (.A1(\miso_capture[0] ),
    .A2(_038_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _169_ (.A1(_035_),
    .A2(\state[0] ),
    .A3(net3),
    .A4(_034_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _170_ (.A1(_047_),
    .A2(_050_),
    .A3(_055_),
    .A4(_058_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _171_ (.A1(\miso_capture[0] ),
    .A2(_037_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _172_ (.A1(_056_),
    .A2(_057_),
    .B(_059_),
    .C(_060_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _173_ (.A1(_043_),
    .A2(_048_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _174_ (.A1(_051_),
    .A2(_052_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _175_ (.A1(\bit_counter[0] ),
    .A2(_049_),
    .A3(_062_),
    .A4(_058_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _176_ (.A1(\state[1] ),
    .A2(\state[0] ),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _177_ (.A1(\miso_capture[1] ),
    .A2(_064_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _178_ (.A1(_112_),
    .A2(_039_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _179_ (.A1(_046_),
    .A2(_036_),
    .A3(_066_),
    .A4(_061_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _180_ (.A1(_046_),
    .A2(_061_),
    .A3(_063_),
    .B1(_065_),
    .B2(_067_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _181_ (.A1(_121_),
    .A2(_118_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _182_ (.A1(\bit_counter[0] ),
    .A2(_127_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _183_ (.A1(_068_),
    .A2(_051_),
    .A3(_052_),
    .A4(_069_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _184_ (.A1(\miso_capture[2] ),
    .A2(_064_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _185_ (.A1(_037_),
    .A2(_061_),
    .A3(_070_),
    .B(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _186_ (.A1(_058_),
    .A2(_061_),
    .A3(_070_),
    .B(_072_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _187_ (.A1(\bit_counter[2] ),
    .A2(_126_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _188_ (.A1(_127_),
    .A2(_130_),
    .A3(_073_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _189_ (.A1(_066_),
    .A2(_074_),
    .B(\miso_capture[3] ),
    .C(_038_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _190_ (.A1(\miso_capture[3] ),
    .A2(_037_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _191_ (.A1(_063_),
    .A2(_074_),
    .B(_075_),
    .C(_076_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _192_ (.A1(\miso_capture[4] ),
    .A2(_038_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _193_ (.A1(\bit_counter[0] ),
    .A2(_068_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _194_ (.A1(_078_),
    .A2(_062_),
    .A3(_074_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _195_ (.A1(_078_),
    .A2(_062_),
    .A3(_058_),
    .A4(_074_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _196_ (.A1(\miso_capture[4] ),
    .A2(_037_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _197_ (.A1(_077_),
    .A2(_079_),
    .B(_080_),
    .C(_081_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _198_ (.A1(_043_),
    .A2(_073_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _199_ (.A1(_046_),
    .A2(_037_),
    .A3(_066_),
    .A4(_082_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _200_ (.A1(\miso_capture[5] ),
    .A2(_064_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _201_ (.A1(_046_),
    .A2(_063_),
    .A3(_082_),
    .B1(_083_),
    .B2(_084_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _202_ (.A1(\miso_capture[6] ),
    .A2(_064_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _203_ (.A1(_037_),
    .A2(_070_),
    .A3(_082_),
    .B(_085_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _204_ (.A1(_058_),
    .A2(_070_),
    .A3(_082_),
    .B(_086_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _205_ (.A1(_127_),
    .A2(_130_),
    .A3(_048_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _206_ (.A1(\miso_capture[7] ),
    .A2(_064_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _207_ (.A1(_037_),
    .A2(_066_),
    .A3(_087_),
    .B(_088_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _208_ (.A1(_063_),
    .A2(_087_),
    .B(_089_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _209_ (.I0(\miso_capture[0] ),
    .I1(net13),
    .S(_111_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _210_ (.I0(\miso_capture[1] ),
    .I1(net14),
    .S(_111_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _211_ (.I0(\miso_capture[2] ),
    .I1(net15),
    .S(_111_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _212_ (.I0(\miso_capture[3] ),
    .I1(net16),
    .S(_111_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _213_ (.I0(\miso_capture[4] ),
    .I1(net17),
    .S(_111_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _214_ (.I0(\miso_capture[5] ),
    .I1(net18),
    .S(_111_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _215_ (.I0(\miso_capture[6] ),
    .I1(net19),
    .S(_111_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _216_ (.I0(\miso_capture[7] ),
    .I1(net20),
    .S(_111_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _217_ (.A1(\state[1] ),
    .A2(net22),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _218_ (.A1(\state[0] ),
    .A2(_090_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _219_ (.I(net23),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _220_ (.A1(\state[0] ),
    .A2(_091_),
    .B1(_045_),
    .B2(net12),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _221_ (.A1(_035_),
    .A2(\state[0] ),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _222_ (.I0(net11),
    .I1(\tx_shift[6] ),
    .S(_092_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _223_ (.A1(net22),
    .A2(_116_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _224_ (.I0(net12),
    .I1(_094_),
    .S(\state[0] ),
    .Z(_095_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _225_ (.A1(_035_),
    .A2(_095_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _226_ (.I0(net24),
    .I1(_093_),
    .S(_096_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _227_ (.A1(_110_),
    .A2(net22),
    .A3(_113_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _228_ (.I(net12),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _229_ (.A1(_110_),
    .A2(_098_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _230_ (.A1(_035_),
    .A2(_097_),
    .A3(_099_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _231_ (.A1(\bit_counter[2] ),
    .A2(_126_),
    .A3(_038_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _232_ (.I0(_098_),
    .I1(net25),
    .S(_064_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _233_ (.I(\tx_shift[0] ),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _234_ (.A1(net12),
    .A2(net4),
    .A3(_045_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _235_ (.A1(_100_),
    .A2(_096_),
    .B(_101_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _236_ (.I0(net5),
    .I1(\tx_shift[0] ),
    .S(_092_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _237_ (.I0(\tx_shift[1] ),
    .I1(_102_),
    .S(_096_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _238_ (.I0(net6),
    .I1(\tx_shift[1] ),
    .S(_092_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _239_ (.I0(\tx_shift[2] ),
    .I1(_103_),
    .S(_096_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _240_ (.I0(net7),
    .I1(\tx_shift[2] ),
    .S(_092_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _241_ (.I0(\tx_shift[3] ),
    .I1(_104_),
    .S(_096_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _242_ (.I0(net8),
    .I1(\tx_shift[3] ),
    .S(_092_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _243_ (.I0(\tx_shift[4] ),
    .I1(_105_),
    .S(_096_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _244_ (.I0(net9),
    .I1(\tx_shift[4] ),
    .S(_092_),
    .Z(_106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _245_ (.I0(\tx_shift[5] ),
    .I1(_106_),
    .S(_096_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _246_ (.I0(net10),
    .I1(\tx_shift[5] ),
    .S(_092_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _247_ (.I0(\tx_shift[6] ),
    .I1(_107_),
    .S(_096_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _248_ (.A(_112_),
    .B(_113_),
    .CO(_114_),
    .S(_115_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _249_ (.A(_112_),
    .B(_113_),
    .CO(_116_),
    .S(_117_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _250_ (.A(\bit_counter[3] ),
    .B(_113_),
    .CO(_118_),
    .S(_119_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _251_ (.A(\bit_counter[3] ),
    .B(_120_),
    .CO(_121_),
    .S(_122_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _252_ (.A(_112_),
    .B(_123_),
    .CO(_124_),
    .S(_125_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _253_ (.A(\bit_counter[0] ),
    .B(\bit_counter[1] ),
    .CO(_126_),
    .S(_127_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _254_ (.A(_112_),
    .B(_128_),
    .CO(_129_),
    .S(_130_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[0]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\bit_counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[1]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\bit_counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[2]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\bit_counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[3]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \miso_capture[0]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\miso_capture[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \miso_capture[1]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\miso_capture[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \miso_capture[2]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\miso_capture[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \miso_capture[3]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\miso_capture[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \miso_capture[4]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\miso_capture[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \miso_capture[5]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\miso_capture[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \miso_capture[6]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\miso_capture[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \miso_capture[7]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\miso_capture[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[0]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[1]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[2]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[3]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[4]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[5]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[6]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[7]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_valid$_DFF_PN0_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_clk$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \spi_cs_n$_DFFE_PN1P_  (.D(_022_),
    .SETN(net2),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_mosi$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[0]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[1]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \tx_ready$_DFFE_PN1P_  (.D(_026_),
    .SETN(net2),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[0]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[1]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[2]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[3]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\tx_shift[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[4]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\tx_shift[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[5]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\tx_shift[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[6]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\tx_shift[6] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 hold1 (.I(net2),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_65 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(net26),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(spi_miso),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(tx_data[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(tx_data[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(tx_data[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(tx_data[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(tx_data[4]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(tx_data[5]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(tx_data[6]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(tx_data[7]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input11 (.I(tx_valid),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(rx_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(rx_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(rx_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(rx_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(rx_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(rx_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(rx_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(rx_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(rx_valid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(spi_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(spi_cs_n));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(spi_mosi));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net25),
    .Z(tx_ready));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload1 (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload2 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_246 ();
endmodule
