module clock_domain_crossing_fifo (rd_almost_empty,
    rd_clk,
    rd_empty,
    rd_en,
    rd_rst_n,
    wr_almost_full,
    wr_clk,
    wr_en,
    wr_full,
    wr_rst_n,
    rd_count,
    rd_data,
    wr_count,
    wr_data);
 output rd_almost_empty;
 input rd_clk;
 output rd_empty;
 input rd_en;
 input rd_rst_n;
 output wr_almost_full;
 input wr_clk;
 input wr_en;
 output wr_full;
 input wr_rst_n;
 output [4:0] rd_count;
 output [31:0] rd_data;
 output [4:0] wr_count;
 input [31:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire \rd_ptr_bin[0] ;
 wire \rd_ptr_bin[1] ;
 wire \rd_ptr_bin[2] ;
 wire \rd_ptr_bin[3] ;
 wire \rd_ptr_bin[4] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray[3] ;
 wire \rd_ptr_gray_sync1[0] ;
 wire \rd_ptr_gray_sync1[1] ;
 wire \rd_ptr_gray_sync1[2] ;
 wire \rd_ptr_gray_sync1[3] ;
 wire \rd_ptr_gray_sync1[4] ;
 wire \rd_ptr_gray_sync2[0] ;
 wire \rd_ptr_gray_sync2[1] ;
 wire \rd_ptr_gray_sync2[2] ;
 wire \rd_ptr_gray_sync2[3] ;
 wire \rd_ptr_gray_sync2[4] ;
 wire \wr_ptr_bin[0] ;
 wire \wr_ptr_bin[1] ;
 wire \wr_ptr_bin[2] ;
 wire \wr_ptr_bin[3] ;
 wire \wr_ptr_bin[4] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray[3] ;
 wire \wr_ptr_gray_sync1[0] ;
 wire \wr_ptr_gray_sync1[1] ;
 wire \wr_ptr_gray_sync1[2] ;
 wire \wr_ptr_gray_sync1[3] ;
 wire \wr_ptr_gray_sync1[4] ;
 wire \wr_ptr_gray_sync2[0] ;
 wire \wr_ptr_gray_sync2[1] ;
 wire \wr_ptr_gray_sync2[2] ;
 wire \wr_ptr_gray_sync2[3] ;
 wire \wr_ptr_gray_sync2[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;

 sky130_fd_sc_hd__xnor2_1 _0889_ (.A(\rd_ptr_gray_sync2[3] ),
    .B(\rd_ptr_gray_sync2[4] ),
    .Y(_0856_));
 sky130_fd_sc_hd__xor2_1 _0890_ (.A(\rd_ptr_gray_sync2[2] ),
    .B(_0856_),
    .X(_0853_));
 sky130_fd_sc_hd__xor2_1 _0891_ (.A(\rd_ptr_gray_sync2[1] ),
    .B(_0853_),
    .X(_0846_));
 sky130_fd_sc_hd__inv_1 _0892_ (.A(_0888_),
    .Y(net79));
 sky130_fd_sc_hd__xnor2_4 _0893_ (.A(\rd_ptr_gray_sync2[4] ),
    .B(\wr_ptr_bin[4] ),
    .Y(_0590_));
 sky130_fd_sc_hd__nand4_2 _0894_ (.A(_0858_),
    .B(_0855_),
    .C(_0852_),
    .D(_0888_),
    .Y(_0591_));
 sky130_fd_sc_hd__nor2_1 _0895_ (.A(_0590_),
    .B(_0591_),
    .Y(net84));
 sky130_fd_sc_hd__clkbuf_4 _0896_ (.A(\wr_ptr_bin[2] ),
    .X(_0592_));
 sky130_fd_sc_hd__clkbuf_4 _0897_ (.A(\wr_ptr_bin[3] ),
    .X(_0593_));
 sky130_fd_sc_hd__nor2b_1 _0898_ (.A(net84),
    .B_N(net37),
    .Y(_0594_));
 sky130_fd_sc_hd__clkbuf_4 _0899_ (.A(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__nand3_4 _0900_ (.A(_0592_),
    .B(_0593_),
    .C(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_8 _0901_ (.A(net38),
    .B(_0872_),
    .Y(_0597_));
 sky130_fd_sc_hd__nor2_8 _0902_ (.A(_0596_),
    .B(_0597_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_1 _0903_ (.A(_0842_),
    .Y(_0598_));
 sky130_fd_sc_hd__a21o_1 _0904_ (.A1(_0598_),
    .A2(_0852_),
    .B1(_0851_),
    .X(_0599_));
 sky130_fd_sc_hd__a21oi_1 _0905_ (.A1(_0855_),
    .A2(_0599_),
    .B1(_0854_),
    .Y(_0600_));
 sky130_fd_sc_hd__xnor2_1 _0906_ (.A(_0858_),
    .B(_0600_),
    .Y(net82));
 sky130_fd_sc_hd__inv_1 _0907_ (.A(_0844_),
    .Y(_0601_));
 sky130_fd_sc_hd__a21o_1 _0908_ (.A1(_0601_),
    .A2(_0855_),
    .B1(_0854_),
    .X(_0602_));
 sky130_fd_sc_hd__a21oi_1 _0909_ (.A1(_0858_),
    .A2(_0602_),
    .B1(_0857_),
    .Y(_0603_));
 sky130_fd_sc_hd__xnor2_1 _0910_ (.A(_0590_),
    .B(_0603_),
    .Y(net83));
 sky130_fd_sc_hd__nand2_8 _0911_ (.A(net38),
    .B(_0871_),
    .Y(_0604_));
 sky130_fd_sc_hd__o21ai_4 _0912_ (.A1(_0590_),
    .A2(_0591_),
    .B1(net37),
    .Y(_0605_));
 sky130_fd_sc_hd__or3_4 _0913_ (.A(_0592_),
    .B(_0593_),
    .C(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__nor2_8 _0914_ (.A(_0604_),
    .B(_0606_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_8 _0915_ (.A(net38),
    .B(_0874_),
    .Y(_0607_));
 sky130_fd_sc_hd__nor2_8 _0916_ (.A(_0606_),
    .B(_0607_),
    .Y(_0014_));
 sky130_fd_sc_hd__nor2_8 _0917_ (.A(_0597_),
    .B(_0606_),
    .Y(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _0918_ (.A(_0876_),
    .X(_0608_));
 sky130_fd_sc_hd__nand2_8 _0919_ (.A(net38),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor2_8 _0920_ (.A(_0606_),
    .B(_0609_),
    .Y(_0012_));
 sky130_fd_sc_hd__nand3b_4 _0921_ (.A_N(_0593_),
    .B(_0595_),
    .C(_0592_),
    .Y(_0610_));
 sky130_fd_sc_hd__nor2_8 _0922_ (.A(_0604_),
    .B(_0610_),
    .Y(_0011_));
 sky130_fd_sc_hd__nor2_8 _0923_ (.A(_0607_),
    .B(_0610_),
    .Y(_0010_));
 sky130_fd_sc_hd__nor2_8 _0924_ (.A(_0597_),
    .B(_0610_),
    .Y(_0009_));
 sky130_fd_sc_hd__nor2_8 _0925_ (.A(_0609_),
    .B(_0610_),
    .Y(_0008_));
 sky130_fd_sc_hd__nand3b_4 _0926_ (.A_N(_0592_),
    .B(_0593_),
    .C(_0595_),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_8 _0927_ (.A(_0604_),
    .B(_0611_),
    .Y(_0007_));
 sky130_fd_sc_hd__nor2_8 _0928_ (.A(_0607_),
    .B(_0611_),
    .Y(_0006_));
 sky130_fd_sc_hd__nor2_8 _0929_ (.A(_0597_),
    .B(_0611_),
    .Y(_0005_));
 sky130_fd_sc_hd__nor2_8 _0930_ (.A(_0609_),
    .B(_0611_),
    .Y(_0004_));
 sky130_fd_sc_hd__nor2_8 _0931_ (.A(_0596_),
    .B(_0604_),
    .Y(_0003_));
 sky130_fd_sc_hd__nor2_8 _0932_ (.A(_0596_),
    .B(_0609_),
    .Y(_0000_));
 sky130_fd_sc_hd__nor2_8 _0933_ (.A(_0596_),
    .B(_0607_),
    .Y(_0002_));
 sky130_fd_sc_hd__xor2_1 _0934_ (.A(\wr_ptr_gray_sync2[3] ),
    .B(\wr_ptr_gray_sync2[4] ),
    .X(_0864_));
 sky130_fd_sc_hd__xnor2_1 _0935_ (.A(\wr_ptr_gray_sync2[2] ),
    .B(_0864_),
    .Y(_0612_));
 sky130_fd_sc_hd__xor2_2 _0936_ (.A(\wr_ptr_gray_sync2[1] ),
    .B(_0612_),
    .X(_0848_));
 sky130_fd_sc_hd__inv_1 _0937_ (.A(_0850_),
    .Y(net41));
 sky130_fd_sc_hd__xnor2_1 _0938_ (.A(_0849_),
    .B(_0870_),
    .Y(net42));
 sky130_fd_sc_hd__inv_1 _0939_ (.A(_0847_),
    .Y(_0613_));
 sky130_fd_sc_hd__a21o_1 _0940_ (.A1(_0862_),
    .A2(_0613_),
    .B1(_0861_),
    .X(_0614_));
 sky130_fd_sc_hd__a21oi_1 _0941_ (.A1(_0870_),
    .A2(_0614_),
    .B1(_0869_),
    .Y(_0615_));
 sky130_fd_sc_hd__xnor2_1 _0942_ (.A(_0866_),
    .B(_0615_),
    .Y(net43));
 sky130_fd_sc_hd__xor2_1 _0943_ (.A(\wr_ptr_gray_sync2[4] ),
    .B(\rd_ptr_bin[4] ),
    .X(_0616_));
 sky130_fd_sc_hd__inv_1 _0944_ (.A(_0849_),
    .Y(_0617_));
 sky130_fd_sc_hd__a21o_1 _0945_ (.A1(_0617_),
    .A2(_0870_),
    .B1(_0869_),
    .X(_0618_));
 sky130_fd_sc_hd__a21oi_1 _0946_ (.A1(_0866_),
    .A2(_0618_),
    .B1(_0865_),
    .Y(_0619_));
 sky130_fd_sc_hd__xor2_1 _0947_ (.A(_0616_),
    .B(_0619_),
    .X(net44));
 sky130_fd_sc_hd__xor2_1 _0948_ (.A(\wr_ptr_gray_sync2[2] ),
    .B(\rd_ptr_gray[2] ),
    .X(_0620_));
 sky130_fd_sc_hd__xor2_1 _0949_ (.A(\wr_ptr_gray_sync2[1] ),
    .B(\rd_ptr_gray[1] ),
    .X(_0621_));
 sky130_fd_sc_hd__xor2_1 _0950_ (.A(\wr_ptr_gray_sync2[0] ),
    .B(\rd_ptr_gray[0] ),
    .X(_0622_));
 sky130_fd_sc_hd__xor2_1 _0951_ (.A(\wr_ptr_gray_sync2[3] ),
    .B(\rd_ptr_gray[3] ),
    .X(_0623_));
 sky130_fd_sc_hd__or3_1 _0952_ (.A(_0616_),
    .B(_0622_),
    .C(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__or3_1 _0953_ (.A(_0620_),
    .B(_0621_),
    .C(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__inv_1 _0954_ (.A(_0625_),
    .Y(net77));
 sky130_fd_sc_hd__buf_4 _0955_ (.A(\rd_ptr_bin[2] ),
    .X(_0626_));
 sky130_fd_sc_hd__inv_2 _0956_ (.A(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__clkbuf_4 _0957_ (.A(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__clkbuf_8 _0958_ (.A(_0628_),
    .X(_0867_));
 sky130_fd_sc_hd__buf_4 _0959_ (.A(\rd_ptr_bin[3] ),
    .X(_0629_));
 sky130_fd_sc_hd__clkinv_2 _0960_ (.A(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__buf_6 _0961_ (.A(_0630_),
    .X(_0863_));
 sky130_fd_sc_hd__inv_1 _0962_ (.A(_0846_),
    .Y(_0843_));
 sky130_fd_sc_hd__clkbuf_2 _0963_ (.A(\wr_ptr_bin[0] ),
    .X(_0631_));
 sky130_fd_sc_hd__inv_1 _0964_ (.A(_0631_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_1 _0965_ (.A(\rd_ptr_bin[0] ),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_1 _0966_ (.A(_0848_),
    .Y(_0860_));
 sky130_fd_sc_hd__inv_1 _0967_ (.A(_0612_),
    .Y(_0868_));
 sky130_fd_sc_hd__clkinvlp_4 _0968_ (.A(\wr_ptr_bin[1] ),
    .Y(_0841_));
 sky130_fd_sc_hd__inv_1 _0969_ (.A(\rd_ptr_bin[1] ),
    .Y(_0859_));
 sky130_fd_sc_hd__xor2_1 _0970_ (.A(\wr_ptr_gray_sync2[0] ),
    .B(_0848_),
    .X(_0885_));
 sky130_fd_sc_hd__xnor2_1 _0971_ (.A(\rd_ptr_gray_sync2[0] ),
    .B(_0846_),
    .Y(_0887_));
 sky130_fd_sc_hd__inv_1 _0972_ (.A(_0886_),
    .Y(net40));
 sky130_fd_sc_hd__o31ai_4 _0973_ (.A1(_0620_),
    .A2(_0621_),
    .A3(_0624_),
    .B1(net2),
    .Y(_0632_));
 sky130_fd_sc_hd__buf_6 _0974_ (.A(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_4 _0975_ (.A(_0878_),
    .X(_0634_));
 sky130_fd_sc_hd__o21ai_2 _0976_ (.A1(\rd_ptr_bin[3] ),
    .A2(\rd_ptr_bin[2] ),
    .B1(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__buf_4 _0977_ (.A(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_4 _0978_ (.A(_0883_),
    .X(_0637_));
 sky130_fd_sc_hd__buf_4 _0979_ (.A(_0881_),
    .X(_0638_));
 sky130_fd_sc_hd__nor3_2 _0980_ (.A(_0637_),
    .B(_0879_),
    .C(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__buf_4 _0981_ (.A(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__nand2_2 _0982_ (.A(_0636_),
    .B(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__nor2_1 _0983_ (.A(\mem[0][0] ),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nor2_1 _0984_ (.A(_0633_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__clkbuf_8 _0985_ (.A(_0629_),
    .X(_0644_));
 sky130_fd_sc_hd__buf_4 _0986_ (.A(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__buf_4 _0987_ (.A(_0879_),
    .X(_0646_));
 sky130_fd_sc_hd__buf_4 _0988_ (.A(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__buf_6 _0989_ (.A(_0626_),
    .X(_0648_));
 sky130_fd_sc_hd__clkbuf_4 _0990_ (.A(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__a21oi_1 _0991_ (.A1(\mem[10][0] ),
    .A2(_0647_),
    .B1(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__clkbuf_8 _0992_ (.A(_0634_),
    .X(_0651_));
 sky130_fd_sc_hd__buf_4 _0993_ (.A(_0638_),
    .X(_0652_));
 sky130_fd_sc_hd__a22oi_1 _0994_ (.A1(\mem[12][0] ),
    .A2(_0651_),
    .B1(_0652_),
    .B2(\mem[13][0] ),
    .Y(_0653_));
 sky130_fd_sc_hd__buf_4 _0995_ (.A(_0648_),
    .X(_0654_));
 sky130_fd_sc_hd__buf_4 _0996_ (.A(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__nor2b_1 _0997_ (.A(_0626_),
    .B_N(_0637_),
    .Y(_0656_));
 sky130_fd_sc_hd__buf_6 _0998_ (.A(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__buf_6 _0999_ (.A(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_4 _1000_ (.A(_0629_),
    .X(_0659_));
 sky130_fd_sc_hd__buf_4 _1001_ (.A(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__a21oi_1 _1002_ (.A1(\mem[3][0] ),
    .A2(_0658_),
    .B1(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__a221o_1 _1003_ (.A1(_0645_),
    .A2(_0650_),
    .B1(_0653_),
    .B2(_0655_),
    .C1(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__buf_6 _1004_ (.A(_0644_),
    .X(_0663_));
 sky130_fd_sc_hd__clkbuf_4 _1005_ (.A(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__buf_4 _1006_ (.A(_0649_),
    .X(_0665_));
 sky130_fd_sc_hd__clkbuf_8 _1007_ (.A(_0879_),
    .X(_0666_));
 sky130_fd_sc_hd__clkbuf_4 _1008_ (.A(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__nand2_1 _1009_ (.A(\mem[2][0] ),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__buf_4 _1010_ (.A(_0634_),
    .X(_0669_));
 sky130_fd_sc_hd__buf_4 _1011_ (.A(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__nand3_1 _1012_ (.A(_0665_),
    .B(\mem[4][0] ),
    .C(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__o21ai_0 _1013_ (.A1(_0665_),
    .A2(_0668_),
    .B1(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__buf_4 _1014_ (.A(_0649_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_4 _1015_ (.A(_0638_),
    .X(_0674_));
 sky130_fd_sc_hd__buf_4 _1016_ (.A(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__nand2_1 _1017_ (.A(\mem[9][0] ),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__buf_6 _1018_ (.A(_0646_),
    .X(_0677_));
 sky130_fd_sc_hd__buf_4 _1019_ (.A(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__nand3_1 _1020_ (.A(_0665_),
    .B(\mem[14][0] ),
    .C(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__o211ai_1 _1021_ (.A1(_0673_),
    .A2(_0676_),
    .B1(_0679_),
    .C1(_0664_),
    .Y(_0680_));
 sky130_fd_sc_hd__o21ai_0 _1022_ (.A1(_0664_),
    .A2(_0672_),
    .B1(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__buf_4 _1023_ (.A(_0630_),
    .X(_0682_));
 sky130_fd_sc_hd__buf_4 _1024_ (.A(_0646_),
    .X(_0683_));
 sky130_fd_sc_hd__and2_0 _1025_ (.A(\rd_ptr_bin[3] ),
    .B(_0637_),
    .X(_0684_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1026_ (.A(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__buf_4 _1027_ (.A(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__a32o_1 _1028_ (.A1(_0682_),
    .A2(\mem[6][0] ),
    .A3(_0683_),
    .B1(_0686_),
    .B2(\mem[15][0] ),
    .X(_0687_));
 sky130_fd_sc_hd__buf_4 _1029_ (.A(_0663_),
    .X(_0688_));
 sky130_fd_sc_hd__nand2_1 _1030_ (.A(\mem[1][0] ),
    .B(_0675_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand3_1 _1031_ (.A(_0645_),
    .B(\mem[8][0] ),
    .C(_0670_),
    .Y(_0690_));
 sky130_fd_sc_hd__o211ai_1 _1032_ (.A1(_0688_),
    .A2(_0689_),
    .B1(_0690_),
    .C1(_0867_),
    .Y(_0691_));
 sky130_fd_sc_hd__o21ai_0 _1033_ (.A1(_0867_),
    .A2(_0687_),
    .B1(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__and3b_1 _1034_ (.A_N(_0629_),
    .B(_0648_),
    .C(_0638_),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_8 _1035_ (.A(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__nor2b_1 _1036_ (.A(_0629_),
    .B_N(_0626_),
    .Y(_0695_));
 sky130_fd_sc_hd__nor2b_4 _1037_ (.A(_0626_),
    .B_N(_0629_),
    .Y(_0696_));
 sky130_fd_sc_hd__a22o_1 _1038_ (.A1(\mem[7][0] ),
    .A2(_0695_),
    .B1(_0696_),
    .B2(\mem[11][0] ),
    .X(_0697_));
 sky130_fd_sc_hd__buf_4 _1039_ (.A(_0637_),
    .X(_0698_));
 sky130_fd_sc_hd__and2_0 _1040_ (.A(_0635_),
    .B(_0639_),
    .X(_0699_));
 sky130_fd_sc_hd__a221oi_1 _1041_ (.A1(\mem[5][0] ),
    .A2(_0694_),
    .B1(_0697_),
    .B2(_0698_),
    .C1(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__nand4_1 _1042_ (.A(_0662_),
    .B(_0681_),
    .C(_0692_),
    .D(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__a22o_1 _1043_ (.A1(net45),
    .A2(_0633_),
    .B1(_0643_),
    .B2(_0701_),
    .X(_0020_));
 sky130_fd_sc_hd__buf_4 _1044_ (.A(_0632_),
    .X(_0702_));
 sky130_fd_sc_hd__clkbuf_4 _1045_ (.A(_0648_),
    .X(_0703_));
 sky130_fd_sc_hd__clkbuf_4 _1046_ (.A(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__a22oi_1 _1047_ (.A1(_0698_),
    .A2(\mem[15][10] ),
    .B1(\mem[14][10] ),
    .B2(_0647_),
    .Y(_0705_));
 sky130_fd_sc_hd__buf_4 _1048_ (.A(_0646_),
    .X(_0706_));
 sky130_fd_sc_hd__a221oi_1 _1049_ (.A1(_0698_),
    .A2(\mem[7][10] ),
    .B1(\mem[6][10] ),
    .B2(_0706_),
    .C1(_0663_),
    .Y(_0707_));
 sky130_fd_sc_hd__a21oi_1 _1050_ (.A1(_0660_),
    .A2(_0705_),
    .B1(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__buf_4 _1051_ (.A(_0634_),
    .X(_0709_));
 sky130_fd_sc_hd__buf_4 _1052_ (.A(_0638_),
    .X(_0710_));
 sky130_fd_sc_hd__buf_4 _1053_ (.A(_0629_),
    .X(_0711_));
 sky130_fd_sc_hd__clkbuf_4 _1054_ (.A(_0626_),
    .X(_0712_));
 sky130_fd_sc_hd__nand2_4 _1055_ (.A(_0711_),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__a221oi_1 _1056_ (.A1(\mem[12][10] ),
    .A2(_0709_),
    .B1(_0710_),
    .B2(\mem[13][10] ),
    .C1(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__nand2b_2 _1057_ (.A_N(_0629_),
    .B(_0648_),
    .Y(_0715_));
 sky130_fd_sc_hd__a221oi_1 _1058_ (.A1(\mem[4][10] ),
    .A2(_0709_),
    .B1(_0710_),
    .B2(\mem[5][10] ),
    .C1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__buf_4 _1059_ (.A(_0638_),
    .X(_0717_));
 sky130_fd_sc_hd__a22oi_1 _1060_ (.A1(\mem[10][10] ),
    .A2(_0646_),
    .B1(_0717_),
    .B2(\mem[9][10] ),
    .Y(_0718_));
 sky130_fd_sc_hd__buf_6 _1061_ (.A(_0637_),
    .X(_0719_));
 sky130_fd_sc_hd__a22oi_1 _1062_ (.A1(_0719_),
    .A2(\mem[3][10] ),
    .B1(\mem[2][10] ),
    .B2(_0666_),
    .Y(_0720_));
 sky130_fd_sc_hd__nor2_4 _1063_ (.A(_0644_),
    .B(_0648_),
    .Y(_0721_));
 sky130_fd_sc_hd__a22o_1 _1064_ (.A1(_0696_),
    .A2(_0718_),
    .B1(_0720_),
    .B2(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__nor3_1 _1065_ (.A(_0714_),
    .B(_0716_),
    .C(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__a32oi_1 _1066_ (.A1(_0682_),
    .A2(\mem[1][10] ),
    .A3(_0652_),
    .B1(_0686_),
    .B2(\mem[11][10] ),
    .Y(_0724_));
 sky130_fd_sc_hd__nand3_1 _1067_ (.A(_0660_),
    .B(\mem[8][10] ),
    .C(_0670_),
    .Y(_0725_));
 sky130_fd_sc_hd__a21oi_1 _1068_ (.A1(_0724_),
    .A2(_0725_),
    .B1(_0673_),
    .Y(_0726_));
 sky130_fd_sc_hd__clkbuf_8 _1069_ (.A(_0699_),
    .X(_0727_));
 sky130_fd_sc_hd__a2111oi_0 _1070_ (.A1(_0704_),
    .A2(_0708_),
    .B1(_0723_),
    .C1(_0726_),
    .D1(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__buf_4 _1071_ (.A(_0641_),
    .X(_0729_));
 sky130_fd_sc_hd__nor2_1 _1072_ (.A(\mem[0][10] ),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__buf_4 _1073_ (.A(_0633_),
    .X(_0731_));
 sky130_fd_sc_hd__nand2_1 _1074_ (.A(net46),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__o31ai_1 _1075_ (.A1(_0702_),
    .A2(_0728_),
    .A3(_0730_),
    .B1(_0732_),
    .Y(_0021_));
 sky130_fd_sc_hd__buf_6 _1076_ (.A(_0657_),
    .X(_0733_));
 sky130_fd_sc_hd__clkbuf_4 _1077_ (.A(_0644_),
    .X(_0734_));
 sky130_fd_sc_hd__a21oi_1 _1078_ (.A1(\mem[3][11] ),
    .A2(_0733_),
    .B1(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__buf_6 _1079_ (.A(_0637_),
    .X(_0736_));
 sky130_fd_sc_hd__buf_4 _1080_ (.A(_0646_),
    .X(_0737_));
 sky130_fd_sc_hd__a222oi_1 _1081_ (.A1(_0736_),
    .A2(\mem[7][11] ),
    .B1(\mem[4][11] ),
    .B2(_0669_),
    .C1(_0737_),
    .C2(\mem[6][11] ),
    .Y(_0738_));
 sky130_fd_sc_hd__nor2b_1 _1082_ (.A(\rd_ptr_bin[2] ),
    .B_N(_0879_),
    .Y(_0739_));
 sky130_fd_sc_hd__buf_2 _1083_ (.A(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__clkbuf_4 _1084_ (.A(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__buf_4 _1085_ (.A(_0630_),
    .X(_0742_));
 sky130_fd_sc_hd__a21oi_1 _1086_ (.A1(\mem[10][11] ),
    .A2(_0741_),
    .B1(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__clkbuf_4 _1087_ (.A(_0638_),
    .X(_0744_));
 sky130_fd_sc_hd__a222oi_1 _1088_ (.A1(\mem[14][11] ),
    .A2(_0677_),
    .B1(_0744_),
    .B2(\mem[13][11] ),
    .C1(\mem[12][11] ),
    .C2(_0651_),
    .Y(_0745_));
 sky130_fd_sc_hd__a22oi_1 _1089_ (.A1(_0735_),
    .A2(_0738_),
    .B1(_0743_),
    .B2(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__o21ai_0 _1090_ (.A1(_0735_),
    .A2(_0743_),
    .B1(_0867_),
    .Y(_0747_));
 sky130_fd_sc_hd__buf_4 _1091_ (.A(_0630_),
    .X(_0748_));
 sky130_fd_sc_hd__buf_4 _1092_ (.A(_0685_),
    .X(_0749_));
 sky130_fd_sc_hd__a32oi_1 _1093_ (.A1(_0748_),
    .A2(\mem[1][11] ),
    .A3(_0652_),
    .B1(_0749_),
    .B2(\mem[11][11] ),
    .Y(_0750_));
 sky130_fd_sc_hd__clkbuf_4 _1094_ (.A(_0628_),
    .X(_0751_));
 sky130_fd_sc_hd__buf_4 _1095_ (.A(_0626_),
    .X(_0752_));
 sky130_fd_sc_hd__buf_2 _1096_ (.A(_0638_),
    .X(_0753_));
 sky130_fd_sc_hd__and3_1 _1097_ (.A(_0752_),
    .B(\mem[5][11] ),
    .C(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__a31oi_1 _1098_ (.A1(_0751_),
    .A2(\mem[2][11] ),
    .A3(_0683_),
    .B1(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__o22ai_1 _1099_ (.A1(_0665_),
    .A2(_0750_),
    .B1(_0755_),
    .B2(_0664_),
    .Y(_0756_));
 sky130_fd_sc_hd__nand2_4 _1100_ (.A(_0629_),
    .B(_0627_),
    .Y(_0757_));
 sky130_fd_sc_hd__buf_4 _1101_ (.A(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__buf_4 _1102_ (.A(_0634_),
    .X(_0759_));
 sky130_fd_sc_hd__buf_6 _1103_ (.A(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__a22oi_1 _1104_ (.A1(\mem[8][11] ),
    .A2(_0760_),
    .B1(_0675_),
    .B2(\mem[9][11] ),
    .Y(_0761_));
 sky130_fd_sc_hd__and3_1 _1105_ (.A(_0629_),
    .B(_0626_),
    .C(_0637_),
    .X(_0762_));
 sky130_fd_sc_hd__buf_4 _1106_ (.A(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__buf_4 _1107_ (.A(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__nand2_1 _1108_ (.A(\mem[15][11] ),
    .B(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__o21ai_0 _1109_ (.A1(_0758_),
    .A2(_0761_),
    .B1(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__a2111oi_1 _1110_ (.A1(_0746_),
    .A2(_0747_),
    .B1(_0727_),
    .C1(_0756_),
    .D1(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__nor2_1 _1111_ (.A(\mem[0][11] ),
    .B(_0729_),
    .Y(_0768_));
 sky130_fd_sc_hd__nand2_1 _1112_ (.A(net47),
    .B(_0731_),
    .Y(_0769_));
 sky130_fd_sc_hd__o31ai_1 _1113_ (.A1(_0702_),
    .A2(_0767_),
    .A3(_0768_),
    .B1(_0769_),
    .Y(_0022_));
 sky130_fd_sc_hd__buf_4 _1114_ (.A(_0644_),
    .X(_0770_));
 sky130_fd_sc_hd__and3_1 _1115_ (.A(_0770_),
    .B(_0703_),
    .C(\mem[14][12] ),
    .X(_0771_));
 sky130_fd_sc_hd__nor3b_1 _1116_ (.A(_0663_),
    .B(_0649_),
    .C_N(\mem[2][12] ),
    .Y(_0772_));
 sky130_fd_sc_hd__o21ai_0 _1117_ (.A1(_0771_),
    .A2(_0772_),
    .B1(_0678_),
    .Y(_0773_));
 sky130_fd_sc_hd__and3_1 _1118_ (.A(_0770_),
    .B(\mem[12][12] ),
    .C(_0709_),
    .X(_0774_));
 sky130_fd_sc_hd__and3b_1 _1119_ (.A_N(_0711_),
    .B(\mem[6][12] ),
    .C(_0677_),
    .X(_0775_));
 sky130_fd_sc_hd__o21ai_0 _1120_ (.A1(_0774_),
    .A2(_0775_),
    .B1(_0673_),
    .Y(_0776_));
 sky130_fd_sc_hd__a32oi_1 _1121_ (.A1(\mem[1][12] ),
    .A2(_0675_),
    .A3(_0721_),
    .B1(_0636_),
    .B2(_0640_),
    .Y(_0777_));
 sky130_fd_sc_hd__and3b_1 _1122_ (.A_N(_0711_),
    .B(_0703_),
    .C(\mem[7][12] ),
    .X(_0778_));
 sky130_fd_sc_hd__and3b_1 _1123_ (.A_N(_0703_),
    .B(\mem[11][12] ),
    .C(_0659_),
    .X(_0779_));
 sky130_fd_sc_hd__o21ai_0 _1124_ (.A1(_0778_),
    .A2(_0779_),
    .B1(_0698_),
    .Y(_0780_));
 sky130_fd_sc_hd__nand4_1 _1125_ (.A(_0773_),
    .B(_0776_),
    .C(_0777_),
    .D(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__a22oi_1 _1126_ (.A1(\mem[8][12] ),
    .A2(_0670_),
    .B1(_0675_),
    .B2(\mem[9][12] ),
    .Y(_0782_));
 sky130_fd_sc_hd__buf_4 _1127_ (.A(_0752_),
    .X(_0783_));
 sky130_fd_sc_hd__a32oi_1 _1128_ (.A1(_0783_),
    .A2(\mem[4][12] ),
    .A3(_0760_),
    .B1(_0658_),
    .B2(\mem[3][12] ),
    .Y(_0784_));
 sky130_fd_sc_hd__nand2_1 _1129_ (.A(\mem[15][12] ),
    .B(_0764_),
    .Y(_0785_));
 sky130_fd_sc_hd__o221ai_1 _1130_ (.A1(_0758_),
    .A2(_0782_),
    .B1(_0784_),
    .B2(_0664_),
    .C1(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__nand2_1 _1131_ (.A(\mem[10][12] ),
    .B(_0683_),
    .Y(_0787_));
 sky130_fd_sc_hd__nand3_1 _1132_ (.A(_0649_),
    .B(\mem[13][12] ),
    .C(_0652_),
    .Y(_0788_));
 sky130_fd_sc_hd__o21ai_0 _1133_ (.A1(_0783_),
    .A2(_0787_),
    .B1(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__a22o_1 _1134_ (.A1(\mem[5][12] ),
    .A2(_0694_),
    .B1(_0789_),
    .B2(_0664_),
    .X(_0790_));
 sky130_fd_sc_hd__nor3_1 _1135_ (.A(_0781_),
    .B(_0786_),
    .C(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__nor2_1 _1136_ (.A(\mem[0][12] ),
    .B(_0729_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand2_1 _1137_ (.A(net48),
    .B(_0731_),
    .Y(_0793_));
 sky130_fd_sc_hd__o31ai_1 _1138_ (.A1(_0702_),
    .A2(_0791_),
    .A3(_0792_),
    .B1(_0793_),
    .Y(_0023_));
 sky130_fd_sc_hd__a21oi_1 _1139_ (.A1(\mem[3][13] ),
    .A2(_0733_),
    .B1(_0734_),
    .Y(_0794_));
 sky130_fd_sc_hd__a222oi_1 _1140_ (.A1(_0736_),
    .A2(\mem[7][13] ),
    .B1(\mem[4][13] ),
    .B2(_0669_),
    .C1(_0737_),
    .C2(\mem[6][13] ),
    .Y(_0795_));
 sky130_fd_sc_hd__a21oi_1 _1141_ (.A1(\mem[10][13] ),
    .A2(_0741_),
    .B1(_0742_),
    .Y(_0796_));
 sky130_fd_sc_hd__a222oi_1 _1142_ (.A1(\mem[14][13] ),
    .A2(_0677_),
    .B1(_0744_),
    .B2(\mem[13][13] ),
    .C1(\mem[12][13] ),
    .C2(_0651_),
    .Y(_0797_));
 sky130_fd_sc_hd__a22oi_1 _1143_ (.A1(_0794_),
    .A2(_0795_),
    .B1(_0796_),
    .B2(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__o21ai_0 _1144_ (.A1(_0794_),
    .A2(_0796_),
    .B1(_0867_),
    .Y(_0799_));
 sky130_fd_sc_hd__a32oi_1 _1145_ (.A1(_0748_),
    .A2(\mem[1][13] ),
    .A3(_0652_),
    .B1(_0749_),
    .B2(\mem[11][13] ),
    .Y(_0800_));
 sky130_fd_sc_hd__and3_1 _1146_ (.A(_0752_),
    .B(\mem[5][13] ),
    .C(_0753_),
    .X(_0801_));
 sky130_fd_sc_hd__a31oi_1 _1147_ (.A1(_0751_),
    .A2(\mem[2][13] ),
    .A3(_0683_),
    .B1(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__o22ai_1 _1148_ (.A1(_0665_),
    .A2(_0800_),
    .B1(_0802_),
    .B2(_0664_),
    .Y(_0803_));
 sky130_fd_sc_hd__a22oi_1 _1149_ (.A1(\mem[8][13] ),
    .A2(_0760_),
    .B1(_0675_),
    .B2(\mem[9][13] ),
    .Y(_0804_));
 sky130_fd_sc_hd__nand2_1 _1150_ (.A(\mem[15][13] ),
    .B(_0764_),
    .Y(_0805_));
 sky130_fd_sc_hd__o21ai_0 _1151_ (.A1(_0758_),
    .A2(_0804_),
    .B1(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__a2111oi_1 _1152_ (.A1(_0798_),
    .A2(_0799_),
    .B1(_0727_),
    .C1(_0803_),
    .D1(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__nor2_1 _1153_ (.A(\mem[0][13] ),
    .B(_0729_),
    .Y(_0808_));
 sky130_fd_sc_hd__nand2_1 _1154_ (.A(net49),
    .B(_0731_),
    .Y(_0809_));
 sky130_fd_sc_hd__o31ai_1 _1155_ (.A1(_0702_),
    .A2(_0807_),
    .A3(_0808_),
    .B1(_0809_),
    .Y(_0024_));
 sky130_fd_sc_hd__a32o_1 _1156_ (.A1(_0682_),
    .A2(\mem[6][14] ),
    .A3(_0647_),
    .B1(_0686_),
    .B2(\mem[15][14] ),
    .X(_0810_));
 sky130_fd_sc_hd__clkbuf_4 _1157_ (.A(_0711_),
    .X(_0811_));
 sky130_fd_sc_hd__nand3_1 _1158_ (.A(_0811_),
    .B(\mem[8][14] ),
    .C(_0670_),
    .Y(_0812_));
 sky130_fd_sc_hd__buf_2 _1159_ (.A(_0638_),
    .X(_0813_));
 sky130_fd_sc_hd__clkbuf_4 _1160_ (.A(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__nand3_1 _1161_ (.A(_0863_),
    .B(\mem[1][14] ),
    .C(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__clkbuf_4 _1162_ (.A(_0649_),
    .X(_0816_));
 sky130_fd_sc_hd__a21oi_1 _1163_ (.A1(_0812_),
    .A2(_0815_),
    .B1(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__clkbuf_4 _1164_ (.A(_0813_),
    .X(_0818_));
 sky130_fd_sc_hd__nand3_1 _1165_ (.A(_0783_),
    .B(\mem[13][14] ),
    .C(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__buf_4 _1166_ (.A(_0628_),
    .X(_0820_));
 sky130_fd_sc_hd__nand3_1 _1167_ (.A(_0820_),
    .B(\mem[10][14] ),
    .C(_0667_),
    .Y(_0821_));
 sky130_fd_sc_hd__clkbuf_4 _1168_ (.A(_0626_),
    .X(_0822_));
 sky130_fd_sc_hd__clkbuf_4 _1169_ (.A(_0634_),
    .X(_0823_));
 sky130_fd_sc_hd__and3_1 _1170_ (.A(_0822_),
    .B(\mem[4][14] ),
    .C(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__clkbuf_4 _1171_ (.A(_0711_),
    .X(_0825_));
 sky130_fd_sc_hd__a211oi_1 _1172_ (.A1(\mem[3][14] ),
    .A2(_0658_),
    .B1(_0824_),
    .C1(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__a31oi_1 _1173_ (.A1(_0688_),
    .A2(_0819_),
    .A3(_0821_),
    .B1(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__inv_1 _1174_ (.A(_0736_),
    .Y(_0828_));
 sky130_fd_sc_hd__buf_8 _1175_ (.A(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__buf_6 _1176_ (.A(_0695_),
    .X(_0830_));
 sky130_fd_sc_hd__buf_6 _1177_ (.A(_0696_),
    .X(_0831_));
 sky130_fd_sc_hd__a22oi_4 _1178_ (.A1(\mem[7][14] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][14] ),
    .Y(_0832_));
 sky130_fd_sc_hd__buf_2 _1179_ (.A(_0626_),
    .X(_0833_));
 sky130_fd_sc_hd__and3_1 _1180_ (.A(_0711_),
    .B(_0833_),
    .C(\mem[14][14] ),
    .X(_0834_));
 sky130_fd_sc_hd__nor3b_1 _1181_ (.A(_0770_),
    .B(_0654_),
    .C_N(\mem[2][14] ),
    .Y(_0835_));
 sky130_fd_sc_hd__o21ai_1 _1182_ (.A1(_0834_),
    .A2(_0835_),
    .B1(_0678_),
    .Y(_0836_));
 sky130_fd_sc_hd__a22oi_2 _1183_ (.A1(_0636_),
    .A2(_0640_),
    .B1(_0694_),
    .B2(\mem[5][14] ),
    .Y(_0837_));
 sky130_fd_sc_hd__and3_1 _1184_ (.A(_0703_),
    .B(\mem[12][14] ),
    .C(_0759_),
    .X(_0838_));
 sky130_fd_sc_hd__and3b_1 _1185_ (.A_N(_0712_),
    .B(\mem[9][14] ),
    .C(_0674_),
    .X(_0839_));
 sky130_fd_sc_hd__o21ai_1 _1186_ (.A1(_0838_),
    .A2(_0839_),
    .B1(_0645_),
    .Y(_0840_));
 sky130_fd_sc_hd__o2111ai_4 _1187_ (.A1(_0829_),
    .A2(_0832_),
    .B1(_0836_),
    .C1(_0837_),
    .D1(_0840_),
    .Y(_0070_));
 sky130_fd_sc_hd__a2111oi_0 _1188_ (.A1(_0704_),
    .A2(_0810_),
    .B1(_0817_),
    .C1(_0827_),
    .D1(_0070_),
    .Y(_0071_));
 sky130_fd_sc_hd__nor2_1 _1189_ (.A(\mem[0][14] ),
    .B(_0729_),
    .Y(_0072_));
 sky130_fd_sc_hd__nand2_1 _1190_ (.A(net50),
    .B(_0731_),
    .Y(_0073_));
 sky130_fd_sc_hd__o31ai_1 _1191_ (.A1(_0702_),
    .A2(_0071_),
    .A3(_0072_),
    .B1(_0073_),
    .Y(_0025_));
 sky130_fd_sc_hd__a21oi_1 _1192_ (.A1(\mem[3][15] ),
    .A2(_0733_),
    .B1(_0734_),
    .Y(_0074_));
 sky130_fd_sc_hd__a222oi_1 _1193_ (.A1(_0736_),
    .A2(\mem[7][15] ),
    .B1(\mem[4][15] ),
    .B2(_0669_),
    .C1(_0737_),
    .C2(\mem[6][15] ),
    .Y(_0075_));
 sky130_fd_sc_hd__a21oi_1 _1194_ (.A1(\mem[10][15] ),
    .A2(_0741_),
    .B1(_0742_),
    .Y(_0076_));
 sky130_fd_sc_hd__buf_4 _1195_ (.A(_0646_),
    .X(_0077_));
 sky130_fd_sc_hd__a222oi_1 _1196_ (.A1(\mem[14][15] ),
    .A2(_0077_),
    .B1(_0744_),
    .B2(\mem[13][15] ),
    .C1(\mem[12][15] ),
    .C2(_0651_),
    .Y(_0078_));
 sky130_fd_sc_hd__a22oi_1 _1197_ (.A1(_0074_),
    .A2(_0075_),
    .B1(_0076_),
    .B2(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__o21ai_0 _1198_ (.A1(_0074_),
    .A2(_0076_),
    .B1(_0867_),
    .Y(_0080_));
 sky130_fd_sc_hd__clkbuf_4 _1199_ (.A(_0630_),
    .X(_0081_));
 sky130_fd_sc_hd__a32oi_1 _1200_ (.A1(_0081_),
    .A2(\mem[1][15] ),
    .A3(_0652_),
    .B1(_0749_),
    .B2(\mem[11][15] ),
    .Y(_0082_));
 sky130_fd_sc_hd__and3_1 _1201_ (.A(_0752_),
    .B(\mem[5][15] ),
    .C(_0753_),
    .X(_0083_));
 sky130_fd_sc_hd__a31oi_1 _1202_ (.A1(_0751_),
    .A2(\mem[2][15] ),
    .A3(_0683_),
    .B1(_0083_),
    .Y(_0084_));
 sky130_fd_sc_hd__o22ai_1 _1203_ (.A1(_0665_),
    .A2(_0082_),
    .B1(_0084_),
    .B2(_0664_),
    .Y(_0085_));
 sky130_fd_sc_hd__buf_4 _1204_ (.A(_0759_),
    .X(_0086_));
 sky130_fd_sc_hd__a22oi_1 _1205_ (.A1(\mem[8][15] ),
    .A2(_0086_),
    .B1(_0675_),
    .B2(\mem[9][15] ),
    .Y(_0087_));
 sky130_fd_sc_hd__nand2_1 _1206_ (.A(\mem[15][15] ),
    .B(_0764_),
    .Y(_0088_));
 sky130_fd_sc_hd__o21ai_0 _1207_ (.A1(_0758_),
    .A2(_0087_),
    .B1(_0088_),
    .Y(_0089_));
 sky130_fd_sc_hd__a2111oi_0 _1208_ (.A1(_0079_),
    .A2(_0080_),
    .B1(_0727_),
    .C1(_0085_),
    .D1(_0089_),
    .Y(_0090_));
 sky130_fd_sc_hd__nor2_1 _1209_ (.A(\mem[0][15] ),
    .B(_0729_),
    .Y(_0091_));
 sky130_fd_sc_hd__nand2_1 _1210_ (.A(net51),
    .B(_0731_),
    .Y(_0092_));
 sky130_fd_sc_hd__o31ai_1 _1211_ (.A1(_0702_),
    .A2(_0090_),
    .A3(_0091_),
    .B1(_0092_),
    .Y(_0026_));
 sky130_fd_sc_hd__a22oi_1 _1212_ (.A1(_0698_),
    .A2(\mem[15][16] ),
    .B1(\mem[14][16] ),
    .B2(_0647_),
    .Y(_0093_));
 sky130_fd_sc_hd__a221oi_1 _1213_ (.A1(_0698_),
    .A2(\mem[7][16] ),
    .B1(\mem[6][16] ),
    .B2(_0706_),
    .C1(_0663_),
    .Y(_0094_));
 sky130_fd_sc_hd__a21oi_1 _1214_ (.A1(_0660_),
    .A2(_0093_),
    .B1(_0094_),
    .Y(_0095_));
 sky130_fd_sc_hd__a221oi_1 _1215_ (.A1(\mem[12][16] ),
    .A2(_0709_),
    .B1(_0710_),
    .B2(\mem[13][16] ),
    .C1(_0713_),
    .Y(_0096_));
 sky130_fd_sc_hd__a221oi_1 _1216_ (.A1(\mem[4][16] ),
    .A2(_0709_),
    .B1(_0710_),
    .B2(\mem[5][16] ),
    .C1(_0715_),
    .Y(_0097_));
 sky130_fd_sc_hd__a22oi_1 _1217_ (.A1(\mem[10][16] ),
    .A2(_0646_),
    .B1(_0717_),
    .B2(\mem[9][16] ),
    .Y(_0098_));
 sky130_fd_sc_hd__a22oi_1 _1218_ (.A1(_0719_),
    .A2(\mem[3][16] ),
    .B1(\mem[2][16] ),
    .B2(_0666_),
    .Y(_0099_));
 sky130_fd_sc_hd__a22o_1 _1219_ (.A1(_0696_),
    .A2(_0098_),
    .B1(_0099_),
    .B2(_0721_),
    .X(_0100_));
 sky130_fd_sc_hd__nor3_1 _1220_ (.A(_0096_),
    .B(_0097_),
    .C(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hd__a32oi_1 _1221_ (.A1(_0682_),
    .A2(\mem[1][16] ),
    .A3(_0652_),
    .B1(_0686_),
    .B2(\mem[11][16] ),
    .Y(_0102_));
 sky130_fd_sc_hd__nand3_1 _1222_ (.A(_0660_),
    .B(\mem[8][16] ),
    .C(_0670_),
    .Y(_0103_));
 sky130_fd_sc_hd__a21oi_1 _1223_ (.A1(_0102_),
    .A2(_0103_),
    .B1(_0673_),
    .Y(_0104_));
 sky130_fd_sc_hd__a2111oi_0 _1224_ (.A1(_0704_),
    .A2(_0095_),
    .B1(_0101_),
    .C1(_0104_),
    .D1(_0727_),
    .Y(_0105_));
 sky130_fd_sc_hd__nor2_1 _1225_ (.A(\mem[0][16] ),
    .B(_0729_),
    .Y(_0106_));
 sky130_fd_sc_hd__nand2_1 _1226_ (.A(net52),
    .B(_0731_),
    .Y(_0107_));
 sky130_fd_sc_hd__o31ai_1 _1227_ (.A1(_0702_),
    .A2(_0105_),
    .A3(_0106_),
    .B1(_0107_),
    .Y(_0027_));
 sky130_fd_sc_hd__a21oi_1 _1228_ (.A1(\mem[3][17] ),
    .A2(_0733_),
    .B1(_0734_),
    .Y(_0108_));
 sky130_fd_sc_hd__a222oi_1 _1229_ (.A1(_0736_),
    .A2(\mem[7][17] ),
    .B1(\mem[4][17] ),
    .B2(_0669_),
    .C1(_0737_),
    .C2(\mem[6][17] ),
    .Y(_0109_));
 sky130_fd_sc_hd__a21oi_1 _1230_ (.A1(\mem[10][17] ),
    .A2(_0741_),
    .B1(_0742_),
    .Y(_0110_));
 sky130_fd_sc_hd__a222oi_1 _1231_ (.A1(\mem[14][17] ),
    .A2(_0077_),
    .B1(_0744_),
    .B2(\mem[13][17] ),
    .C1(\mem[12][17] ),
    .C2(_0651_),
    .Y(_0111_));
 sky130_fd_sc_hd__a22oi_1 _1232_ (.A1(_0108_),
    .A2(_0109_),
    .B1(_0110_),
    .B2(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__o21ai_0 _1233_ (.A1(_0108_),
    .A2(_0110_),
    .B1(_0867_),
    .Y(_0113_));
 sky130_fd_sc_hd__a32oi_1 _1234_ (.A1(_0081_),
    .A2(\mem[1][17] ),
    .A3(_0652_),
    .B1(_0749_),
    .B2(\mem[11][17] ),
    .Y(_0114_));
 sky130_fd_sc_hd__and3_1 _1235_ (.A(_0752_),
    .B(\mem[5][17] ),
    .C(_0753_),
    .X(_0115_));
 sky130_fd_sc_hd__a31oi_1 _1236_ (.A1(_0751_),
    .A2(\mem[2][17] ),
    .A3(_0683_),
    .B1(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__o22ai_1 _1237_ (.A1(_0665_),
    .A2(_0114_),
    .B1(_0116_),
    .B2(_0664_),
    .Y(_0117_));
 sky130_fd_sc_hd__a22oi_1 _1238_ (.A1(\mem[8][17] ),
    .A2(_0086_),
    .B1(_0675_),
    .B2(\mem[9][17] ),
    .Y(_0118_));
 sky130_fd_sc_hd__nand2_1 _1239_ (.A(\mem[15][17] ),
    .B(_0764_),
    .Y(_0119_));
 sky130_fd_sc_hd__o21ai_0 _1240_ (.A1(_0758_),
    .A2(_0118_),
    .B1(_0119_),
    .Y(_0120_));
 sky130_fd_sc_hd__a2111oi_0 _1241_ (.A1(_0112_),
    .A2(_0113_),
    .B1(_0727_),
    .C1(_0117_),
    .D1(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hd__nor2_1 _1242_ (.A(\mem[0][17] ),
    .B(_0729_),
    .Y(_0122_));
 sky130_fd_sc_hd__nand2_1 _1243_ (.A(net53),
    .B(_0731_),
    .Y(_0123_));
 sky130_fd_sc_hd__o31ai_1 _1244_ (.A1(_0702_),
    .A2(_0121_),
    .A3(_0122_),
    .B1(_0123_),
    .Y(_0028_));
 sky130_fd_sc_hd__a22oi_1 _1245_ (.A1(_0698_),
    .A2(\mem[15][18] ),
    .B1(\mem[14][18] ),
    .B2(_0647_),
    .Y(_0124_));
 sky130_fd_sc_hd__a221oi_1 _1246_ (.A1(_0698_),
    .A2(\mem[7][18] ),
    .B1(\mem[6][18] ),
    .B2(_0706_),
    .C1(_0663_),
    .Y(_0125_));
 sky130_fd_sc_hd__a21oi_1 _1247_ (.A1(_0660_),
    .A2(_0124_),
    .B1(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__a221oi_1 _1248_ (.A1(\mem[12][18] ),
    .A2(_0709_),
    .B1(_0710_),
    .B2(\mem[13][18] ),
    .C1(_0713_),
    .Y(_0127_));
 sky130_fd_sc_hd__a221oi_1 _1249_ (.A1(\mem[4][18] ),
    .A2(_0709_),
    .B1(_0710_),
    .B2(\mem[5][18] ),
    .C1(_0715_),
    .Y(_0128_));
 sky130_fd_sc_hd__a22oi_1 _1250_ (.A1(\mem[10][18] ),
    .A2(_0646_),
    .B1(_0717_),
    .B2(\mem[9][18] ),
    .Y(_0129_));
 sky130_fd_sc_hd__a22oi_1 _1251_ (.A1(_0637_),
    .A2(\mem[3][18] ),
    .B1(\mem[2][18] ),
    .B2(_0666_),
    .Y(_0130_));
 sky130_fd_sc_hd__a22o_1 _1252_ (.A1(_0696_),
    .A2(_0129_),
    .B1(_0130_),
    .B2(_0721_),
    .X(_0131_));
 sky130_fd_sc_hd__nor3_1 _1253_ (.A(_0127_),
    .B(_0128_),
    .C(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__a32oi_1 _1254_ (.A1(_0682_),
    .A2(\mem[1][18] ),
    .A3(_0652_),
    .B1(_0686_),
    .B2(\mem[11][18] ),
    .Y(_0133_));
 sky130_fd_sc_hd__nand3_1 _1255_ (.A(_0811_),
    .B(\mem[8][18] ),
    .C(_0670_),
    .Y(_0134_));
 sky130_fd_sc_hd__a21oi_1 _1256_ (.A1(_0133_),
    .A2(_0134_),
    .B1(_0673_),
    .Y(_0135_));
 sky130_fd_sc_hd__a2111oi_0 _1257_ (.A1(_0704_),
    .A2(_0126_),
    .B1(_0132_),
    .C1(_0135_),
    .D1(_0727_),
    .Y(_0136_));
 sky130_fd_sc_hd__nor2_1 _1258_ (.A(\mem[0][18] ),
    .B(_0729_),
    .Y(_0137_));
 sky130_fd_sc_hd__nand2_1 _1259_ (.A(net54),
    .B(_0731_),
    .Y(_0138_));
 sky130_fd_sc_hd__o31ai_1 _1260_ (.A1(_0702_),
    .A2(_0136_),
    .A3(_0137_),
    .B1(_0138_),
    .Y(_0029_));
 sky130_fd_sc_hd__a21oi_1 _1261_ (.A1(\mem[3][19] ),
    .A2(_0733_),
    .B1(_0734_),
    .Y(_0139_));
 sky130_fd_sc_hd__a222oi_1 _1262_ (.A1(_0736_),
    .A2(\mem[7][19] ),
    .B1(\mem[4][19] ),
    .B2(_0669_),
    .C1(_0737_),
    .C2(\mem[6][19] ),
    .Y(_0140_));
 sky130_fd_sc_hd__a21oi_1 _1263_ (.A1(\mem[10][19] ),
    .A2(_0741_),
    .B1(_0742_),
    .Y(_0141_));
 sky130_fd_sc_hd__a222oi_1 _1264_ (.A1(\mem[14][19] ),
    .A2(_0077_),
    .B1(_0744_),
    .B2(\mem[13][19] ),
    .C1(\mem[12][19] ),
    .C2(_0651_),
    .Y(_0142_));
 sky130_fd_sc_hd__a22oi_1 _1265_ (.A1(_0139_),
    .A2(_0140_),
    .B1(_0141_),
    .B2(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__o21ai_0 _1266_ (.A1(_0139_),
    .A2(_0141_),
    .B1(_0867_),
    .Y(_0144_));
 sky130_fd_sc_hd__clkbuf_4 _1267_ (.A(_0638_),
    .X(_0145_));
 sky130_fd_sc_hd__a32oi_1 _1268_ (.A1(_0081_),
    .A2(\mem[1][19] ),
    .A3(_0145_),
    .B1(_0749_),
    .B2(\mem[11][19] ),
    .Y(_0146_));
 sky130_fd_sc_hd__clkbuf_4 _1269_ (.A(_0648_),
    .X(_0147_));
 sky130_fd_sc_hd__and3_1 _1270_ (.A(_0147_),
    .B(\mem[5][19] ),
    .C(_0753_),
    .X(_0148_));
 sky130_fd_sc_hd__a31oi_1 _1271_ (.A1(_0751_),
    .A2(\mem[2][19] ),
    .A3(_0683_),
    .B1(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__o22ai_1 _1272_ (.A1(_0665_),
    .A2(_0146_),
    .B1(_0149_),
    .B2(_0664_),
    .Y(_0150_));
 sky130_fd_sc_hd__a22oi_1 _1273_ (.A1(\mem[8][19] ),
    .A2(_0086_),
    .B1(_0675_),
    .B2(\mem[9][19] ),
    .Y(_0151_));
 sky130_fd_sc_hd__nand2_1 _1274_ (.A(\mem[15][19] ),
    .B(_0764_),
    .Y(_0152_));
 sky130_fd_sc_hd__o21ai_0 _1275_ (.A1(_0758_),
    .A2(_0151_),
    .B1(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__a2111oi_1 _1276_ (.A1(_0143_),
    .A2(_0144_),
    .B1(_0727_),
    .C1(_0150_),
    .D1(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__nor2_1 _1277_ (.A(\mem[0][19] ),
    .B(_0729_),
    .Y(_0155_));
 sky130_fd_sc_hd__nand2_1 _1278_ (.A(net55),
    .B(_0731_),
    .Y(_0156_));
 sky130_fd_sc_hd__o31ai_1 _1279_ (.A1(_0702_),
    .A2(_0154_),
    .A3(_0155_),
    .B1(_0156_),
    .Y(_0030_));
 sky130_fd_sc_hd__buf_6 _1280_ (.A(_0632_),
    .X(_0157_));
 sky130_fd_sc_hd__a21oi_1 _1281_ (.A1(\mem[3][1] ),
    .A2(_0733_),
    .B1(_0734_),
    .Y(_0158_));
 sky130_fd_sc_hd__a222oi_1 _1282_ (.A1(_0736_),
    .A2(\mem[7][1] ),
    .B1(\mem[4][1] ),
    .B2(_0669_),
    .C1(_0737_),
    .C2(\mem[6][1] ),
    .Y(_0159_));
 sky130_fd_sc_hd__a21oi_1 _1283_ (.A1(\mem[10][1] ),
    .A2(_0741_),
    .B1(_0742_),
    .Y(_0160_));
 sky130_fd_sc_hd__clkbuf_4 _1284_ (.A(_0634_),
    .X(_0161_));
 sky130_fd_sc_hd__buf_6 _1285_ (.A(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__a222oi_1 _1286_ (.A1(\mem[14][1] ),
    .A2(_0077_),
    .B1(_0744_),
    .B2(\mem[13][1] ),
    .C1(\mem[12][1] ),
    .C2(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__a22oi_1 _1287_ (.A1(_0158_),
    .A2(_0159_),
    .B1(_0160_),
    .B2(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__o21ai_0 _1288_ (.A1(_0158_),
    .A2(_0160_),
    .B1(_0867_),
    .Y(_0165_));
 sky130_fd_sc_hd__clkbuf_4 _1289_ (.A(_0685_),
    .X(_0166_));
 sky130_fd_sc_hd__a32oi_1 _1290_ (.A1(_0081_),
    .A2(\mem[1][1] ),
    .A3(_0145_),
    .B1(_0166_),
    .B2(\mem[11][1] ),
    .Y(_0167_));
 sky130_fd_sc_hd__clkbuf_4 _1291_ (.A(_0666_),
    .X(_0168_));
 sky130_fd_sc_hd__and3_1 _1292_ (.A(_0147_),
    .B(\mem[5][1] ),
    .C(_0753_),
    .X(_0169_));
 sky130_fd_sc_hd__a31oi_1 _1293_ (.A1(_0751_),
    .A2(\mem[2][1] ),
    .A3(_0168_),
    .B1(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__o22ai_2 _1294_ (.A1(_0665_),
    .A2(_0167_),
    .B1(_0170_),
    .B2(_0664_),
    .Y(_0171_));
 sky130_fd_sc_hd__a22oi_1 _1295_ (.A1(\mem[8][1] ),
    .A2(_0086_),
    .B1(_0675_),
    .B2(\mem[9][1] ),
    .Y(_0172_));
 sky130_fd_sc_hd__nand2_1 _1296_ (.A(\mem[15][1] ),
    .B(_0764_),
    .Y(_0173_));
 sky130_fd_sc_hd__o21ai_0 _1297_ (.A1(_0758_),
    .A2(_0172_),
    .B1(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__a2111oi_2 _1298_ (.A1(_0164_),
    .A2(_0165_),
    .B1(_0727_),
    .C1(_0171_),
    .D1(_0174_),
    .Y(_0175_));
 sky130_fd_sc_hd__buf_6 _1299_ (.A(_0641_),
    .X(_0176_));
 sky130_fd_sc_hd__nor2_1 _1300_ (.A(\mem[0][1] ),
    .B(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__buf_6 _1301_ (.A(_0633_),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _1302_ (.A(net56),
    .B(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__o31ai_1 _1303_ (.A1(_0157_),
    .A2(_0175_),
    .A3(_0177_),
    .B1(_0179_),
    .Y(_0031_));
 sky130_fd_sc_hd__a32o_1 _1304_ (.A1(_0682_),
    .A2(\mem[6][20] ),
    .A3(_0647_),
    .B1(_0686_),
    .B2(\mem[15][20] ),
    .X(_0180_));
 sky130_fd_sc_hd__nand3_1 _1305_ (.A(_0811_),
    .B(\mem[8][20] ),
    .C(_0670_),
    .Y(_0181_));
 sky130_fd_sc_hd__nand3_1 _1306_ (.A(_0863_),
    .B(\mem[1][20] ),
    .C(_0814_),
    .Y(_0182_));
 sky130_fd_sc_hd__a21oi_1 _1307_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_0816_),
    .Y(_0183_));
 sky130_fd_sc_hd__nand3_1 _1308_ (.A(_0783_),
    .B(\mem[13][20] ),
    .C(_0818_),
    .Y(_0184_));
 sky130_fd_sc_hd__nand3_1 _1309_ (.A(_0820_),
    .B(\mem[10][20] ),
    .C(_0667_),
    .Y(_0185_));
 sky130_fd_sc_hd__and3_1 _1310_ (.A(_0822_),
    .B(\mem[4][20] ),
    .C(_0161_),
    .X(_0186_));
 sky130_fd_sc_hd__a211oi_1 _1311_ (.A1(\mem[3][20] ),
    .A2(_0658_),
    .B1(_0186_),
    .C1(_0825_),
    .Y(_0187_));
 sky130_fd_sc_hd__a31oi_1 _1312_ (.A1(_0688_),
    .A2(_0184_),
    .A3(_0185_),
    .B1(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__a22oi_2 _1313_ (.A1(\mem[7][20] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][20] ),
    .Y(_0189_));
 sky130_fd_sc_hd__and3_1 _1314_ (.A(_0711_),
    .B(_0833_),
    .C(\mem[14][20] ),
    .X(_0190_));
 sky130_fd_sc_hd__nor3b_1 _1315_ (.A(_0770_),
    .B(_0654_),
    .C_N(\mem[2][20] ),
    .Y(_0191_));
 sky130_fd_sc_hd__o21ai_2 _1316_ (.A1(_0190_),
    .A2(_0191_),
    .B1(_0678_),
    .Y(_0192_));
 sky130_fd_sc_hd__a22oi_2 _1317_ (.A1(_0636_),
    .A2(_0640_),
    .B1(_0694_),
    .B2(\mem[5][20] ),
    .Y(_0193_));
 sky130_fd_sc_hd__and3_1 _1318_ (.A(_0703_),
    .B(\mem[12][20] ),
    .C(_0823_),
    .X(_0194_));
 sky130_fd_sc_hd__and3b_1 _1319_ (.A_N(_0712_),
    .B(\mem[9][20] ),
    .C(_0674_),
    .X(_0195_));
 sky130_fd_sc_hd__o21ai_2 _1320_ (.A1(_0194_),
    .A2(_0195_),
    .B1(_0645_),
    .Y(_0196_));
 sky130_fd_sc_hd__o2111ai_4 _1321_ (.A1(_0829_),
    .A2(_0189_),
    .B1(_0192_),
    .C1(_0193_),
    .D1(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__a2111oi_1 _1322_ (.A1(_0704_),
    .A2(_0180_),
    .B1(_0183_),
    .C1(_0188_),
    .D1(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__nor2_1 _1323_ (.A(\mem[0][20] ),
    .B(_0176_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand2_1 _1324_ (.A(net57),
    .B(_0178_),
    .Y(_0200_));
 sky130_fd_sc_hd__o31ai_1 _1325_ (.A1(_0157_),
    .A2(_0198_),
    .A3(_0199_),
    .B1(_0200_),
    .Y(_0032_));
 sky130_fd_sc_hd__a21oi_1 _1326_ (.A1(\mem[3][21] ),
    .A2(_0733_),
    .B1(_0734_),
    .Y(_0201_));
 sky130_fd_sc_hd__a222oi_1 _1327_ (.A1(_0736_),
    .A2(\mem[7][21] ),
    .B1(\mem[4][21] ),
    .B2(_0669_),
    .C1(_0737_),
    .C2(\mem[6][21] ),
    .Y(_0202_));
 sky130_fd_sc_hd__buf_4 _1328_ (.A(_0630_),
    .X(_0203_));
 sky130_fd_sc_hd__a21oi_1 _1329_ (.A1(\mem[10][21] ),
    .A2(_0741_),
    .B1(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__a222oi_1 _1330_ (.A1(\mem[14][21] ),
    .A2(_0077_),
    .B1(_0744_),
    .B2(\mem[13][21] ),
    .C1(\mem[12][21] ),
    .C2(_0162_),
    .Y(_0205_));
 sky130_fd_sc_hd__a22oi_1 _1331_ (.A1(_0201_),
    .A2(_0202_),
    .B1(_0204_),
    .B2(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__buf_4 _1332_ (.A(_0628_),
    .X(_0207_));
 sky130_fd_sc_hd__o21ai_0 _1333_ (.A1(_0201_),
    .A2(_0204_),
    .B1(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__buf_4 _1334_ (.A(_0699_),
    .X(_0209_));
 sky130_fd_sc_hd__a32oi_1 _1335_ (.A1(_0081_),
    .A2(\mem[1][21] ),
    .A3(_0145_),
    .B1(_0166_),
    .B2(\mem[11][21] ),
    .Y(_0210_));
 sky130_fd_sc_hd__and3_1 _1336_ (.A(_0147_),
    .B(\mem[5][21] ),
    .C(_0753_),
    .X(_0211_));
 sky130_fd_sc_hd__a31oi_1 _1337_ (.A1(_0751_),
    .A2(\mem[2][21] ),
    .A3(_0168_),
    .B1(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__buf_4 _1338_ (.A(_0663_),
    .X(_0213_));
 sky130_fd_sc_hd__o22ai_1 _1339_ (.A1(_0665_),
    .A2(_0210_),
    .B1(_0212_),
    .B2(_0213_),
    .Y(_0214_));
 sky130_fd_sc_hd__buf_4 _1340_ (.A(_0674_),
    .X(_0215_));
 sky130_fd_sc_hd__a22oi_1 _1341_ (.A1(\mem[8][21] ),
    .A2(_0086_),
    .B1(_0215_),
    .B2(\mem[9][21] ),
    .Y(_0216_));
 sky130_fd_sc_hd__nand2_1 _1342_ (.A(\mem[15][21] ),
    .B(_0764_),
    .Y(_0217_));
 sky130_fd_sc_hd__o21ai_0 _1343_ (.A1(_0758_),
    .A2(_0216_),
    .B1(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__a2111oi_1 _1344_ (.A1(_0206_),
    .A2(_0208_),
    .B1(_0209_),
    .C1(_0214_),
    .D1(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__nor2_1 _1345_ (.A(\mem[0][21] ),
    .B(_0176_),
    .Y(_0220_));
 sky130_fd_sc_hd__nand2_1 _1346_ (.A(net58),
    .B(_0178_),
    .Y(_0221_));
 sky130_fd_sc_hd__o31ai_1 _1347_ (.A1(_0157_),
    .A2(_0219_),
    .A3(_0220_),
    .B1(_0221_),
    .Y(_0033_));
 sky130_fd_sc_hd__a32o_1 _1348_ (.A1(_0748_),
    .A2(\mem[6][22] ),
    .A3(_0647_),
    .B1(_0686_),
    .B2(\mem[15][22] ),
    .X(_0222_));
 sky130_fd_sc_hd__nand3_1 _1349_ (.A(_0811_),
    .B(\mem[8][22] ),
    .C(_0670_),
    .Y(_0223_));
 sky130_fd_sc_hd__nand3_1 _1350_ (.A(_0863_),
    .B(\mem[1][22] ),
    .C(_0814_),
    .Y(_0224_));
 sky130_fd_sc_hd__a21oi_1 _1351_ (.A1(_0223_),
    .A2(_0224_),
    .B1(_0816_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand3_1 _1352_ (.A(_0783_),
    .B(\mem[13][22] ),
    .C(_0818_),
    .Y(_0226_));
 sky130_fd_sc_hd__nand3_1 _1353_ (.A(_0820_),
    .B(\mem[10][22] ),
    .C(_0667_),
    .Y(_0227_));
 sky130_fd_sc_hd__and3_1 _1354_ (.A(_0822_),
    .B(\mem[4][22] ),
    .C(_0161_),
    .X(_0228_));
 sky130_fd_sc_hd__a211oi_1 _1355_ (.A1(\mem[3][22] ),
    .A2(_0658_),
    .B1(_0228_),
    .C1(_0825_),
    .Y(_0229_));
 sky130_fd_sc_hd__a31oi_1 _1356_ (.A1(_0688_),
    .A2(_0226_),
    .A3(_0227_),
    .B1(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__a22oi_2 _1357_ (.A1(\mem[7][22] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][22] ),
    .Y(_0231_));
 sky130_fd_sc_hd__and3_1 _1358_ (.A(_0711_),
    .B(_0833_),
    .C(\mem[14][22] ),
    .X(_0232_));
 sky130_fd_sc_hd__nor3b_1 _1359_ (.A(_0659_),
    .B(_0654_),
    .C_N(\mem[2][22] ),
    .Y(_0233_));
 sky130_fd_sc_hd__o21ai_1 _1360_ (.A1(_0232_),
    .A2(_0233_),
    .B1(_0678_),
    .Y(_0234_));
 sky130_fd_sc_hd__a22oi_2 _1361_ (.A1(_0636_),
    .A2(_0640_),
    .B1(_0694_),
    .B2(\mem[5][22] ),
    .Y(_0235_));
 sky130_fd_sc_hd__and3_1 _1362_ (.A(_0703_),
    .B(\mem[12][22] ),
    .C(_0823_),
    .X(_0236_));
 sky130_fd_sc_hd__and3b_1 _1363_ (.A_N(_0712_),
    .B(\mem[9][22] ),
    .C(_0813_),
    .X(_0237_));
 sky130_fd_sc_hd__o21ai_1 _1364_ (.A1(_0236_),
    .A2(_0237_),
    .B1(_0645_),
    .Y(_0238_));
 sky130_fd_sc_hd__o2111ai_4 _1365_ (.A1(_0829_),
    .A2(_0231_),
    .B1(_0234_),
    .C1(_0235_),
    .D1(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__a2111oi_1 _1366_ (.A1(_0704_),
    .A2(_0222_),
    .B1(_0225_),
    .C1(_0230_),
    .D1(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__nor2_1 _1367_ (.A(\mem[0][22] ),
    .B(_0176_),
    .Y(_0241_));
 sky130_fd_sc_hd__nand2_1 _1368_ (.A(net59),
    .B(_0178_),
    .Y(_0242_));
 sky130_fd_sc_hd__o31ai_1 _1369_ (.A1(_0157_),
    .A2(_0240_),
    .A3(_0241_),
    .B1(_0242_),
    .Y(_0034_));
 sky130_fd_sc_hd__a21oi_1 _1370_ (.A1(\mem[3][23] ),
    .A2(_0733_),
    .B1(_0734_),
    .Y(_0243_));
 sky130_fd_sc_hd__a222oi_1 _1371_ (.A1(_0736_),
    .A2(\mem[7][23] ),
    .B1(\mem[4][23] ),
    .B2(_0669_),
    .C1(_0737_),
    .C2(\mem[6][23] ),
    .Y(_0244_));
 sky130_fd_sc_hd__a21oi_1 _1372_ (.A1(\mem[10][23] ),
    .A2(_0741_),
    .B1(_0203_),
    .Y(_0245_));
 sky130_fd_sc_hd__a222oi_1 _1373_ (.A1(\mem[14][23] ),
    .A2(_0077_),
    .B1(_0744_),
    .B2(\mem[13][23] ),
    .C1(\mem[12][23] ),
    .C2(_0162_),
    .Y(_0246_));
 sky130_fd_sc_hd__a22oi_1 _1374_ (.A1(_0243_),
    .A2(_0244_),
    .B1(_0245_),
    .B2(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__o21ai_0 _1375_ (.A1(_0243_),
    .A2(_0245_),
    .B1(_0207_),
    .Y(_0248_));
 sky130_fd_sc_hd__a32oi_1 _1376_ (.A1(_0081_),
    .A2(\mem[1][23] ),
    .A3(_0145_),
    .B1(_0166_),
    .B2(\mem[11][23] ),
    .Y(_0249_));
 sky130_fd_sc_hd__and3_1 _1377_ (.A(_0147_),
    .B(\mem[5][23] ),
    .C(_0753_),
    .X(_0250_));
 sky130_fd_sc_hd__a31oi_1 _1378_ (.A1(_0751_),
    .A2(\mem[2][23] ),
    .A3(_0168_),
    .B1(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__o22ai_1 _1379_ (.A1(_0655_),
    .A2(_0249_),
    .B1(_0251_),
    .B2(_0213_),
    .Y(_0252_));
 sky130_fd_sc_hd__a22oi_1 _1380_ (.A1(\mem[8][23] ),
    .A2(_0086_),
    .B1(_0215_),
    .B2(\mem[9][23] ),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_1 _1381_ (.A(\mem[15][23] ),
    .B(_0763_),
    .Y(_0254_));
 sky130_fd_sc_hd__o21ai_0 _1382_ (.A1(_0758_),
    .A2(_0253_),
    .B1(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__a2111oi_1 _1383_ (.A1(_0247_),
    .A2(_0248_),
    .B1(_0209_),
    .C1(_0252_),
    .D1(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__nor2_1 _1384_ (.A(\mem[0][23] ),
    .B(_0176_),
    .Y(_0257_));
 sky130_fd_sc_hd__nand2_1 _1385_ (.A(net60),
    .B(_0178_),
    .Y(_0258_));
 sky130_fd_sc_hd__o31ai_1 _1386_ (.A1(_0157_),
    .A2(_0256_),
    .A3(_0257_),
    .B1(_0258_),
    .Y(_0035_));
 sky130_fd_sc_hd__a32o_1 _1387_ (.A1(_0748_),
    .A2(\mem[6][24] ),
    .A3(_0647_),
    .B1(_0686_),
    .B2(\mem[15][24] ),
    .X(_0259_));
 sky130_fd_sc_hd__nand3_1 _1388_ (.A(_0811_),
    .B(\mem[8][24] ),
    .C(_0760_),
    .Y(_0260_));
 sky130_fd_sc_hd__nand3_1 _1389_ (.A(_0863_),
    .B(\mem[1][24] ),
    .C(_0814_),
    .Y(_0261_));
 sky130_fd_sc_hd__a21oi_1 _1390_ (.A1(_0260_),
    .A2(_0261_),
    .B1(_0816_),
    .Y(_0262_));
 sky130_fd_sc_hd__nand3_1 _1391_ (.A(_0783_),
    .B(\mem[13][24] ),
    .C(_0818_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand3_1 _1392_ (.A(_0820_),
    .B(\mem[10][24] ),
    .C(_0667_),
    .Y(_0264_));
 sky130_fd_sc_hd__and3_1 _1393_ (.A(_0822_),
    .B(\mem[4][24] ),
    .C(_0161_),
    .X(_0265_));
 sky130_fd_sc_hd__a211oi_1 _1394_ (.A1(\mem[3][24] ),
    .A2(_0658_),
    .B1(_0265_),
    .C1(_0825_),
    .Y(_0266_));
 sky130_fd_sc_hd__a31oi_1 _1395_ (.A1(_0688_),
    .A2(_0263_),
    .A3(_0264_),
    .B1(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__a22oi_2 _1396_ (.A1(\mem[7][24] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][24] ),
    .Y(_0268_));
 sky130_fd_sc_hd__and3_1 _1397_ (.A(_0711_),
    .B(_0833_),
    .C(\mem[14][24] ),
    .X(_0269_));
 sky130_fd_sc_hd__nor3b_1 _1398_ (.A(_0659_),
    .B(_0654_),
    .C_N(\mem[2][24] ),
    .Y(_0270_));
 sky130_fd_sc_hd__o21ai_1 _1399_ (.A1(_0269_),
    .A2(_0270_),
    .B1(_0678_),
    .Y(_0271_));
 sky130_fd_sc_hd__a22oi_2 _1400_ (.A1(_0636_),
    .A2(_0640_),
    .B1(_0694_),
    .B2(\mem[5][24] ),
    .Y(_0272_));
 sky130_fd_sc_hd__and3_1 _1401_ (.A(_0703_),
    .B(\mem[12][24] ),
    .C(_0823_),
    .X(_0273_));
 sky130_fd_sc_hd__and3b_1 _1402_ (.A_N(_0712_),
    .B(\mem[9][24] ),
    .C(_0813_),
    .X(_0274_));
 sky130_fd_sc_hd__o21ai_1 _1403_ (.A1(_0273_),
    .A2(_0274_),
    .B1(_0645_),
    .Y(_0275_));
 sky130_fd_sc_hd__o2111ai_4 _1404_ (.A1(_0829_),
    .A2(_0268_),
    .B1(_0271_),
    .C1(_0272_),
    .D1(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__a2111oi_1 _1405_ (.A1(_0704_),
    .A2(_0259_),
    .B1(_0262_),
    .C1(_0267_),
    .D1(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__nor2_1 _1406_ (.A(\mem[0][24] ),
    .B(_0176_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand2_1 _1407_ (.A(net61),
    .B(_0178_),
    .Y(_0279_));
 sky130_fd_sc_hd__o31ai_1 _1408_ (.A1(_0157_),
    .A2(_0277_),
    .A3(_0278_),
    .B1(_0279_),
    .Y(_0036_));
 sky130_fd_sc_hd__a21oi_1 _1409_ (.A1(\mem[3][25] ),
    .A2(_0657_),
    .B1(_0734_),
    .Y(_0280_));
 sky130_fd_sc_hd__a222oi_1 _1410_ (.A1(_0719_),
    .A2(\mem[7][25] ),
    .B1(\mem[4][25] ),
    .B2(_0669_),
    .C1(_0737_),
    .C2(\mem[6][25] ),
    .Y(_0281_));
 sky130_fd_sc_hd__a21oi_1 _1411_ (.A1(\mem[10][25] ),
    .A2(_0741_),
    .B1(_0203_),
    .Y(_0282_));
 sky130_fd_sc_hd__a222oi_1 _1412_ (.A1(\mem[14][25] ),
    .A2(_0077_),
    .B1(_0744_),
    .B2(\mem[13][25] ),
    .C1(\mem[12][25] ),
    .C2(_0162_),
    .Y(_0283_));
 sky130_fd_sc_hd__a22oi_1 _1413_ (.A1(_0280_),
    .A2(_0281_),
    .B1(_0282_),
    .B2(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_0 _1414_ (.A1(_0280_),
    .A2(_0282_),
    .B1(_0207_),
    .Y(_0285_));
 sky130_fd_sc_hd__a32oi_1 _1415_ (.A1(_0081_),
    .A2(\mem[1][25] ),
    .A3(_0145_),
    .B1(_0166_),
    .B2(\mem[11][25] ),
    .Y(_0286_));
 sky130_fd_sc_hd__and3_1 _1416_ (.A(_0147_),
    .B(\mem[5][25] ),
    .C(_0753_),
    .X(_0287_));
 sky130_fd_sc_hd__a31oi_1 _1417_ (.A1(_0751_),
    .A2(\mem[2][25] ),
    .A3(_0168_),
    .B1(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__o22ai_1 _1418_ (.A1(_0655_),
    .A2(_0286_),
    .B1(_0288_),
    .B2(_0213_),
    .Y(_0289_));
 sky130_fd_sc_hd__a22oi_1 _1419_ (.A1(\mem[8][25] ),
    .A2(_0086_),
    .B1(_0215_),
    .B2(\mem[9][25] ),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_1 _1420_ (.A(\mem[15][25] ),
    .B(_0763_),
    .Y(_0291_));
 sky130_fd_sc_hd__o21ai_0 _1421_ (.A1(_0758_),
    .A2(_0290_),
    .B1(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__a2111oi_1 _1422_ (.A1(_0284_),
    .A2(_0285_),
    .B1(_0209_),
    .C1(_0289_),
    .D1(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__nor2_1 _1423_ (.A(\mem[0][25] ),
    .B(_0176_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _1424_ (.A(net62),
    .B(_0178_),
    .Y(_0295_));
 sky130_fd_sc_hd__o31ai_1 _1425_ (.A1(_0157_),
    .A2(_0293_),
    .A3(_0294_),
    .B1(_0295_),
    .Y(_0037_));
 sky130_fd_sc_hd__a32o_1 _1426_ (.A1(_0748_),
    .A2(\mem[6][26] ),
    .A3(_0706_),
    .B1(_0686_),
    .B2(\mem[15][26] ),
    .X(_0296_));
 sky130_fd_sc_hd__nand3_1 _1427_ (.A(_0811_),
    .B(\mem[8][26] ),
    .C(_0760_),
    .Y(_0297_));
 sky130_fd_sc_hd__nand3_1 _1428_ (.A(_0863_),
    .B(\mem[1][26] ),
    .C(_0814_),
    .Y(_0298_));
 sky130_fd_sc_hd__a21oi_1 _1429_ (.A1(_0297_),
    .A2(_0298_),
    .B1(_0816_),
    .Y(_0299_));
 sky130_fd_sc_hd__nand3_1 _1430_ (.A(_0783_),
    .B(\mem[13][26] ),
    .C(_0818_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand3_1 _1431_ (.A(_0820_),
    .B(\mem[10][26] ),
    .C(_0667_),
    .Y(_0301_));
 sky130_fd_sc_hd__and3_1 _1432_ (.A(_0822_),
    .B(\mem[4][26] ),
    .C(_0161_),
    .X(_0302_));
 sky130_fd_sc_hd__a211oi_1 _1433_ (.A1(\mem[3][26] ),
    .A2(_0658_),
    .B1(_0302_),
    .C1(_0825_),
    .Y(_0303_));
 sky130_fd_sc_hd__a31oi_1 _1434_ (.A1(_0688_),
    .A2(_0300_),
    .A3(_0301_),
    .B1(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__a22oi_2 _1435_ (.A1(\mem[7][26] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][26] ),
    .Y(_0305_));
 sky130_fd_sc_hd__and3_1 _1436_ (.A(_0711_),
    .B(_0833_),
    .C(\mem[14][26] ),
    .X(_0306_));
 sky130_fd_sc_hd__nor3b_1 _1437_ (.A(_0659_),
    .B(_0654_),
    .C_N(\mem[2][26] ),
    .Y(_0307_));
 sky130_fd_sc_hd__o21ai_1 _1438_ (.A1(_0306_),
    .A2(_0307_),
    .B1(_0678_),
    .Y(_0308_));
 sky130_fd_sc_hd__a22oi_2 _1439_ (.A1(_0636_),
    .A2(_0640_),
    .B1(_0694_),
    .B2(\mem[5][26] ),
    .Y(_0309_));
 sky130_fd_sc_hd__and3_1 _1440_ (.A(_0703_),
    .B(\mem[12][26] ),
    .C(_0823_),
    .X(_0310_));
 sky130_fd_sc_hd__and3b_1 _1441_ (.A_N(_0712_),
    .B(\mem[9][26] ),
    .C(_0813_),
    .X(_0311_));
 sky130_fd_sc_hd__o21ai_1 _1442_ (.A1(_0310_),
    .A2(_0311_),
    .B1(_0645_),
    .Y(_0312_));
 sky130_fd_sc_hd__o2111ai_4 _1443_ (.A1(_0829_),
    .A2(_0305_),
    .B1(_0308_),
    .C1(_0309_),
    .D1(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__a2111oi_1 _1444_ (.A1(_0704_),
    .A2(_0296_),
    .B1(_0299_),
    .C1(_0304_),
    .D1(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__nor2_1 _1445_ (.A(\mem[0][26] ),
    .B(_0176_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand2_1 _1446_ (.A(net63),
    .B(_0178_),
    .Y(_0316_));
 sky130_fd_sc_hd__o31ai_1 _1447_ (.A1(_0157_),
    .A2(_0314_),
    .A3(_0315_),
    .B1(_0316_),
    .Y(_0038_));
 sky130_fd_sc_hd__a21oi_1 _1448_ (.A1(\mem[3][27] ),
    .A2(_0657_),
    .B1(_0734_),
    .Y(_0317_));
 sky130_fd_sc_hd__a222oi_1 _1449_ (.A1(_0719_),
    .A2(\mem[7][27] ),
    .B1(\mem[4][27] ),
    .B2(_0759_),
    .C1(_0737_),
    .C2(\mem[6][27] ),
    .Y(_0318_));
 sky130_fd_sc_hd__a21oi_1 _1450_ (.A1(\mem[10][27] ),
    .A2(_0741_),
    .B1(_0203_),
    .Y(_0319_));
 sky130_fd_sc_hd__a222oi_1 _1451_ (.A1(\mem[14][27] ),
    .A2(_0077_),
    .B1(_0744_),
    .B2(\mem[13][27] ),
    .C1(\mem[12][27] ),
    .C2(_0162_),
    .Y(_0320_));
 sky130_fd_sc_hd__a22oi_1 _1452_ (.A1(_0317_),
    .A2(_0318_),
    .B1(_0319_),
    .B2(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__o21ai_0 _1453_ (.A1(_0317_),
    .A2(_0319_),
    .B1(_0207_),
    .Y(_0322_));
 sky130_fd_sc_hd__a32oi_1 _1454_ (.A1(_0081_),
    .A2(\mem[1][27] ),
    .A3(_0145_),
    .B1(_0166_),
    .B2(\mem[11][27] ),
    .Y(_0323_));
 sky130_fd_sc_hd__and3_1 _1455_ (.A(_0147_),
    .B(\mem[5][27] ),
    .C(_0753_),
    .X(_0324_));
 sky130_fd_sc_hd__a31oi_1 _1456_ (.A1(_0751_),
    .A2(\mem[2][27] ),
    .A3(_0168_),
    .B1(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__o22ai_2 _1457_ (.A1(_0655_),
    .A2(_0323_),
    .B1(_0325_),
    .B2(_0213_),
    .Y(_0326_));
 sky130_fd_sc_hd__a22oi_1 _1458_ (.A1(\mem[8][27] ),
    .A2(_0086_),
    .B1(_0215_),
    .B2(\mem[9][27] ),
    .Y(_0327_));
 sky130_fd_sc_hd__nand2_1 _1459_ (.A(\mem[15][27] ),
    .B(_0763_),
    .Y(_0328_));
 sky130_fd_sc_hd__o21ai_1 _1460_ (.A1(_0757_),
    .A2(_0327_),
    .B1(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__a2111oi_2 _1461_ (.A1(_0321_),
    .A2(_0322_),
    .B1(_0209_),
    .C1(_0326_),
    .D1(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__nor2_1 _1462_ (.A(\mem[0][27] ),
    .B(_0176_),
    .Y(_0331_));
 sky130_fd_sc_hd__nand2_1 _1463_ (.A(net64),
    .B(_0178_),
    .Y(_0332_));
 sky130_fd_sc_hd__o31ai_1 _1464_ (.A1(_0157_),
    .A2(_0330_),
    .A3(_0331_),
    .B1(_0332_),
    .Y(_0039_));
 sky130_fd_sc_hd__a32o_1 _1465_ (.A1(_0748_),
    .A2(\mem[6][28] ),
    .A3(_0706_),
    .B1(_0749_),
    .B2(\mem[15][28] ),
    .X(_0333_));
 sky130_fd_sc_hd__nand3_1 _1466_ (.A(_0811_),
    .B(\mem[8][28] ),
    .C(_0760_),
    .Y(_0334_));
 sky130_fd_sc_hd__nand3_1 _1467_ (.A(_0863_),
    .B(\mem[1][28] ),
    .C(_0814_),
    .Y(_0335_));
 sky130_fd_sc_hd__a21oi_1 _1468_ (.A1(_0334_),
    .A2(_0335_),
    .B1(_0816_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand3_1 _1469_ (.A(_0783_),
    .B(\mem[13][28] ),
    .C(_0818_),
    .Y(_0337_));
 sky130_fd_sc_hd__nand3_1 _1470_ (.A(_0820_),
    .B(\mem[10][28] ),
    .C(_0667_),
    .Y(_0338_));
 sky130_fd_sc_hd__and3_1 _1471_ (.A(_0822_),
    .B(\mem[4][28] ),
    .C(_0161_),
    .X(_0339_));
 sky130_fd_sc_hd__a211oi_1 _1472_ (.A1(\mem[3][28] ),
    .A2(_0658_),
    .B1(_0339_),
    .C1(_0825_),
    .Y(_0340_));
 sky130_fd_sc_hd__a31oi_1 _1473_ (.A1(_0688_),
    .A2(_0337_),
    .A3(_0338_),
    .B1(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__a22oi_2 _1474_ (.A1(\mem[7][28] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][28] ),
    .Y(_0342_));
 sky130_fd_sc_hd__and3_1 _1475_ (.A(_0644_),
    .B(_0833_),
    .C(\mem[14][28] ),
    .X(_0343_));
 sky130_fd_sc_hd__nor3b_1 _1476_ (.A(_0659_),
    .B(_0654_),
    .C_N(\mem[2][28] ),
    .Y(_0344_));
 sky130_fd_sc_hd__o21ai_1 _1477_ (.A1(_0343_),
    .A2(_0344_),
    .B1(_0678_),
    .Y(_0345_));
 sky130_fd_sc_hd__a22oi_2 _1478_ (.A1(_0636_),
    .A2(_0640_),
    .B1(_0694_),
    .B2(\mem[5][28] ),
    .Y(_0346_));
 sky130_fd_sc_hd__and3_1 _1479_ (.A(_0752_),
    .B(\mem[12][28] ),
    .C(_0823_),
    .X(_0347_));
 sky130_fd_sc_hd__and3b_1 _1480_ (.A_N(_0712_),
    .B(\mem[9][28] ),
    .C(_0813_),
    .X(_0348_));
 sky130_fd_sc_hd__o21ai_1 _1481_ (.A1(_0347_),
    .A2(_0348_),
    .B1(_0645_),
    .Y(_0349_));
 sky130_fd_sc_hd__o2111ai_4 _1482_ (.A1(_0829_),
    .A2(_0342_),
    .B1(_0345_),
    .C1(_0346_),
    .D1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__a2111oi_2 _1483_ (.A1(_0704_),
    .A2(_0333_),
    .B1(_0336_),
    .C1(_0341_),
    .D1(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__nor2_1 _1484_ (.A(\mem[0][28] ),
    .B(_0176_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _1485_ (.A(net65),
    .B(_0178_),
    .Y(_0353_));
 sky130_fd_sc_hd__o31ai_1 _1486_ (.A1(_0157_),
    .A2(_0351_),
    .A3(_0352_),
    .B1(_0353_),
    .Y(_0040_));
 sky130_fd_sc_hd__buf_6 _1487_ (.A(_0632_),
    .X(_0354_));
 sky130_fd_sc_hd__a21oi_1 _1488_ (.A1(\mem[3][29] ),
    .A2(_0657_),
    .B1(_0770_),
    .Y(_0355_));
 sky130_fd_sc_hd__a222oi_1 _1489_ (.A1(_0719_),
    .A2(\mem[7][29] ),
    .B1(\mem[4][29] ),
    .B2(_0759_),
    .C1(_0677_),
    .C2(\mem[6][29] ),
    .Y(_0356_));
 sky130_fd_sc_hd__a21oi_1 _1490_ (.A1(\mem[10][29] ),
    .A2(_0740_),
    .B1(_0203_),
    .Y(_0357_));
 sky130_fd_sc_hd__a222oi_1 _1491_ (.A1(\mem[14][29] ),
    .A2(_0077_),
    .B1(_0674_),
    .B2(\mem[13][29] ),
    .C1(\mem[12][29] ),
    .C2(_0162_),
    .Y(_0358_));
 sky130_fd_sc_hd__a22oi_1 _1492_ (.A1(_0355_),
    .A2(_0356_),
    .B1(_0357_),
    .B2(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__o21ai_0 _1493_ (.A1(_0355_),
    .A2(_0357_),
    .B1(_0207_),
    .Y(_0360_));
 sky130_fd_sc_hd__a32oi_1 _1494_ (.A1(_0081_),
    .A2(\mem[1][29] ),
    .A3(_0145_),
    .B1(_0166_),
    .B2(\mem[11][29] ),
    .Y(_0361_));
 sky130_fd_sc_hd__and3_1 _1495_ (.A(_0147_),
    .B(\mem[5][29] ),
    .C(_0717_),
    .X(_0362_));
 sky130_fd_sc_hd__a31oi_1 _1496_ (.A1(_0628_),
    .A2(\mem[2][29] ),
    .A3(_0168_),
    .B1(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__o22ai_2 _1497_ (.A1(_0655_),
    .A2(_0361_),
    .B1(_0363_),
    .B2(_0213_),
    .Y(_0364_));
 sky130_fd_sc_hd__a22oi_1 _1498_ (.A1(\mem[8][29] ),
    .A2(_0086_),
    .B1(_0215_),
    .B2(\mem[9][29] ),
    .Y(_0365_));
 sky130_fd_sc_hd__nand2_1 _1499_ (.A(\mem[15][29] ),
    .B(_0763_),
    .Y(_0366_));
 sky130_fd_sc_hd__o21ai_1 _1500_ (.A1(_0757_),
    .A2(_0365_),
    .B1(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__a2111oi_2 _1501_ (.A1(_0359_),
    .A2(_0360_),
    .B1(_0209_),
    .C1(_0364_),
    .D1(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__buf_6 _1502_ (.A(_0641_),
    .X(_0369_));
 sky130_fd_sc_hd__nor2_1 _1503_ (.A(\mem[0][29] ),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__buf_6 _1504_ (.A(_0633_),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_1 _1505_ (.A(net66),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__o31ai_1 _1506_ (.A1(_0354_),
    .A2(_0368_),
    .A3(_0370_),
    .B1(_0372_),
    .Y(_0041_));
 sky130_fd_sc_hd__a32o_1 _1507_ (.A1(_0748_),
    .A2(\mem[6][2] ),
    .A3(_0706_),
    .B1(_0749_),
    .B2(\mem[15][2] ),
    .X(_0373_));
 sky130_fd_sc_hd__nand3_1 _1508_ (.A(_0811_),
    .B(\mem[8][2] ),
    .C(_0760_),
    .Y(_0374_));
 sky130_fd_sc_hd__nand3_1 _1509_ (.A(_0863_),
    .B(\mem[1][2] ),
    .C(_0814_),
    .Y(_0375_));
 sky130_fd_sc_hd__a21oi_1 _1510_ (.A1(_0374_),
    .A2(_0375_),
    .B1(_0816_),
    .Y(_0376_));
 sky130_fd_sc_hd__nand3_1 _1511_ (.A(_0783_),
    .B(\mem[13][2] ),
    .C(_0818_),
    .Y(_0377_));
 sky130_fd_sc_hd__nand3_1 _1512_ (.A(_0820_),
    .B(\mem[10][2] ),
    .C(_0667_),
    .Y(_0378_));
 sky130_fd_sc_hd__and3_1 _1513_ (.A(_0822_),
    .B(\mem[4][2] ),
    .C(_0161_),
    .X(_0379_));
 sky130_fd_sc_hd__a211oi_1 _1514_ (.A1(\mem[3][2] ),
    .A2(_0658_),
    .B1(_0379_),
    .C1(_0825_),
    .Y(_0380_));
 sky130_fd_sc_hd__a31oi_1 _1515_ (.A1(_0688_),
    .A2(_0377_),
    .A3(_0378_),
    .B1(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__a22oi_2 _1516_ (.A1(\mem[7][2] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][2] ),
    .Y(_0382_));
 sky130_fd_sc_hd__and3_1 _1517_ (.A(_0644_),
    .B(_0833_),
    .C(\mem[14][2] ),
    .X(_0383_));
 sky130_fd_sc_hd__nor3b_1 _1518_ (.A(_0659_),
    .B(_0654_),
    .C_N(\mem[2][2] ),
    .Y(_0384_));
 sky130_fd_sc_hd__o21ai_1 _1519_ (.A1(_0383_),
    .A2(_0384_),
    .B1(_0678_),
    .Y(_0385_));
 sky130_fd_sc_hd__a22oi_2 _1520_ (.A1(_0636_),
    .A2(_0640_),
    .B1(_0694_),
    .B2(\mem[5][2] ),
    .Y(_0386_));
 sky130_fd_sc_hd__and3_1 _1521_ (.A(_0752_),
    .B(\mem[12][2] ),
    .C(_0823_),
    .X(_0387_));
 sky130_fd_sc_hd__and3b_1 _1522_ (.A_N(_0712_),
    .B(\mem[9][2] ),
    .C(_0813_),
    .X(_0388_));
 sky130_fd_sc_hd__o21ai_1 _1523_ (.A1(_0387_),
    .A2(_0388_),
    .B1(_0645_),
    .Y(_0389_));
 sky130_fd_sc_hd__o2111ai_4 _1524_ (.A1(_0829_),
    .A2(_0382_),
    .B1(_0385_),
    .C1(_0386_),
    .D1(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__a2111oi_1 _1525_ (.A1(_0704_),
    .A2(_0373_),
    .B1(_0376_),
    .C1(_0381_),
    .D1(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__nor2_1 _1526_ (.A(\mem[0][2] ),
    .B(_0369_),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_1 _1527_ (.A(net67),
    .B(_0371_),
    .Y(_0393_));
 sky130_fd_sc_hd__o31ai_1 _1528_ (.A1(_0354_),
    .A2(_0391_),
    .A3(_0392_),
    .B1(_0393_),
    .Y(_0042_));
 sky130_fd_sc_hd__a22oi_1 _1529_ (.A1(_0698_),
    .A2(\mem[15][30] ),
    .B1(\mem[14][30] ),
    .B2(_0647_),
    .Y(_0394_));
 sky130_fd_sc_hd__a221oi_1 _1530_ (.A1(_0736_),
    .A2(\mem[7][30] ),
    .B1(\mem[6][30] ),
    .B2(_0706_),
    .C1(_0663_),
    .Y(_0395_));
 sky130_fd_sc_hd__a21oi_1 _1531_ (.A1(_0660_),
    .A2(_0394_),
    .B1(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__a221oi_1 _1532_ (.A1(\mem[12][30] ),
    .A2(_0709_),
    .B1(_0710_),
    .B2(\mem[13][30] ),
    .C1(_0713_),
    .Y(_0397_));
 sky130_fd_sc_hd__a221oi_1 _1533_ (.A1(\mem[4][30] ),
    .A2(_0709_),
    .B1(_0710_),
    .B2(\mem[5][30] ),
    .C1(_0715_),
    .Y(_0398_));
 sky130_fd_sc_hd__a22oi_1 _1534_ (.A1(\mem[10][30] ),
    .A2(_0646_),
    .B1(_0717_),
    .B2(\mem[9][30] ),
    .Y(_0399_));
 sky130_fd_sc_hd__a22oi_1 _1535_ (.A1(_0637_),
    .A2(\mem[3][30] ),
    .B1(\mem[2][30] ),
    .B2(_0666_),
    .Y(_0400_));
 sky130_fd_sc_hd__a22o_1 _1536_ (.A1(_0696_),
    .A2(_0399_),
    .B1(_0400_),
    .B2(_0721_),
    .X(_0401_));
 sky130_fd_sc_hd__nor3_1 _1537_ (.A(_0397_),
    .B(_0398_),
    .C(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__a32oi_1 _1538_ (.A1(_0682_),
    .A2(\mem[1][30] ),
    .A3(_0652_),
    .B1(_0686_),
    .B2(\mem[11][30] ),
    .Y(_0403_));
 sky130_fd_sc_hd__nand3_1 _1539_ (.A(_0811_),
    .B(\mem[8][30] ),
    .C(_0670_),
    .Y(_0404_));
 sky130_fd_sc_hd__a21oi_1 _1540_ (.A1(_0403_),
    .A2(_0404_),
    .B1(_0673_),
    .Y(_0405_));
 sky130_fd_sc_hd__a2111oi_1 _1541_ (.A1(_0673_),
    .A2(_0396_),
    .B1(_0402_),
    .C1(_0405_),
    .D1(_0727_),
    .Y(_0406_));
 sky130_fd_sc_hd__nor2_1 _1542_ (.A(\mem[0][30] ),
    .B(_0369_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _1543_ (.A(net68),
    .B(_0371_),
    .Y(_0408_));
 sky130_fd_sc_hd__o31ai_1 _1544_ (.A1(_0354_),
    .A2(_0406_),
    .A3(_0407_),
    .B1(_0408_),
    .Y(_0043_));
 sky130_fd_sc_hd__a21oi_1 _1545_ (.A1(\mem[3][31] ),
    .A2(_0657_),
    .B1(_0770_),
    .Y(_0409_));
 sky130_fd_sc_hd__a222oi_1 _1546_ (.A1(_0719_),
    .A2(\mem[7][31] ),
    .B1(\mem[4][31] ),
    .B2(_0759_),
    .C1(_0677_),
    .C2(\mem[6][31] ),
    .Y(_0410_));
 sky130_fd_sc_hd__a21oi_1 _1547_ (.A1(\mem[10][31] ),
    .A2(_0740_),
    .B1(_0203_),
    .Y(_0411_));
 sky130_fd_sc_hd__a222oi_1 _1548_ (.A1(\mem[14][31] ),
    .A2(_0077_),
    .B1(_0674_),
    .B2(\mem[13][31] ),
    .C1(\mem[12][31] ),
    .C2(_0162_),
    .Y(_0412_));
 sky130_fd_sc_hd__a22oi_1 _1549_ (.A1(_0409_),
    .A2(_0410_),
    .B1(_0411_),
    .B2(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__o21ai_0 _1550_ (.A1(_0409_),
    .A2(_0411_),
    .B1(_0207_),
    .Y(_0414_));
 sky130_fd_sc_hd__a32oi_1 _1551_ (.A1(_0081_),
    .A2(\mem[1][31] ),
    .A3(_0145_),
    .B1(_0166_),
    .B2(\mem[11][31] ),
    .Y(_0415_));
 sky130_fd_sc_hd__and3_1 _1552_ (.A(_0147_),
    .B(\mem[5][31] ),
    .C(_0717_),
    .X(_0416_));
 sky130_fd_sc_hd__a31oi_1 _1553_ (.A1(_0628_),
    .A2(\mem[2][31] ),
    .A3(_0168_),
    .B1(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__o22ai_2 _1554_ (.A1(_0655_),
    .A2(_0415_),
    .B1(_0417_),
    .B2(_0213_),
    .Y(_0418_));
 sky130_fd_sc_hd__a22oi_1 _1555_ (.A1(\mem[8][31] ),
    .A2(_0086_),
    .B1(_0215_),
    .B2(\mem[9][31] ),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _1556_ (.A(\mem[15][31] ),
    .B(_0763_),
    .Y(_0420_));
 sky130_fd_sc_hd__o21ai_1 _1557_ (.A1(_0757_),
    .A2(_0419_),
    .B1(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__a2111oi_2 _1558_ (.A1(_0413_),
    .A2(_0414_),
    .B1(_0209_),
    .C1(_0418_),
    .D1(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__nor2_1 _1559_ (.A(\mem[0][31] ),
    .B(_0369_),
    .Y(_0423_));
 sky130_fd_sc_hd__nand2_1 _1560_ (.A(net69),
    .B(_0371_),
    .Y(_0424_));
 sky130_fd_sc_hd__o31ai_1 _1561_ (.A1(_0354_),
    .A2(_0422_),
    .A3(_0423_),
    .B1(_0424_),
    .Y(_0044_));
 sky130_fd_sc_hd__a21oi_1 _1562_ (.A1(\mem[3][3] ),
    .A2(_0657_),
    .B1(_0770_),
    .Y(_0425_));
 sky130_fd_sc_hd__a222oi_1 _1563_ (.A1(_0719_),
    .A2(\mem[7][3] ),
    .B1(\mem[4][3] ),
    .B2(_0759_),
    .C1(_0677_),
    .C2(\mem[6][3] ),
    .Y(_0426_));
 sky130_fd_sc_hd__a21oi_1 _1564_ (.A1(\mem[10][3] ),
    .A2(_0740_),
    .B1(_0203_),
    .Y(_0427_));
 sky130_fd_sc_hd__a222oi_1 _1565_ (.A1(\mem[14][3] ),
    .A2(_0666_),
    .B1(_0674_),
    .B2(\mem[13][3] ),
    .C1(\mem[12][3] ),
    .C2(_0162_),
    .Y(_0428_));
 sky130_fd_sc_hd__a22oi_1 _1566_ (.A1(_0425_),
    .A2(_0426_),
    .B1(_0427_),
    .B2(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__o21ai_0 _1567_ (.A1(_0425_),
    .A2(_0427_),
    .B1(_0207_),
    .Y(_0430_));
 sky130_fd_sc_hd__a32oi_1 _1568_ (.A1(_0742_),
    .A2(\mem[1][3] ),
    .A3(_0145_),
    .B1(_0166_),
    .B2(\mem[11][3] ),
    .Y(_0431_));
 sky130_fd_sc_hd__and3_1 _1569_ (.A(_0147_),
    .B(\mem[5][3] ),
    .C(_0717_),
    .X(_0432_));
 sky130_fd_sc_hd__a31oi_1 _1570_ (.A1(_0628_),
    .A2(\mem[2][3] ),
    .A3(_0168_),
    .B1(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__o22ai_2 _1571_ (.A1(_0655_),
    .A2(_0431_),
    .B1(_0433_),
    .B2(_0213_),
    .Y(_0434_));
 sky130_fd_sc_hd__a22oi_1 _1572_ (.A1(\mem[8][3] ),
    .A2(_0651_),
    .B1(_0215_),
    .B2(\mem[9][3] ),
    .Y(_0435_));
 sky130_fd_sc_hd__nand2_1 _1573_ (.A(\mem[15][3] ),
    .B(_0763_),
    .Y(_0436_));
 sky130_fd_sc_hd__o21ai_0 _1574_ (.A1(_0757_),
    .A2(_0435_),
    .B1(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__a2111oi_1 _1575_ (.A1(_0429_),
    .A2(_0430_),
    .B1(_0209_),
    .C1(_0434_),
    .D1(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__nor2_1 _1576_ (.A(\mem[0][3] ),
    .B(_0369_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand2_1 _1577_ (.A(net70),
    .B(_0371_),
    .Y(_0440_));
 sky130_fd_sc_hd__o31ai_1 _1578_ (.A1(_0354_),
    .A2(_0438_),
    .A3(_0439_),
    .B1(_0440_),
    .Y(_0045_));
 sky130_fd_sc_hd__a32o_1 _1579_ (.A1(_0748_),
    .A2(\mem[6][4] ),
    .A3(_0706_),
    .B1(_0749_),
    .B2(\mem[15][4] ),
    .X(_0441_));
 sky130_fd_sc_hd__nand3_1 _1580_ (.A(_0811_),
    .B(\mem[8][4] ),
    .C(_0760_),
    .Y(_0442_));
 sky130_fd_sc_hd__nand3_1 _1581_ (.A(_0682_),
    .B(\mem[1][4] ),
    .C(_0814_),
    .Y(_0443_));
 sky130_fd_sc_hd__a21oi_1 _1582_ (.A1(_0442_),
    .A2(_0443_),
    .B1(_0816_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand3_1 _1583_ (.A(_0649_),
    .B(\mem[13][4] ),
    .C(_0818_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand3_1 _1584_ (.A(_0820_),
    .B(\mem[10][4] ),
    .C(_0683_),
    .Y(_0446_));
 sky130_fd_sc_hd__and3_1 _1585_ (.A(_0648_),
    .B(\mem[4][4] ),
    .C(_0161_),
    .X(_0447_));
 sky130_fd_sc_hd__a211oi_1 _1586_ (.A1(\mem[3][4] ),
    .A2(_0658_),
    .B1(_0447_),
    .C1(_0825_),
    .Y(_0448_));
 sky130_fd_sc_hd__a31oi_1 _1587_ (.A1(_0688_),
    .A2(_0445_),
    .A3(_0446_),
    .B1(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__a22oi_2 _1588_ (.A1(\mem[7][4] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][4] ),
    .Y(_0450_));
 sky130_fd_sc_hd__and3_1 _1589_ (.A(_0644_),
    .B(_0822_),
    .C(\mem[14][4] ),
    .X(_0451_));
 sky130_fd_sc_hd__nor3b_1 _1590_ (.A(_0659_),
    .B(_0654_),
    .C_N(\mem[2][4] ),
    .Y(_0452_));
 sky130_fd_sc_hd__o21ai_0 _1591_ (.A1(_0451_),
    .A2(_0452_),
    .B1(_0678_),
    .Y(_0453_));
 sky130_fd_sc_hd__a22oi_1 _1592_ (.A1(_0636_),
    .A2(_0640_),
    .B1(_0694_),
    .B2(\mem[5][4] ),
    .Y(_0454_));
 sky130_fd_sc_hd__and3_1 _1593_ (.A(_0752_),
    .B(\mem[12][4] ),
    .C(_0823_),
    .X(_0455_));
 sky130_fd_sc_hd__and3b_1 _1594_ (.A_N(_0833_),
    .B(\mem[9][4] ),
    .C(_0813_),
    .X(_0456_));
 sky130_fd_sc_hd__o21ai_0 _1595_ (.A1(_0455_),
    .A2(_0456_),
    .B1(_0660_),
    .Y(_0457_));
 sky130_fd_sc_hd__o2111ai_2 _1596_ (.A1(_0829_),
    .A2(_0450_),
    .B1(_0453_),
    .C1(_0454_),
    .D1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__a2111oi_2 _1597_ (.A1(_0673_),
    .A2(_0441_),
    .B1(_0444_),
    .C1(_0449_),
    .D1(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor2_1 _1598_ (.A(\mem[0][4] ),
    .B(_0369_),
    .Y(_0460_));
 sky130_fd_sc_hd__nand2_1 _1599_ (.A(net71),
    .B(_0371_),
    .Y(_0461_));
 sky130_fd_sc_hd__o31ai_1 _1600_ (.A1(_0354_),
    .A2(_0459_),
    .A3(_0460_),
    .B1(_0461_),
    .Y(_0046_));
 sky130_fd_sc_hd__a21oi_1 _1601_ (.A1(\mem[3][5] ),
    .A2(_0657_),
    .B1(_0770_),
    .Y(_0462_));
 sky130_fd_sc_hd__a222oi_1 _1602_ (.A1(_0719_),
    .A2(\mem[7][5] ),
    .B1(\mem[4][5] ),
    .B2(_0759_),
    .C1(_0677_),
    .C2(\mem[6][5] ),
    .Y(_0463_));
 sky130_fd_sc_hd__a21oi_1 _1603_ (.A1(\mem[10][5] ),
    .A2(_0740_),
    .B1(_0203_),
    .Y(_0464_));
 sky130_fd_sc_hd__a222oi_1 _1604_ (.A1(\mem[14][5] ),
    .A2(_0666_),
    .B1(_0674_),
    .B2(\mem[13][5] ),
    .C1(\mem[12][5] ),
    .C2(_0162_),
    .Y(_0465_));
 sky130_fd_sc_hd__a22oi_1 _1605_ (.A1(_0462_),
    .A2(_0463_),
    .B1(_0464_),
    .B2(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__o21ai_0 _1606_ (.A1(_0462_),
    .A2(_0464_),
    .B1(_0207_),
    .Y(_0467_));
 sky130_fd_sc_hd__a32oi_1 _1607_ (.A1(_0742_),
    .A2(\mem[1][5] ),
    .A3(_0145_),
    .B1(_0166_),
    .B2(\mem[11][5] ),
    .Y(_0468_));
 sky130_fd_sc_hd__and3_1 _1608_ (.A(_0147_),
    .B(\mem[5][5] ),
    .C(_0717_),
    .X(_0469_));
 sky130_fd_sc_hd__a31oi_1 _1609_ (.A1(_0628_),
    .A2(\mem[2][5] ),
    .A3(_0168_),
    .B1(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__o22ai_1 _1610_ (.A1(_0655_),
    .A2(_0468_),
    .B1(_0470_),
    .B2(_0213_),
    .Y(_0471_));
 sky130_fd_sc_hd__a22oi_1 _1611_ (.A1(\mem[8][5] ),
    .A2(_0651_),
    .B1(_0215_),
    .B2(\mem[9][5] ),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _1612_ (.A(\mem[15][5] ),
    .B(_0763_),
    .Y(_0473_));
 sky130_fd_sc_hd__o21ai_0 _1613_ (.A1(_0757_),
    .A2(_0472_),
    .B1(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__a2111oi_0 _1614_ (.A1(_0466_),
    .A2(_0467_),
    .B1(_0209_),
    .C1(_0471_),
    .D1(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__nor2_1 _1615_ (.A(\mem[0][5] ),
    .B(_0369_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_1 _1616_ (.A(net72),
    .B(_0371_),
    .Y(_0477_));
 sky130_fd_sc_hd__o31ai_1 _1617_ (.A1(_0354_),
    .A2(_0475_),
    .A3(_0476_),
    .B1(_0477_),
    .Y(_0047_));
 sky130_fd_sc_hd__a32o_1 _1618_ (.A1(_0748_),
    .A2(\mem[6][6] ),
    .A3(_0706_),
    .B1(_0749_),
    .B2(\mem[15][6] ),
    .X(_0478_));
 sky130_fd_sc_hd__nand3_1 _1619_ (.A(_0825_),
    .B(\mem[8][6] ),
    .C(_0760_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand3_1 _1620_ (.A(_0682_),
    .B(\mem[1][6] ),
    .C(_0814_),
    .Y(_0480_));
 sky130_fd_sc_hd__a21oi_1 _1621_ (.A1(_0479_),
    .A2(_0480_),
    .B1(_0816_),
    .Y(_0481_));
 sky130_fd_sc_hd__nand3_1 _1622_ (.A(_0649_),
    .B(\mem[13][6] ),
    .C(_0818_),
    .Y(_0482_));
 sky130_fd_sc_hd__nand3_1 _1623_ (.A(_0820_),
    .B(\mem[10][6] ),
    .C(_0683_),
    .Y(_0483_));
 sky130_fd_sc_hd__and3_1 _1624_ (.A(_0648_),
    .B(\mem[4][6] ),
    .C(_0161_),
    .X(_0484_));
 sky130_fd_sc_hd__a211oi_1 _1625_ (.A1(\mem[3][6] ),
    .A2(_0733_),
    .B1(_0484_),
    .C1(_0663_),
    .Y(_0485_));
 sky130_fd_sc_hd__a31oi_1 _1626_ (.A1(_0688_),
    .A2(_0482_),
    .A3(_0483_),
    .B1(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__a22oi_4 _1627_ (.A1(\mem[7][6] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][6] ),
    .Y(_0487_));
 sky130_fd_sc_hd__and3_1 _1628_ (.A(_0644_),
    .B(_0822_),
    .C(\mem[14][6] ),
    .X(_0488_));
 sky130_fd_sc_hd__nor3b_1 _1629_ (.A(_0659_),
    .B(_0654_),
    .C_N(\mem[2][6] ),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_1 _1630_ (.A1(_0488_),
    .A2(_0489_),
    .B1(_0667_),
    .Y(_0490_));
 sky130_fd_sc_hd__a22oi_2 _1631_ (.A1(_0635_),
    .A2(_0639_),
    .B1(_0693_),
    .B2(\mem[5][6] ),
    .Y(_0491_));
 sky130_fd_sc_hd__and3_1 _1632_ (.A(_0752_),
    .B(\mem[12][6] ),
    .C(_0823_),
    .X(_0492_));
 sky130_fd_sc_hd__and3b_1 _1633_ (.A_N(_0833_),
    .B(\mem[9][6] ),
    .C(_0813_),
    .X(_0493_));
 sky130_fd_sc_hd__o21ai_1 _1634_ (.A1(_0492_),
    .A2(_0493_),
    .B1(_0660_),
    .Y(_0494_));
 sky130_fd_sc_hd__o2111ai_4 _1635_ (.A1(_0829_),
    .A2(_0487_),
    .B1(_0490_),
    .C1(_0491_),
    .D1(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__a2111oi_2 _1636_ (.A1(_0673_),
    .A2(_0478_),
    .B1(_0481_),
    .C1(_0486_),
    .D1(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__nor2_1 _1637_ (.A(\mem[0][6] ),
    .B(_0369_),
    .Y(_0497_));
 sky130_fd_sc_hd__nand2_1 _1638_ (.A(net73),
    .B(_0371_),
    .Y(_0498_));
 sky130_fd_sc_hd__o31ai_1 _1639_ (.A1(_0354_),
    .A2(_0496_),
    .A3(_0497_),
    .B1(_0498_),
    .Y(_0048_));
 sky130_fd_sc_hd__a21oi_1 _1640_ (.A1(\mem[3][7] ),
    .A2(_0657_),
    .B1(_0770_),
    .Y(_0499_));
 sky130_fd_sc_hd__a222oi_1 _1641_ (.A1(_0719_),
    .A2(\mem[7][7] ),
    .B1(\mem[4][7] ),
    .B2(_0759_),
    .C1(_0677_),
    .C2(\mem[6][7] ),
    .Y(_0500_));
 sky130_fd_sc_hd__a21oi_1 _1642_ (.A1(\mem[10][7] ),
    .A2(_0740_),
    .B1(_0203_),
    .Y(_0501_));
 sky130_fd_sc_hd__a222oi_1 _1643_ (.A1(\mem[14][7] ),
    .A2(_0666_),
    .B1(_0674_),
    .B2(\mem[13][7] ),
    .C1(\mem[12][7] ),
    .C2(_0162_),
    .Y(_0502_));
 sky130_fd_sc_hd__a22oi_1 _1644_ (.A1(_0499_),
    .A2(_0500_),
    .B1(_0501_),
    .B2(_0502_),
    .Y(_0503_));
 sky130_fd_sc_hd__o21ai_0 _1645_ (.A1(_0499_),
    .A2(_0501_),
    .B1(_0207_),
    .Y(_0504_));
 sky130_fd_sc_hd__a32oi_1 _1646_ (.A1(_0742_),
    .A2(\mem[1][7] ),
    .A3(_0710_),
    .B1(_0166_),
    .B2(\mem[11][7] ),
    .Y(_0505_));
 sky130_fd_sc_hd__and3_1 _1647_ (.A(_0712_),
    .B(\mem[5][7] ),
    .C(_0717_),
    .X(_0506_));
 sky130_fd_sc_hd__a31oi_1 _1648_ (.A1(_0628_),
    .A2(\mem[2][7] ),
    .A3(_0168_),
    .B1(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__o22ai_1 _1649_ (.A1(_0655_),
    .A2(_0505_),
    .B1(_0507_),
    .B2(_0213_),
    .Y(_0508_));
 sky130_fd_sc_hd__a22oi_1 _1650_ (.A1(\mem[8][7] ),
    .A2(_0651_),
    .B1(_0215_),
    .B2(\mem[9][7] ),
    .Y(_0509_));
 sky130_fd_sc_hd__nand2_1 _1651_ (.A(\mem[15][7] ),
    .B(_0763_),
    .Y(_0510_));
 sky130_fd_sc_hd__o21ai_0 _1652_ (.A1(_0757_),
    .A2(_0509_),
    .B1(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__a2111oi_1 _1653_ (.A1(_0503_),
    .A2(_0504_),
    .B1(_0209_),
    .C1(_0508_),
    .D1(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__nor2_1 _1654_ (.A(\mem[0][7] ),
    .B(_0369_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_1 _1655_ (.A(net74),
    .B(_0371_),
    .Y(_0514_));
 sky130_fd_sc_hd__o31ai_1 _1656_ (.A1(_0354_),
    .A2(_0512_),
    .A3(_0513_),
    .B1(_0514_),
    .Y(_0049_));
 sky130_fd_sc_hd__a32o_1 _1657_ (.A1(_0748_),
    .A2(\mem[6][8] ),
    .A3(_0706_),
    .B1(_0749_),
    .B2(\mem[15][8] ),
    .X(_0515_));
 sky130_fd_sc_hd__nand3_1 _1658_ (.A(_0825_),
    .B(\mem[8][8] ),
    .C(_0760_),
    .Y(_0516_));
 sky130_fd_sc_hd__nand3_1 _1659_ (.A(_0682_),
    .B(\mem[1][8] ),
    .C(_0814_),
    .Y(_0517_));
 sky130_fd_sc_hd__a21oi_1 _1660_ (.A1(_0516_),
    .A2(_0517_),
    .B1(_0816_),
    .Y(_0518_));
 sky130_fd_sc_hd__nand3_1 _1661_ (.A(_0649_),
    .B(\mem[13][8] ),
    .C(_0818_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand3_1 _1662_ (.A(_0820_),
    .B(\mem[10][8] ),
    .C(_0683_),
    .Y(_0520_));
 sky130_fd_sc_hd__and3_1 _1663_ (.A(_0648_),
    .B(\mem[4][8] ),
    .C(_0161_),
    .X(_0521_));
 sky130_fd_sc_hd__a211oi_1 _1664_ (.A1(\mem[3][8] ),
    .A2(_0733_),
    .B1(_0521_),
    .C1(_0663_),
    .Y(_0522_));
 sky130_fd_sc_hd__a31oi_1 _1665_ (.A1(_0645_),
    .A2(_0519_),
    .A3(_0520_),
    .B1(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__a22oi_2 _1666_ (.A1(\mem[7][8] ),
    .A2(_0830_),
    .B1(_0831_),
    .B2(\mem[11][8] ),
    .Y(_0524_));
 sky130_fd_sc_hd__and3_1 _1667_ (.A(_0644_),
    .B(_0822_),
    .C(\mem[14][8] ),
    .X(_0525_));
 sky130_fd_sc_hd__nor3b_1 _1668_ (.A(_0659_),
    .B(_0703_),
    .C_N(\mem[2][8] ),
    .Y(_0526_));
 sky130_fd_sc_hd__o21ai_1 _1669_ (.A1(_0525_),
    .A2(_0526_),
    .B1(_0667_),
    .Y(_0527_));
 sky130_fd_sc_hd__a22oi_2 _1670_ (.A1(_0635_),
    .A2(_0639_),
    .B1(_0693_),
    .B2(\mem[5][8] ),
    .Y(_0528_));
 sky130_fd_sc_hd__and3_1 _1671_ (.A(_0752_),
    .B(\mem[12][8] ),
    .C(_0823_),
    .X(_0529_));
 sky130_fd_sc_hd__and3b_1 _1672_ (.A_N(_0833_),
    .B(\mem[9][8] ),
    .C(_0813_),
    .X(_0530_));
 sky130_fd_sc_hd__o21ai_1 _1673_ (.A1(_0529_),
    .A2(_0530_),
    .B1(_0660_),
    .Y(_0531_));
 sky130_fd_sc_hd__o2111ai_4 _1674_ (.A1(_0828_),
    .A2(_0524_),
    .B1(_0527_),
    .C1(_0528_),
    .D1(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__a2111oi_0 _1675_ (.A1(_0673_),
    .A2(_0515_),
    .B1(_0518_),
    .C1(_0523_),
    .D1(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__nor2_1 _1676_ (.A(\mem[0][8] ),
    .B(_0369_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _1677_ (.A(net75),
    .B(_0371_),
    .Y(_0535_));
 sky130_fd_sc_hd__o31ai_1 _1678_ (.A1(_0354_),
    .A2(_0533_),
    .A3(_0534_),
    .B1(_0535_),
    .Y(_0050_));
 sky130_fd_sc_hd__a21oi_1 _1679_ (.A1(\mem[3][9] ),
    .A2(_0657_),
    .B1(_0770_),
    .Y(_0536_));
 sky130_fd_sc_hd__a222oi_1 _1680_ (.A1(_0719_),
    .A2(\mem[7][9] ),
    .B1(\mem[4][9] ),
    .B2(_0759_),
    .C1(_0677_),
    .C2(\mem[6][9] ),
    .Y(_0537_));
 sky130_fd_sc_hd__a21oi_1 _1681_ (.A1(\mem[10][9] ),
    .A2(_0740_),
    .B1(_0203_),
    .Y(_0538_));
 sky130_fd_sc_hd__a222oi_1 _1682_ (.A1(\mem[14][9] ),
    .A2(_0666_),
    .B1(_0674_),
    .B2(\mem[13][9] ),
    .C1(\mem[12][9] ),
    .C2(_0709_),
    .Y(_0539_));
 sky130_fd_sc_hd__a22oi_1 _1683_ (.A1(_0536_),
    .A2(_0537_),
    .B1(_0538_),
    .B2(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__o21ai_0 _1684_ (.A1(_0536_),
    .A2(_0538_),
    .B1(_0207_),
    .Y(_0541_));
 sky130_fd_sc_hd__a32oi_1 _1685_ (.A1(_0742_),
    .A2(\mem[1][9] ),
    .A3(_0710_),
    .B1(_0685_),
    .B2(\mem[11][9] ),
    .Y(_0542_));
 sky130_fd_sc_hd__and3_1 _1686_ (.A(_0712_),
    .B(\mem[5][9] ),
    .C(_0717_),
    .X(_0543_));
 sky130_fd_sc_hd__a31oi_1 _1687_ (.A1(_0628_),
    .A2(\mem[2][9] ),
    .A3(_0647_),
    .B1(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__o22ai_2 _1688_ (.A1(_0655_),
    .A2(_0542_),
    .B1(_0544_),
    .B2(_0213_),
    .Y(_0545_));
 sky130_fd_sc_hd__a22oi_1 _1689_ (.A1(\mem[8][9] ),
    .A2(_0651_),
    .B1(_0215_),
    .B2(\mem[9][9] ),
    .Y(_0546_));
 sky130_fd_sc_hd__nand2_1 _1690_ (.A(\mem[15][9] ),
    .B(_0763_),
    .Y(_0547_));
 sky130_fd_sc_hd__o21ai_1 _1691_ (.A1(_0757_),
    .A2(_0546_),
    .B1(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__a2111oi_2 _1692_ (.A1(_0540_),
    .A2(_0541_),
    .B1(_0209_),
    .C1(_0545_),
    .D1(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__nor2_1 _1693_ (.A(\mem[0][9] ),
    .B(_0641_),
    .Y(_0550_));
 sky130_fd_sc_hd__buf_6 _1694_ (.A(_0633_),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _1695_ (.A(net76),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__o31ai_1 _1696_ (.A1(_0633_),
    .A2(_0549_),
    .A3(_0550_),
    .B1(_0552_),
    .Y(_0051_));
 sky130_fd_sc_hd__xnor2_1 _1697_ (.A(\rd_ptr_bin[0] ),
    .B(_0551_),
    .Y(_0052_));
 sky130_fd_sc_hd__mux2_1 _1698_ (.A0(_0019_),
    .A1(\rd_ptr_bin[1] ),
    .S(_0633_),
    .X(_0053_));
 sky130_fd_sc_hd__nor2_1 _1699_ (.A(_0829_),
    .B(_0633_),
    .Y(_0553_));
 sky130_fd_sc_hd__xnor2_1 _1700_ (.A(_0867_),
    .B(_0553_),
    .Y(_0054_));
 sky130_fd_sc_hd__nand3_1 _1701_ (.A(_0649_),
    .B(\rd_ptr_bin[0] ),
    .C(\rd_ptr_bin[1] ),
    .Y(_0554_));
 sky130_fd_sc_hd__nor2_1 _1702_ (.A(_0633_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__xnor2_1 _1703_ (.A(_0863_),
    .B(_0555_),
    .Y(_0055_));
 sky130_fd_sc_hd__xor2_1 _1704_ (.A(\rd_ptr_bin[0] ),
    .B(_0019_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_1 _1705_ (.A(\rd_ptr_gray[0] ),
    .B(_0551_),
    .Y(_0557_));
 sky130_fd_sc_hd__o21ai_0 _1706_ (.A1(_0551_),
    .A2(_0556_),
    .B1(_0557_),
    .Y(_0056_));
 sky130_fd_sc_hd__xor2_2 _1707_ (.A(_0783_),
    .B(_0698_),
    .X(_0558_));
 sky130_fd_sc_hd__xnor2_1 _1708_ (.A(_0019_),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _1709_ (.A(\rd_ptr_gray[1] ),
    .B(_0551_),
    .Y(_0560_));
 sky130_fd_sc_hd__o21ai_0 _1710_ (.A1(_0551_),
    .A2(_0559_),
    .B1(_0560_),
    .Y(_0057_));
 sky130_fd_sc_hd__xnor2_1 _1711_ (.A(_0863_),
    .B(_0554_),
    .Y(_0561_));
 sky130_fd_sc_hd__xor2_1 _1712_ (.A(_0558_),
    .B(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__nand2_1 _1713_ (.A(\rd_ptr_gray[2] ),
    .B(_0551_),
    .Y(_0563_));
 sky130_fd_sc_hd__o21ai_0 _1714_ (.A1(_0551_),
    .A2(_0562_),
    .B1(_0563_),
    .Y(_0058_));
 sky130_fd_sc_hd__xnor2_1 _1715_ (.A(\rd_ptr_bin[4] ),
    .B(_0764_),
    .Y(_0564_));
 sky130_fd_sc_hd__xnor2_1 _1716_ (.A(_0561_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__nand2_1 _1717_ (.A(\rd_ptr_gray[3] ),
    .B(_0551_),
    .Y(_0566_));
 sky130_fd_sc_hd__o21ai_0 _1718_ (.A1(_0551_),
    .A2(_0565_),
    .B1(_0566_),
    .Y(_0059_));
 sky130_fd_sc_hd__nand3_1 _1719_ (.A(net2),
    .B(_0625_),
    .C(_0764_),
    .Y(_0567_));
 sky130_fd_sc_hd__xnor2_1 _1720_ (.A(\rd_ptr_bin[4] ),
    .B(_0567_),
    .Y(_0060_));
 sky130_fd_sc_hd__xnor2_1 _1721_ (.A(_0631_),
    .B(_0605_),
    .Y(_0061_));
 sky130_fd_sc_hd__nand2_1 _1722_ (.A(_0017_),
    .B(_0595_),
    .Y(_0568_));
 sky130_fd_sc_hd__o21ai_0 _1723_ (.A1(_0841_),
    .A2(_0595_),
    .B1(_0568_),
    .Y(_0062_));
 sky130_fd_sc_hd__nand2_1 _1724_ (.A(_0608_),
    .B(_0595_),
    .Y(_0569_));
 sky130_fd_sc_hd__xnor2_1 _1725_ (.A(_0592_),
    .B(_0569_),
    .Y(_0063_));
 sky130_fd_sc_hd__nand4_1 _1726_ (.A(_0592_),
    .B(_0631_),
    .C(\wr_ptr_bin[1] ),
    .D(_0595_),
    .Y(_0570_));
 sky130_fd_sc_hd__xnor2_1 _1727_ (.A(_0593_),
    .B(_0570_),
    .Y(_0064_));
 sky130_fd_sc_hd__xor2_1 _1728_ (.A(_0631_),
    .B(_0017_),
    .X(_0571_));
 sky130_fd_sc_hd__nand2_1 _1729_ (.A(\wr_ptr_gray[0] ),
    .B(_0605_),
    .Y(_0572_));
 sky130_fd_sc_hd__o21ai_0 _1730_ (.A1(_0605_),
    .A2(_0571_),
    .B1(_0572_),
    .Y(_0065_));
 sky130_fd_sc_hd__xor2_1 _1731_ (.A(_0608_),
    .B(_0017_),
    .X(_0573_));
 sky130_fd_sc_hd__xnor2_1 _1732_ (.A(_0592_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand2_1 _1733_ (.A(\wr_ptr_gray[1] ),
    .B(_0605_),
    .Y(_0575_));
 sky130_fd_sc_hd__o21ai_0 _1734_ (.A1(_0605_),
    .A2(_0574_),
    .B1(_0575_),
    .Y(_0066_));
 sky130_fd_sc_hd__xnor2_1 _1735_ (.A(_0593_),
    .B(_0608_),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_1 _1736_ (.A(_0631_),
    .B(\wr_ptr_bin[1] ),
    .Y(_0577_));
 sky130_fd_sc_hd__nand2_1 _1737_ (.A(_0592_),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__xnor2_1 _1738_ (.A(_0576_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2_1 _1739_ (.A(\wr_ptr_gray[2] ),
    .B(_0605_),
    .Y(_0580_));
 sky130_fd_sc_hd__o21ai_0 _1740_ (.A1(_0605_),
    .A2(_0579_),
    .B1(_0580_),
    .Y(_0067_));
 sky130_fd_sc_hd__nand2_1 _1741_ (.A(\wr_ptr_bin[2] ),
    .B(_0608_),
    .Y(_0581_));
 sky130_fd_sc_hd__a21boi_0 _1742_ (.A1(_0593_),
    .A2(_0581_),
    .B1_N(_0577_),
    .Y(_0582_));
 sky130_fd_sc_hd__nand4_1 _1743_ (.A(\wr_ptr_bin[2] ),
    .B(_0593_),
    .C(_0631_),
    .D(\wr_ptr_bin[1] ),
    .Y(_0583_));
 sky130_fd_sc_hd__o22ai_1 _1744_ (.A1(_0592_),
    .A2(_0593_),
    .B1(_0608_),
    .B2(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__nor2_1 _1745_ (.A(_0582_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__xnor2_1 _1746_ (.A(\wr_ptr_bin[4] ),
    .B(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_1 _1747_ (.A(\wr_ptr_gray[3] ),
    .B(_0605_),
    .Y(_0587_));
 sky130_fd_sc_hd__o21ai_0 _1748_ (.A1(_0605_),
    .A2(_0586_),
    .B1(_0587_),
    .Y(_0068_));
 sky130_fd_sc_hd__nand4_1 _1749_ (.A(_0592_),
    .B(_0593_),
    .C(_0608_),
    .D(_0595_),
    .Y(_0588_));
 sky130_fd_sc_hd__xnor2_1 _1750_ (.A(\wr_ptr_bin[4] ),
    .B(_0588_),
    .Y(_0069_));
 sky130_fd_sc_hd__a21oi_1 _1751_ (.A1(net40),
    .A2(net41),
    .B1(net42),
    .Y(_0589_));
 sky130_fd_sc_hd__nor4b_1 _1752_ (.A(net43),
    .B(net44),
    .C(net77),
    .D_N(_0589_),
    .Y(net39));
 sky130_fd_sc_hd__inv_1 _1753_ (.A(_0845_),
    .Y(net80));
 sky130_fd_sc_hd__xnor2_1 _1754_ (.A(_0844_),
    .B(_0855_),
    .Y(net81));
 sky130_fd_sc_hd__a31o_1 _1755_ (.A1(net80),
    .A2(net82),
    .A3(net81),
    .B1(net83),
    .X(net78));
 sky130_fd_sc_hd__fa_1 _1756_ (.A(_0841_),
    .B(_0842_),
    .CIN(_0843_),
    .COUT(_0844_),
    .SUM(_0845_));
 sky130_fd_sc_hd__fa_1 _1757_ (.A(\rd_ptr_bin[1] ),
    .B(_0847_),
    .CIN(_0848_),
    .COUT(_0849_),
    .SUM(_0850_));
 sky130_fd_sc_hd__ha_1 _1758_ (.A(\wr_ptr_bin[1] ),
    .B(_0846_),
    .COUT(_0851_),
    .SUM(_0852_));
 sky130_fd_sc_hd__ha_1 _1759_ (.A(\wr_ptr_bin[2] ),
    .B(_0853_),
    .COUT(_0854_),
    .SUM(_0855_));
 sky130_fd_sc_hd__ha_1 _1760_ (.A(\wr_ptr_bin[3] ),
    .B(_0856_),
    .COUT(_0857_),
    .SUM(_0858_));
 sky130_fd_sc_hd__ha_1 _1761_ (.A(_0859_),
    .B(_0860_),
    .COUT(_0861_),
    .SUM(_0862_));
 sky130_fd_sc_hd__ha_1 _1762_ (.A(_0863_),
    .B(_0864_),
    .COUT(_0865_),
    .SUM(_0866_));
 sky130_fd_sc_hd__ha_1 _1763_ (.A(_0867_),
    .B(_0868_),
    .COUT(_0869_),
    .SUM(_0870_));
 sky130_fd_sc_hd__ha_1 _1764_ (.A(_0016_),
    .B(_0841_),
    .COUT(_0871_),
    .SUM(_0017_));
 sky130_fd_sc_hd__ha_1 _1765_ (.A(_0016_),
    .B(\wr_ptr_bin[1] ),
    .COUT(_0872_),
    .SUM(_0873_));
 sky130_fd_sc_hd__ha_1 _1766_ (.A(\wr_ptr_bin[0] ),
    .B(_0841_),
    .COUT(_0874_),
    .SUM(_0875_));
 sky130_fd_sc_hd__ha_1 _1767_ (.A(\wr_ptr_bin[0] ),
    .B(\wr_ptr_bin[1] ),
    .COUT(_0876_),
    .SUM(_0877_));
 sky130_fd_sc_hd__ha_1 _1768_ (.A(_0018_),
    .B(_0859_),
    .COUT(_0878_),
    .SUM(_0019_));
 sky130_fd_sc_hd__ha_2 _1769_ (.A(_0018_),
    .B(\rd_ptr_bin[1] ),
    .COUT(_0879_),
    .SUM(_0880_));
 sky130_fd_sc_hd__ha_1 _1770_ (.A(\rd_ptr_bin[0] ),
    .B(_0859_),
    .COUT(_0881_),
    .SUM(_0882_));
 sky130_fd_sc_hd__ha_1 _1771_ (.A(\rd_ptr_bin[0] ),
    .B(\rd_ptr_bin[1] ),
    .COUT(_0883_),
    .SUM(_0884_));
 sky130_fd_sc_hd__ha_1 _1772_ (.A(\rd_ptr_bin[0] ),
    .B(_0885_),
    .COUT(_0847_),
    .SUM(_0886_));
 sky130_fd_sc_hd__ha_1 _1773_ (.A(_0016_),
    .B(_0887_),
    .COUT(_0842_),
    .SUM(_0888_));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net5),
    .DE(_0015_),
    .Q(\mem[0][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][10]$_DFFE_PP_  (.D(net6),
    .DE(_0015_),
    .Q(\mem[0][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][11]$_DFFE_PP_  (.D(net7),
    .DE(_0015_),
    .Q(\mem[0][11] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][12]$_DFFE_PP_  (.D(net8),
    .DE(_0015_),
    .Q(\mem[0][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][13]$_DFFE_PP_  (.D(net9),
    .DE(_0015_),
    .Q(\mem[0][13] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][14]$_DFFE_PP_  (.D(net10),
    .DE(_0015_),
    .Q(\mem[0][14] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][15]$_DFFE_PP_  (.D(net11),
    .DE(_0015_),
    .Q(\mem[0][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][16]$_DFFE_PP_  (.D(net12),
    .DE(_0015_),
    .Q(\mem[0][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][17]$_DFFE_PP_  (.D(net13),
    .DE(_0015_),
    .Q(\mem[0][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][18]$_DFFE_PP_  (.D(net14),
    .DE(_0015_),
    .Q(\mem[0][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][19]$_DFFE_PP_  (.D(net15),
    .DE(_0015_),
    .Q(\mem[0][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net16),
    .DE(_0015_),
    .Q(\mem[0][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][20]$_DFFE_PP_  (.D(net17),
    .DE(_0015_),
    .Q(\mem[0][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][21]$_DFFE_PP_  (.D(net18),
    .DE(_0015_),
    .Q(\mem[0][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][22]$_DFFE_PP_  (.D(net19),
    .DE(_0015_),
    .Q(\mem[0][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][23]$_DFFE_PP_  (.D(net20),
    .DE(_0015_),
    .Q(\mem[0][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][24]$_DFFE_PP_  (.D(net21),
    .DE(_0015_),
    .Q(\mem[0][24] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][25]$_DFFE_PP_  (.D(net22),
    .DE(_0015_),
    .Q(\mem[0][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][26]$_DFFE_PP_  (.D(net23),
    .DE(_0015_),
    .Q(\mem[0][26] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][27]$_DFFE_PP_  (.D(net24),
    .DE(_0015_),
    .Q(\mem[0][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][28]$_DFFE_PP_  (.D(net25),
    .DE(_0015_),
    .Q(\mem[0][28] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][29]$_DFFE_PP_  (.D(net26),
    .DE(_0015_),
    .Q(\mem[0][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net27),
    .DE(_0015_),
    .Q(\mem[0][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][30]$_DFFE_PP_  (.D(net28),
    .DE(_0015_),
    .Q(\mem[0][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][31]$_DFFE_PP_  (.D(net29),
    .DE(_0015_),
    .Q(\mem[0][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net30),
    .DE(_0015_),
    .Q(\mem[0][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net31),
    .DE(_0015_),
    .Q(\mem[0][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net32),
    .DE(_0015_),
    .Q(\mem[0][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net33),
    .DE(_0015_),
    .Q(\mem[0][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net34),
    .DE(_0015_),
    .Q(\mem[0][7] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][8]$_DFFE_PP_  (.D(net35),
    .DE(_0015_),
    .Q(\mem[0][8] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][9]$_DFFE_PP_  (.D(net36),
    .DE(_0015_),
    .Q(\mem[0][9] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net5),
    .DE(_0005_),
    .Q(\mem[10][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][10]$_DFFE_PP_  (.D(net6),
    .DE(_0005_),
    .Q(\mem[10][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][11]$_DFFE_PP_  (.D(net7),
    .DE(_0005_),
    .Q(\mem[10][11] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][12]$_DFFE_PP_  (.D(net8),
    .DE(_0005_),
    .Q(\mem[10][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][13]$_DFFE_PP_  (.D(net9),
    .DE(_0005_),
    .Q(\mem[10][13] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][14]$_DFFE_PP_  (.D(net10),
    .DE(_0005_),
    .Q(\mem[10][14] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][15]$_DFFE_PP_  (.D(net11),
    .DE(_0005_),
    .Q(\mem[10][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][16]$_DFFE_PP_  (.D(net12),
    .DE(_0005_),
    .Q(\mem[10][16] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][17]$_DFFE_PP_  (.D(net13),
    .DE(_0005_),
    .Q(\mem[10][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][18]$_DFFE_PP_  (.D(net14),
    .DE(_0005_),
    .Q(\mem[10][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][19]$_DFFE_PP_  (.D(net15),
    .DE(_0005_),
    .Q(\mem[10][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net16),
    .DE(_0005_),
    .Q(\mem[10][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][20]$_DFFE_PP_  (.D(net17),
    .DE(_0005_),
    .Q(\mem[10][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][21]$_DFFE_PP_  (.D(net18),
    .DE(_0005_),
    .Q(\mem[10][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][22]$_DFFE_PP_  (.D(net19),
    .DE(_0005_),
    .Q(\mem[10][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][23]$_DFFE_PP_  (.D(net20),
    .DE(_0005_),
    .Q(\mem[10][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][24]$_DFFE_PP_  (.D(net21),
    .DE(_0005_),
    .Q(\mem[10][24] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][25]$_DFFE_PP_  (.D(net22),
    .DE(_0005_),
    .Q(\mem[10][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][26]$_DFFE_PP_  (.D(net23),
    .DE(_0005_),
    .Q(\mem[10][26] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][27]$_DFFE_PP_  (.D(net24),
    .DE(_0005_),
    .Q(\mem[10][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][28]$_DFFE_PP_  (.D(net25),
    .DE(_0005_),
    .Q(\mem[10][28] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][29]$_DFFE_PP_  (.D(net26),
    .DE(_0005_),
    .Q(\mem[10][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net27),
    .DE(_0005_),
    .Q(\mem[10][2] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][30]$_DFFE_PP_  (.D(net28),
    .DE(_0005_),
    .Q(\mem[10][30] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][31]$_DFFE_PP_  (.D(net29),
    .DE(_0005_),
    .Q(\mem[10][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net30),
    .DE(_0005_),
    .Q(\mem[10][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net31),
    .DE(_0005_),
    .Q(\mem[10][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net32),
    .DE(_0005_),
    .Q(\mem[10][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net33),
    .DE(_0005_),
    .Q(\mem[10][6] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net34),
    .DE(_0005_),
    .Q(\mem[10][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][8]$_DFFE_PP_  (.D(net35),
    .DE(_0005_),
    .Q(\mem[10][8] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][9]$_DFFE_PP_  (.D(net36),
    .DE(_0005_),
    .Q(\mem[10][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net5),
    .DE(_0004_),
    .Q(\mem[11][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][10]$_DFFE_PP_  (.D(net6),
    .DE(_0004_),
    .Q(\mem[11][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][11]$_DFFE_PP_  (.D(net7),
    .DE(_0004_),
    .Q(\mem[11][11] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][12]$_DFFE_PP_  (.D(net8),
    .DE(_0004_),
    .Q(\mem[11][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][13]$_DFFE_PP_  (.D(net9),
    .DE(_0004_),
    .Q(\mem[11][13] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][14]$_DFFE_PP_  (.D(net10),
    .DE(_0004_),
    .Q(\mem[11][14] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][15]$_DFFE_PP_  (.D(net11),
    .DE(_0004_),
    .Q(\mem[11][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][16]$_DFFE_PP_  (.D(net12),
    .DE(_0004_),
    .Q(\mem[11][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][17]$_DFFE_PP_  (.D(net13),
    .DE(_0004_),
    .Q(\mem[11][17] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][18]$_DFFE_PP_  (.D(net14),
    .DE(_0004_),
    .Q(\mem[11][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][19]$_DFFE_PP_  (.D(net15),
    .DE(_0004_),
    .Q(\mem[11][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net16),
    .DE(_0004_),
    .Q(\mem[11][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][20]$_DFFE_PP_  (.D(net17),
    .DE(_0004_),
    .Q(\mem[11][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][21]$_DFFE_PP_  (.D(net18),
    .DE(_0004_),
    .Q(\mem[11][21] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][22]$_DFFE_PP_  (.D(net19),
    .DE(_0004_),
    .Q(\mem[11][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][23]$_DFFE_PP_  (.D(net20),
    .DE(_0004_),
    .Q(\mem[11][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][24]$_DFFE_PP_  (.D(net21),
    .DE(_0004_),
    .Q(\mem[11][24] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][25]$_DFFE_PP_  (.D(net22),
    .DE(_0004_),
    .Q(\mem[11][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][26]$_DFFE_PP_  (.D(net23),
    .DE(_0004_),
    .Q(\mem[11][26] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][27]$_DFFE_PP_  (.D(net24),
    .DE(_0004_),
    .Q(\mem[11][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][28]$_DFFE_PP_  (.D(net25),
    .DE(_0004_),
    .Q(\mem[11][28] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][29]$_DFFE_PP_  (.D(net26),
    .DE(_0004_),
    .Q(\mem[11][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net27),
    .DE(_0004_),
    .Q(\mem[11][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][30]$_DFFE_PP_  (.D(net28),
    .DE(_0004_),
    .Q(\mem[11][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][31]$_DFFE_PP_  (.D(net29),
    .DE(_0004_),
    .Q(\mem[11][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net30),
    .DE(_0004_),
    .Q(\mem[11][3] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net31),
    .DE(_0004_),
    .Q(\mem[11][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net32),
    .DE(_0004_),
    .Q(\mem[11][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net33),
    .DE(_0004_),
    .Q(\mem[11][6] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net34),
    .DE(_0004_),
    .Q(\mem[11][7] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][8]$_DFFE_PP_  (.D(net35),
    .DE(_0004_),
    .Q(\mem[11][8] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][9]$_DFFE_PP_  (.D(net36),
    .DE(_0004_),
    .Q(\mem[11][9] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net5),
    .DE(_0003_),
    .Q(\mem[12][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][10]$_DFFE_PP_  (.D(net6),
    .DE(_0003_),
    .Q(\mem[12][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][11]$_DFFE_PP_  (.D(net7),
    .DE(_0003_),
    .Q(\mem[12][11] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][12]$_DFFE_PP_  (.D(net8),
    .DE(_0003_),
    .Q(\mem[12][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][13]$_DFFE_PP_  (.D(net9),
    .DE(_0003_),
    .Q(\mem[12][13] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][14]$_DFFE_PP_  (.D(net10),
    .DE(_0003_),
    .Q(\mem[12][14] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][15]$_DFFE_PP_  (.D(net11),
    .DE(_0003_),
    .Q(\mem[12][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][16]$_DFFE_PP_  (.D(net12),
    .DE(_0003_),
    .Q(\mem[12][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][17]$_DFFE_PP_  (.D(net13),
    .DE(_0003_),
    .Q(\mem[12][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][18]$_DFFE_PP_  (.D(net14),
    .DE(_0003_),
    .Q(\mem[12][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][19]$_DFFE_PP_  (.D(net15),
    .DE(_0003_),
    .Q(\mem[12][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net16),
    .DE(_0003_),
    .Q(\mem[12][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][20]$_DFFE_PP_  (.D(net17),
    .DE(_0003_),
    .Q(\mem[12][20] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][21]$_DFFE_PP_  (.D(net18),
    .DE(_0003_),
    .Q(\mem[12][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][22]$_DFFE_PP_  (.D(net19),
    .DE(_0003_),
    .Q(\mem[12][22] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][23]$_DFFE_PP_  (.D(net20),
    .DE(_0003_),
    .Q(\mem[12][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][24]$_DFFE_PP_  (.D(net21),
    .DE(_0003_),
    .Q(\mem[12][24] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][25]$_DFFE_PP_  (.D(net22),
    .DE(_0003_),
    .Q(\mem[12][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][26]$_DFFE_PP_  (.D(net23),
    .DE(_0003_),
    .Q(\mem[12][26] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][27]$_DFFE_PP_  (.D(net24),
    .DE(_0003_),
    .Q(\mem[12][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][28]$_DFFE_PP_  (.D(net25),
    .DE(_0003_),
    .Q(\mem[12][28] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][29]$_DFFE_PP_  (.D(net26),
    .DE(_0003_),
    .Q(\mem[12][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net27),
    .DE(_0003_),
    .Q(\mem[12][2] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][30]$_DFFE_PP_  (.D(net28),
    .DE(_0003_),
    .Q(\mem[12][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][31]$_DFFE_PP_  (.D(net29),
    .DE(_0003_),
    .Q(\mem[12][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net30),
    .DE(_0003_),
    .Q(\mem[12][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net31),
    .DE(_0003_),
    .Q(\mem[12][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net32),
    .DE(_0003_),
    .Q(\mem[12][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net33),
    .DE(_0003_),
    .Q(\mem[12][6] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net34),
    .DE(_0003_),
    .Q(\mem[12][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][8]$_DFFE_PP_  (.D(net35),
    .DE(_0003_),
    .Q(\mem[12][8] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][9]$_DFFE_PP_  (.D(net36),
    .DE(_0003_),
    .Q(\mem[12][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net5),
    .DE(_0002_),
    .Q(\mem[13][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][10]$_DFFE_PP_  (.D(net6),
    .DE(_0002_),
    .Q(\mem[13][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][11]$_DFFE_PP_  (.D(net7),
    .DE(_0002_),
    .Q(\mem[13][11] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][12]$_DFFE_PP_  (.D(net8),
    .DE(_0002_),
    .Q(\mem[13][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][13]$_DFFE_PP_  (.D(net9),
    .DE(_0002_),
    .Q(\mem[13][13] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][14]$_DFFE_PP_  (.D(net10),
    .DE(_0002_),
    .Q(\mem[13][14] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][15]$_DFFE_PP_  (.D(net11),
    .DE(_0002_),
    .Q(\mem[13][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][16]$_DFFE_PP_  (.D(net12),
    .DE(_0002_),
    .Q(\mem[13][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][17]$_DFFE_PP_  (.D(net13),
    .DE(_0002_),
    .Q(\mem[13][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][18]$_DFFE_PP_  (.D(net14),
    .DE(_0002_),
    .Q(\mem[13][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][19]$_DFFE_PP_  (.D(net15),
    .DE(_0002_),
    .Q(\mem[13][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net16),
    .DE(_0002_),
    .Q(\mem[13][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][20]$_DFFE_PP_  (.D(net17),
    .DE(_0002_),
    .Q(\mem[13][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][21]$_DFFE_PP_  (.D(net18),
    .DE(_0002_),
    .Q(\mem[13][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][22]$_DFFE_PP_  (.D(net19),
    .DE(_0002_),
    .Q(\mem[13][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][23]$_DFFE_PP_  (.D(net20),
    .DE(_0002_),
    .Q(\mem[13][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][24]$_DFFE_PP_  (.D(net21),
    .DE(_0002_),
    .Q(\mem[13][24] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][25]$_DFFE_PP_  (.D(net22),
    .DE(_0002_),
    .Q(\mem[13][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][26]$_DFFE_PP_  (.D(net23),
    .DE(_0002_),
    .Q(\mem[13][26] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][27]$_DFFE_PP_  (.D(net24),
    .DE(_0002_),
    .Q(\mem[13][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][28]$_DFFE_PP_  (.D(net25),
    .DE(_0002_),
    .Q(\mem[13][28] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][29]$_DFFE_PP_  (.D(net26),
    .DE(_0002_),
    .Q(\mem[13][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net27),
    .DE(_0002_),
    .Q(\mem[13][2] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][30]$_DFFE_PP_  (.D(net28),
    .DE(_0002_),
    .Q(\mem[13][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][31]$_DFFE_PP_  (.D(net29),
    .DE(_0002_),
    .Q(\mem[13][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net30),
    .DE(_0002_),
    .Q(\mem[13][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net31),
    .DE(_0002_),
    .Q(\mem[13][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net32),
    .DE(_0002_),
    .Q(\mem[13][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net33),
    .DE(_0002_),
    .Q(\mem[13][6] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net34),
    .DE(_0002_),
    .Q(\mem[13][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][8]$_DFFE_PP_  (.D(net35),
    .DE(_0002_),
    .Q(\mem[13][8] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][9]$_DFFE_PP_  (.D(net36),
    .DE(_0002_),
    .Q(\mem[13][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net5),
    .DE(_0001_),
    .Q(\mem[14][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][10]$_DFFE_PP_  (.D(net6),
    .DE(_0001_),
    .Q(\mem[14][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][11]$_DFFE_PP_  (.D(net7),
    .DE(_0001_),
    .Q(\mem[14][11] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][12]$_DFFE_PP_  (.D(net8),
    .DE(_0001_),
    .Q(\mem[14][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][13]$_DFFE_PP_  (.D(net9),
    .DE(_0001_),
    .Q(\mem[14][13] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][14]$_DFFE_PP_  (.D(net10),
    .DE(_0001_),
    .Q(\mem[14][14] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][15]$_DFFE_PP_  (.D(net11),
    .DE(_0001_),
    .Q(\mem[14][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][16]$_DFFE_PP_  (.D(net12),
    .DE(_0001_),
    .Q(\mem[14][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][17]$_DFFE_PP_  (.D(net13),
    .DE(_0001_),
    .Q(\mem[14][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][18]$_DFFE_PP_  (.D(net14),
    .DE(_0001_),
    .Q(\mem[14][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][19]$_DFFE_PP_  (.D(net15),
    .DE(_0001_),
    .Q(\mem[14][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net16),
    .DE(_0001_),
    .Q(\mem[14][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][20]$_DFFE_PP_  (.D(net17),
    .DE(_0001_),
    .Q(\mem[14][20] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][21]$_DFFE_PP_  (.D(net18),
    .DE(_0001_),
    .Q(\mem[14][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][22]$_DFFE_PP_  (.D(net19),
    .DE(_0001_),
    .Q(\mem[14][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][23]$_DFFE_PP_  (.D(net20),
    .DE(_0001_),
    .Q(\mem[14][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][24]$_DFFE_PP_  (.D(net21),
    .DE(_0001_),
    .Q(\mem[14][24] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][25]$_DFFE_PP_  (.D(net22),
    .DE(_0001_),
    .Q(\mem[14][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][26]$_DFFE_PP_  (.D(net23),
    .DE(_0001_),
    .Q(\mem[14][26] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][27]$_DFFE_PP_  (.D(net24),
    .DE(_0001_),
    .Q(\mem[14][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][28]$_DFFE_PP_  (.D(net25),
    .DE(_0001_),
    .Q(\mem[14][28] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][29]$_DFFE_PP_  (.D(net26),
    .DE(_0001_),
    .Q(\mem[14][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net27),
    .DE(_0001_),
    .Q(\mem[14][2] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][30]$_DFFE_PP_  (.D(net28),
    .DE(_0001_),
    .Q(\mem[14][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][31]$_DFFE_PP_  (.D(net29),
    .DE(_0001_),
    .Q(\mem[14][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net30),
    .DE(_0001_),
    .Q(\mem[14][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net31),
    .DE(_0001_),
    .Q(\mem[14][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net32),
    .DE(_0001_),
    .Q(\mem[14][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net33),
    .DE(_0001_),
    .Q(\mem[14][6] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net34),
    .DE(_0001_),
    .Q(\mem[14][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][8]$_DFFE_PP_  (.D(net35),
    .DE(_0001_),
    .Q(\mem[14][8] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][9]$_DFFE_PP_  (.D(net36),
    .DE(_0001_),
    .Q(\mem[14][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net5),
    .DE(_0000_),
    .Q(\mem[15][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][10]$_DFFE_PP_  (.D(net6),
    .DE(_0000_),
    .Q(\mem[15][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][11]$_DFFE_PP_  (.D(net7),
    .DE(_0000_),
    .Q(\mem[15][11] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][12]$_DFFE_PP_  (.D(net8),
    .DE(_0000_),
    .Q(\mem[15][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][13]$_DFFE_PP_  (.D(net9),
    .DE(_0000_),
    .Q(\mem[15][13] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][14]$_DFFE_PP_  (.D(net10),
    .DE(_0000_),
    .Q(\mem[15][14] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][15]$_DFFE_PP_  (.D(net11),
    .DE(_0000_),
    .Q(\mem[15][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][16]$_DFFE_PP_  (.D(net12),
    .DE(_0000_),
    .Q(\mem[15][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][17]$_DFFE_PP_  (.D(net13),
    .DE(_0000_),
    .Q(\mem[15][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][18]$_DFFE_PP_  (.D(net14),
    .DE(_0000_),
    .Q(\mem[15][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][19]$_DFFE_PP_  (.D(net15),
    .DE(_0000_),
    .Q(\mem[15][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net16),
    .DE(_0000_),
    .Q(\mem[15][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][20]$_DFFE_PP_  (.D(net17),
    .DE(_0000_),
    .Q(\mem[15][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][21]$_DFFE_PP_  (.D(net18),
    .DE(_0000_),
    .Q(\mem[15][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][22]$_DFFE_PP_  (.D(net19),
    .DE(_0000_),
    .Q(\mem[15][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][23]$_DFFE_PP_  (.D(net20),
    .DE(_0000_),
    .Q(\mem[15][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][24]$_DFFE_PP_  (.D(net21),
    .DE(_0000_),
    .Q(\mem[15][24] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][25]$_DFFE_PP_  (.D(net22),
    .DE(_0000_),
    .Q(\mem[15][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][26]$_DFFE_PP_  (.D(net23),
    .DE(_0000_),
    .Q(\mem[15][26] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][27]$_DFFE_PP_  (.D(net24),
    .DE(_0000_),
    .Q(\mem[15][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][28]$_DFFE_PP_  (.D(net25),
    .DE(_0000_),
    .Q(\mem[15][28] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][29]$_DFFE_PP_  (.D(net26),
    .DE(_0000_),
    .Q(\mem[15][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net27),
    .DE(_0000_),
    .Q(\mem[15][2] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][30]$_DFFE_PP_  (.D(net28),
    .DE(_0000_),
    .Q(\mem[15][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][31]$_DFFE_PP_  (.D(net29),
    .DE(_0000_),
    .Q(\mem[15][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net30),
    .DE(_0000_),
    .Q(\mem[15][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net31),
    .DE(_0000_),
    .Q(\mem[15][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net32),
    .DE(_0000_),
    .Q(\mem[15][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net33),
    .DE(_0000_),
    .Q(\mem[15][6] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net34),
    .DE(_0000_),
    .Q(\mem[15][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][8]$_DFFE_PP_  (.D(net35),
    .DE(_0000_),
    .Q(\mem[15][8] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][9]$_DFFE_PP_  (.D(net36),
    .DE(_0000_),
    .Q(\mem[15][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net5),
    .DE(_0014_),
    .Q(\mem[1][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][10]$_DFFE_PP_  (.D(net6),
    .DE(_0014_),
    .Q(\mem[1][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][11]$_DFFE_PP_  (.D(net7),
    .DE(_0014_),
    .Q(\mem[1][11] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][12]$_DFFE_PP_  (.D(net8),
    .DE(_0014_),
    .Q(\mem[1][12] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][13]$_DFFE_PP_  (.D(net9),
    .DE(_0014_),
    .Q(\mem[1][13] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][14]$_DFFE_PP_  (.D(net10),
    .DE(_0014_),
    .Q(\mem[1][14] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][15]$_DFFE_PP_  (.D(net11),
    .DE(_0014_),
    .Q(\mem[1][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][16]$_DFFE_PP_  (.D(net12),
    .DE(_0014_),
    .Q(\mem[1][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][17]$_DFFE_PP_  (.D(net13),
    .DE(_0014_),
    .Q(\mem[1][17] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][18]$_DFFE_PP_  (.D(net14),
    .DE(_0014_),
    .Q(\mem[1][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][19]$_DFFE_PP_  (.D(net15),
    .DE(_0014_),
    .Q(\mem[1][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net16),
    .DE(_0014_),
    .Q(\mem[1][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][20]$_DFFE_PP_  (.D(net17),
    .DE(_0014_),
    .Q(\mem[1][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][21]$_DFFE_PP_  (.D(net18),
    .DE(_0014_),
    .Q(\mem[1][21] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][22]$_DFFE_PP_  (.D(net19),
    .DE(_0014_),
    .Q(\mem[1][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][23]$_DFFE_PP_  (.D(net20),
    .DE(_0014_),
    .Q(\mem[1][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][24]$_DFFE_PP_  (.D(net21),
    .DE(_0014_),
    .Q(\mem[1][24] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][25]$_DFFE_PP_  (.D(net22),
    .DE(_0014_),
    .Q(\mem[1][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][26]$_DFFE_PP_  (.D(net23),
    .DE(_0014_),
    .Q(\mem[1][26] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][27]$_DFFE_PP_  (.D(net24),
    .DE(_0014_),
    .Q(\mem[1][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][28]$_DFFE_PP_  (.D(net25),
    .DE(_0014_),
    .Q(\mem[1][28] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][29]$_DFFE_PP_  (.D(net26),
    .DE(_0014_),
    .Q(\mem[1][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net27),
    .DE(_0014_),
    .Q(\mem[1][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][30]$_DFFE_PP_  (.D(net28),
    .DE(_0014_),
    .Q(\mem[1][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][31]$_DFFE_PP_  (.D(net29),
    .DE(_0014_),
    .Q(\mem[1][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net30),
    .DE(_0014_),
    .Q(\mem[1][3] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net31),
    .DE(_0014_),
    .Q(\mem[1][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net32),
    .DE(_0014_),
    .Q(\mem[1][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net33),
    .DE(_0014_),
    .Q(\mem[1][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net34),
    .DE(_0014_),
    .Q(\mem[1][7] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][8]$_DFFE_PP_  (.D(net35),
    .DE(_0014_),
    .Q(\mem[1][8] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][9]$_DFFE_PP_  (.D(net36),
    .DE(_0014_),
    .Q(\mem[1][9] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net5),
    .DE(_0013_),
    .Q(\mem[2][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][10]$_DFFE_PP_  (.D(net6),
    .DE(_0013_),
    .Q(\mem[2][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][11]$_DFFE_PP_  (.D(net7),
    .DE(_0013_),
    .Q(\mem[2][11] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][12]$_DFFE_PP_  (.D(net8),
    .DE(_0013_),
    .Q(\mem[2][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][13]$_DFFE_PP_  (.D(net9),
    .DE(_0013_),
    .Q(\mem[2][13] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][14]$_DFFE_PP_  (.D(net10),
    .DE(_0013_),
    .Q(\mem[2][14] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][15]$_DFFE_PP_  (.D(net11),
    .DE(_0013_),
    .Q(\mem[2][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][16]$_DFFE_PP_  (.D(net12),
    .DE(_0013_),
    .Q(\mem[2][16] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][17]$_DFFE_PP_  (.D(net13),
    .DE(_0013_),
    .Q(\mem[2][17] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][18]$_DFFE_PP_  (.D(net14),
    .DE(_0013_),
    .Q(\mem[2][18] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][19]$_DFFE_PP_  (.D(net15),
    .DE(_0013_),
    .Q(\mem[2][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net16),
    .DE(_0013_),
    .Q(\mem[2][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][20]$_DFFE_PP_  (.D(net17),
    .DE(_0013_),
    .Q(\mem[2][20] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][21]$_DFFE_PP_  (.D(net18),
    .DE(_0013_),
    .Q(\mem[2][21] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][22]$_DFFE_PP_  (.D(net19),
    .DE(_0013_),
    .Q(\mem[2][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][23]$_DFFE_PP_  (.D(net20),
    .DE(_0013_),
    .Q(\mem[2][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][24]$_DFFE_PP_  (.D(net21),
    .DE(_0013_),
    .Q(\mem[2][24] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][25]$_DFFE_PP_  (.D(net22),
    .DE(_0013_),
    .Q(\mem[2][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][26]$_DFFE_PP_  (.D(net23),
    .DE(_0013_),
    .Q(\mem[2][26] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][27]$_DFFE_PP_  (.D(net24),
    .DE(_0013_),
    .Q(\mem[2][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][28]$_DFFE_PP_  (.D(net25),
    .DE(_0013_),
    .Q(\mem[2][28] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][29]$_DFFE_PP_  (.D(net26),
    .DE(_0013_),
    .Q(\mem[2][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net27),
    .DE(_0013_),
    .Q(\mem[2][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][30]$_DFFE_PP_  (.D(net28),
    .DE(_0013_),
    .Q(\mem[2][30] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][31]$_DFFE_PP_  (.D(net29),
    .DE(_0013_),
    .Q(\mem[2][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net30),
    .DE(_0013_),
    .Q(\mem[2][3] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net31),
    .DE(_0013_),
    .Q(\mem[2][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net32),
    .DE(_0013_),
    .Q(\mem[2][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net33),
    .DE(_0013_),
    .Q(\mem[2][6] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net34),
    .DE(_0013_),
    .Q(\mem[2][7] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][8]$_DFFE_PP_  (.D(net35),
    .DE(_0013_),
    .Q(\mem[2][8] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][9]$_DFFE_PP_  (.D(net36),
    .DE(_0013_),
    .Q(\mem[2][9] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net5),
    .DE(_0012_),
    .Q(\mem[3][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][10]$_DFFE_PP_  (.D(net6),
    .DE(_0012_),
    .Q(\mem[3][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][11]$_DFFE_PP_  (.D(net7),
    .DE(_0012_),
    .Q(\mem[3][11] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][12]$_DFFE_PP_  (.D(net8),
    .DE(_0012_),
    .Q(\mem[3][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][13]$_DFFE_PP_  (.D(net9),
    .DE(_0012_),
    .Q(\mem[3][13] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][14]$_DFFE_PP_  (.D(net10),
    .DE(_0012_),
    .Q(\mem[3][14] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][15]$_DFFE_PP_  (.D(net11),
    .DE(_0012_),
    .Q(\mem[3][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][16]$_DFFE_PP_  (.D(net12),
    .DE(_0012_),
    .Q(\mem[3][16] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][17]$_DFFE_PP_  (.D(net13),
    .DE(_0012_),
    .Q(\mem[3][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][18]$_DFFE_PP_  (.D(net14),
    .DE(_0012_),
    .Q(\mem[3][18] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][19]$_DFFE_PP_  (.D(net15),
    .DE(_0012_),
    .Q(\mem[3][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net16),
    .DE(_0012_),
    .Q(\mem[3][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][20]$_DFFE_PP_  (.D(net17),
    .DE(_0012_),
    .Q(\mem[3][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][21]$_DFFE_PP_  (.D(net18),
    .DE(_0012_),
    .Q(\mem[3][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][22]$_DFFE_PP_  (.D(net19),
    .DE(_0012_),
    .Q(\mem[3][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][23]$_DFFE_PP_  (.D(net20),
    .DE(_0012_),
    .Q(\mem[3][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][24]$_DFFE_PP_  (.D(net21),
    .DE(_0012_),
    .Q(\mem[3][24] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][25]$_DFFE_PP_  (.D(net22),
    .DE(_0012_),
    .Q(\mem[3][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][26]$_DFFE_PP_  (.D(net23),
    .DE(_0012_),
    .Q(\mem[3][26] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][27]$_DFFE_PP_  (.D(net24),
    .DE(_0012_),
    .Q(\mem[3][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][28]$_DFFE_PP_  (.D(net25),
    .DE(_0012_),
    .Q(\mem[3][28] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][29]$_DFFE_PP_  (.D(net26),
    .DE(_0012_),
    .Q(\mem[3][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net27),
    .DE(_0012_),
    .Q(\mem[3][2] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][30]$_DFFE_PP_  (.D(net28),
    .DE(_0012_),
    .Q(\mem[3][30] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][31]$_DFFE_PP_  (.D(net29),
    .DE(_0012_),
    .Q(\mem[3][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net30),
    .DE(_0012_),
    .Q(\mem[3][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net31),
    .DE(_0012_),
    .Q(\mem[3][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net32),
    .DE(_0012_),
    .Q(\mem[3][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net33),
    .DE(_0012_),
    .Q(\mem[3][6] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net34),
    .DE(_0012_),
    .Q(\mem[3][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][8]$_DFFE_PP_  (.D(net35),
    .DE(_0012_),
    .Q(\mem[3][8] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][9]$_DFFE_PP_  (.D(net36),
    .DE(_0012_),
    .Q(\mem[3][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net5),
    .DE(_0011_),
    .Q(\mem[4][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][10]$_DFFE_PP_  (.D(net6),
    .DE(_0011_),
    .Q(\mem[4][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][11]$_DFFE_PP_  (.D(net7),
    .DE(_0011_),
    .Q(\mem[4][11] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][12]$_DFFE_PP_  (.D(net8),
    .DE(_0011_),
    .Q(\mem[4][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][13]$_DFFE_PP_  (.D(net9),
    .DE(_0011_),
    .Q(\mem[4][13] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][14]$_DFFE_PP_  (.D(net10),
    .DE(_0011_),
    .Q(\mem[4][14] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][15]$_DFFE_PP_  (.D(net11),
    .DE(_0011_),
    .Q(\mem[4][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][16]$_DFFE_PP_  (.D(net12),
    .DE(_0011_),
    .Q(\mem[4][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][17]$_DFFE_PP_  (.D(net13),
    .DE(_0011_),
    .Q(\mem[4][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][18]$_DFFE_PP_  (.D(net14),
    .DE(_0011_),
    .Q(\mem[4][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][19]$_DFFE_PP_  (.D(net15),
    .DE(_0011_),
    .Q(\mem[4][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net16),
    .DE(_0011_),
    .Q(\mem[4][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][20]$_DFFE_PP_  (.D(net17),
    .DE(_0011_),
    .Q(\mem[4][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][21]$_DFFE_PP_  (.D(net18),
    .DE(_0011_),
    .Q(\mem[4][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][22]$_DFFE_PP_  (.D(net19),
    .DE(_0011_),
    .Q(\mem[4][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][23]$_DFFE_PP_  (.D(net20),
    .DE(_0011_),
    .Q(\mem[4][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][24]$_DFFE_PP_  (.D(net21),
    .DE(_0011_),
    .Q(\mem[4][24] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][25]$_DFFE_PP_  (.D(net22),
    .DE(_0011_),
    .Q(\mem[4][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][26]$_DFFE_PP_  (.D(net23),
    .DE(_0011_),
    .Q(\mem[4][26] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][27]$_DFFE_PP_  (.D(net24),
    .DE(_0011_),
    .Q(\mem[4][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][28]$_DFFE_PP_  (.D(net25),
    .DE(_0011_),
    .Q(\mem[4][28] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][29]$_DFFE_PP_  (.D(net26),
    .DE(_0011_),
    .Q(\mem[4][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net27),
    .DE(_0011_),
    .Q(\mem[4][2] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][30]$_DFFE_PP_  (.D(net28),
    .DE(_0011_),
    .Q(\mem[4][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][31]$_DFFE_PP_  (.D(net29),
    .DE(_0011_),
    .Q(\mem[4][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net30),
    .DE(_0011_),
    .Q(\mem[4][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net31),
    .DE(_0011_),
    .Q(\mem[4][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net32),
    .DE(_0011_),
    .Q(\mem[4][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net33),
    .DE(_0011_),
    .Q(\mem[4][6] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net34),
    .DE(_0011_),
    .Q(\mem[4][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][8]$_DFFE_PP_  (.D(net35),
    .DE(_0011_),
    .Q(\mem[4][8] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][9]$_DFFE_PP_  (.D(net36),
    .DE(_0011_),
    .Q(\mem[4][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net5),
    .DE(_0010_),
    .Q(\mem[5][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][10]$_DFFE_PP_  (.D(net6),
    .DE(_0010_),
    .Q(\mem[5][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][11]$_DFFE_PP_  (.D(net7),
    .DE(_0010_),
    .Q(\mem[5][11] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][12]$_DFFE_PP_  (.D(net8),
    .DE(_0010_),
    .Q(\mem[5][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][13]$_DFFE_PP_  (.D(net9),
    .DE(_0010_),
    .Q(\mem[5][13] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][14]$_DFFE_PP_  (.D(net10),
    .DE(_0010_),
    .Q(\mem[5][14] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][15]$_DFFE_PP_  (.D(net11),
    .DE(_0010_),
    .Q(\mem[5][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][16]$_DFFE_PP_  (.D(net12),
    .DE(_0010_),
    .Q(\mem[5][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][17]$_DFFE_PP_  (.D(net13),
    .DE(_0010_),
    .Q(\mem[5][17] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][18]$_DFFE_PP_  (.D(net14),
    .DE(_0010_),
    .Q(\mem[5][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][19]$_DFFE_PP_  (.D(net15),
    .DE(_0010_),
    .Q(\mem[5][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net16),
    .DE(_0010_),
    .Q(\mem[5][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][20]$_DFFE_PP_  (.D(net17),
    .DE(_0010_),
    .Q(\mem[5][20] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][21]$_DFFE_PP_  (.D(net18),
    .DE(_0010_),
    .Q(\mem[5][21] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][22]$_DFFE_PP_  (.D(net19),
    .DE(_0010_),
    .Q(\mem[5][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][23]$_DFFE_PP_  (.D(net20),
    .DE(_0010_),
    .Q(\mem[5][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][24]$_DFFE_PP_  (.D(net21),
    .DE(_0010_),
    .Q(\mem[5][24] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][25]$_DFFE_PP_  (.D(net22),
    .DE(_0010_),
    .Q(\mem[5][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][26]$_DFFE_PP_  (.D(net23),
    .DE(_0010_),
    .Q(\mem[5][26] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][27]$_DFFE_PP_  (.D(net24),
    .DE(_0010_),
    .Q(\mem[5][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][28]$_DFFE_PP_  (.D(net25),
    .DE(_0010_),
    .Q(\mem[5][28] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][29]$_DFFE_PP_  (.D(net26),
    .DE(_0010_),
    .Q(\mem[5][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net27),
    .DE(_0010_),
    .Q(\mem[5][2] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][30]$_DFFE_PP_  (.D(net28),
    .DE(_0010_),
    .Q(\mem[5][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][31]$_DFFE_PP_  (.D(net29),
    .DE(_0010_),
    .Q(\mem[5][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net30),
    .DE(_0010_),
    .Q(\mem[5][3] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net31),
    .DE(_0010_),
    .Q(\mem[5][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net32),
    .DE(_0010_),
    .Q(\mem[5][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net33),
    .DE(_0010_),
    .Q(\mem[5][6] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net34),
    .DE(_0010_),
    .Q(\mem[5][7] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][8]$_DFFE_PP_  (.D(net35),
    .DE(_0010_),
    .Q(\mem[5][8] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][9]$_DFFE_PP_  (.D(net36),
    .DE(_0010_),
    .Q(\mem[5][9] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net5),
    .DE(_0009_),
    .Q(\mem[6][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][10]$_DFFE_PP_  (.D(net6),
    .DE(_0009_),
    .Q(\mem[6][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][11]$_DFFE_PP_  (.D(net7),
    .DE(_0009_),
    .Q(\mem[6][11] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][12]$_DFFE_PP_  (.D(net8),
    .DE(_0009_),
    .Q(\mem[6][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][13]$_DFFE_PP_  (.D(net9),
    .DE(_0009_),
    .Q(\mem[6][13] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][14]$_DFFE_PP_  (.D(net10),
    .DE(_0009_),
    .Q(\mem[6][14] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][15]$_DFFE_PP_  (.D(net11),
    .DE(_0009_),
    .Q(\mem[6][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][16]$_DFFE_PP_  (.D(net12),
    .DE(_0009_),
    .Q(\mem[6][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][17]$_DFFE_PP_  (.D(net13),
    .DE(_0009_),
    .Q(\mem[6][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][18]$_DFFE_PP_  (.D(net14),
    .DE(_0009_),
    .Q(\mem[6][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][19]$_DFFE_PP_  (.D(net15),
    .DE(_0009_),
    .Q(\mem[6][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net16),
    .DE(_0009_),
    .Q(\mem[6][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][20]$_DFFE_PP_  (.D(net17),
    .DE(_0009_),
    .Q(\mem[6][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][21]$_DFFE_PP_  (.D(net18),
    .DE(_0009_),
    .Q(\mem[6][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][22]$_DFFE_PP_  (.D(net19),
    .DE(_0009_),
    .Q(\mem[6][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][23]$_DFFE_PP_  (.D(net20),
    .DE(_0009_),
    .Q(\mem[6][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][24]$_DFFE_PP_  (.D(net21),
    .DE(_0009_),
    .Q(\mem[6][24] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][25]$_DFFE_PP_  (.D(net22),
    .DE(_0009_),
    .Q(\mem[6][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][26]$_DFFE_PP_  (.D(net23),
    .DE(_0009_),
    .Q(\mem[6][26] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][27]$_DFFE_PP_  (.D(net24),
    .DE(_0009_),
    .Q(\mem[6][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][28]$_DFFE_PP_  (.D(net25),
    .DE(_0009_),
    .Q(\mem[6][28] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][29]$_DFFE_PP_  (.D(net26),
    .DE(_0009_),
    .Q(\mem[6][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net27),
    .DE(_0009_),
    .Q(\mem[6][2] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][30]$_DFFE_PP_  (.D(net28),
    .DE(_0009_),
    .Q(\mem[6][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][31]$_DFFE_PP_  (.D(net29),
    .DE(_0009_),
    .Q(\mem[6][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net30),
    .DE(_0009_),
    .Q(\mem[6][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net31),
    .DE(_0009_),
    .Q(\mem[6][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net32),
    .DE(_0009_),
    .Q(\mem[6][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net33),
    .DE(_0009_),
    .Q(\mem[6][6] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net34),
    .DE(_0009_),
    .Q(\mem[6][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][8]$_DFFE_PP_  (.D(net35),
    .DE(_0009_),
    .Q(\mem[6][8] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][9]$_DFFE_PP_  (.D(net36),
    .DE(_0009_),
    .Q(\mem[6][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net5),
    .DE(_0008_),
    .Q(\mem[7][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][10]$_DFFE_PP_  (.D(net6),
    .DE(_0008_),
    .Q(\mem[7][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][11]$_DFFE_PP_  (.D(net7),
    .DE(_0008_),
    .Q(\mem[7][11] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][12]$_DFFE_PP_  (.D(net8),
    .DE(_0008_),
    .Q(\mem[7][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][13]$_DFFE_PP_  (.D(net9),
    .DE(_0008_),
    .Q(\mem[7][13] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][14]$_DFFE_PP_  (.D(net10),
    .DE(_0008_),
    .Q(\mem[7][14] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][15]$_DFFE_PP_  (.D(net11),
    .DE(_0008_),
    .Q(\mem[7][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][16]$_DFFE_PP_  (.D(net12),
    .DE(_0008_),
    .Q(\mem[7][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][17]$_DFFE_PP_  (.D(net13),
    .DE(_0008_),
    .Q(\mem[7][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][18]$_DFFE_PP_  (.D(net14),
    .DE(_0008_),
    .Q(\mem[7][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][19]$_DFFE_PP_  (.D(net15),
    .DE(_0008_),
    .Q(\mem[7][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net16),
    .DE(_0008_),
    .Q(\mem[7][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][20]$_DFFE_PP_  (.D(net17),
    .DE(_0008_),
    .Q(\mem[7][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][21]$_DFFE_PP_  (.D(net18),
    .DE(_0008_),
    .Q(\mem[7][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][22]$_DFFE_PP_  (.D(net19),
    .DE(_0008_),
    .Q(\mem[7][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][23]$_DFFE_PP_  (.D(net20),
    .DE(_0008_),
    .Q(\mem[7][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][24]$_DFFE_PP_  (.D(net21),
    .DE(_0008_),
    .Q(\mem[7][24] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][25]$_DFFE_PP_  (.D(net22),
    .DE(_0008_),
    .Q(\mem[7][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][26]$_DFFE_PP_  (.D(net23),
    .DE(_0008_),
    .Q(\mem[7][26] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][27]$_DFFE_PP_  (.D(net24),
    .DE(_0008_),
    .Q(\mem[7][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][28]$_DFFE_PP_  (.D(net25),
    .DE(_0008_),
    .Q(\mem[7][28] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][29]$_DFFE_PP_  (.D(net26),
    .DE(_0008_),
    .Q(\mem[7][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net27),
    .DE(_0008_),
    .Q(\mem[7][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][30]$_DFFE_PP_  (.D(net28),
    .DE(_0008_),
    .Q(\mem[7][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][31]$_DFFE_PP_  (.D(net29),
    .DE(_0008_),
    .Q(\mem[7][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net30),
    .DE(_0008_),
    .Q(\mem[7][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net31),
    .DE(_0008_),
    .Q(\mem[7][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net32),
    .DE(_0008_),
    .Q(\mem[7][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net33),
    .DE(_0008_),
    .Q(\mem[7][6] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net34),
    .DE(_0008_),
    .Q(\mem[7][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][8]$_DFFE_PP_  (.D(net35),
    .DE(_0008_),
    .Q(\mem[7][8] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][9]$_DFFE_PP_  (.D(net36),
    .DE(_0008_),
    .Q(\mem[7][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net5),
    .DE(_0007_),
    .Q(\mem[8][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][10]$_DFFE_PP_  (.D(net6),
    .DE(_0007_),
    .Q(\mem[8][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][11]$_DFFE_PP_  (.D(net7),
    .DE(_0007_),
    .Q(\mem[8][11] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][12]$_DFFE_PP_  (.D(net8),
    .DE(_0007_),
    .Q(\mem[8][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][13]$_DFFE_PP_  (.D(net9),
    .DE(_0007_),
    .Q(\mem[8][13] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][14]$_DFFE_PP_  (.D(net10),
    .DE(_0007_),
    .Q(\mem[8][14] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][15]$_DFFE_PP_  (.D(net11),
    .DE(_0007_),
    .Q(\mem[8][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][16]$_DFFE_PP_  (.D(net12),
    .DE(_0007_),
    .Q(\mem[8][16] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][17]$_DFFE_PP_  (.D(net13),
    .DE(_0007_),
    .Q(\mem[8][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][18]$_DFFE_PP_  (.D(net14),
    .DE(_0007_),
    .Q(\mem[8][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][19]$_DFFE_PP_  (.D(net15),
    .DE(_0007_),
    .Q(\mem[8][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net16),
    .DE(_0007_),
    .Q(\mem[8][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][20]$_DFFE_PP_  (.D(net17),
    .DE(_0007_),
    .Q(\mem[8][20] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][21]$_DFFE_PP_  (.D(net18),
    .DE(_0007_),
    .Q(\mem[8][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][22]$_DFFE_PP_  (.D(net19),
    .DE(_0007_),
    .Q(\mem[8][22] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][23]$_DFFE_PP_  (.D(net20),
    .DE(_0007_),
    .Q(\mem[8][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][24]$_DFFE_PP_  (.D(net21),
    .DE(_0007_),
    .Q(\mem[8][24] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][25]$_DFFE_PP_  (.D(net22),
    .DE(_0007_),
    .Q(\mem[8][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][26]$_DFFE_PP_  (.D(net23),
    .DE(_0007_),
    .Q(\mem[8][26] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][27]$_DFFE_PP_  (.D(net24),
    .DE(_0007_),
    .Q(\mem[8][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][28]$_DFFE_PP_  (.D(net25),
    .DE(_0007_),
    .Q(\mem[8][28] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][29]$_DFFE_PP_  (.D(net26),
    .DE(_0007_),
    .Q(\mem[8][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net27),
    .DE(_0007_),
    .Q(\mem[8][2] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][30]$_DFFE_PP_  (.D(net28),
    .DE(_0007_),
    .Q(\mem[8][30] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][31]$_DFFE_PP_  (.D(net29),
    .DE(_0007_),
    .Q(\mem[8][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net30),
    .DE(_0007_),
    .Q(\mem[8][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net31),
    .DE(_0007_),
    .Q(\mem[8][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net32),
    .DE(_0007_),
    .Q(\mem[8][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net33),
    .DE(_0007_),
    .Q(\mem[8][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net34),
    .DE(_0007_),
    .Q(\mem[8][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][8]$_DFFE_PP_  (.D(net35),
    .DE(_0007_),
    .Q(\mem[8][8] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][9]$_DFFE_PP_  (.D(net36),
    .DE(_0007_),
    .Q(\mem[8][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net5),
    .DE(_0006_),
    .Q(\mem[9][0] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][10]$_DFFE_PP_  (.D(net6),
    .DE(_0006_),
    .Q(\mem[9][10] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][11]$_DFFE_PP_  (.D(net7),
    .DE(_0006_),
    .Q(\mem[9][11] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][12]$_DFFE_PP_  (.D(net8),
    .DE(_0006_),
    .Q(\mem[9][12] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][13]$_DFFE_PP_  (.D(net9),
    .DE(_0006_),
    .Q(\mem[9][13] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][14]$_DFFE_PP_  (.D(net10),
    .DE(_0006_),
    .Q(\mem[9][14] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][15]$_DFFE_PP_  (.D(net11),
    .DE(_0006_),
    .Q(\mem[9][15] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][16]$_DFFE_PP_  (.D(net12),
    .DE(_0006_),
    .Q(\mem[9][16] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][17]$_DFFE_PP_  (.D(net13),
    .DE(_0006_),
    .Q(\mem[9][17] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][18]$_DFFE_PP_  (.D(net14),
    .DE(_0006_),
    .Q(\mem[9][18] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][19]$_DFFE_PP_  (.D(net15),
    .DE(_0006_),
    .Q(\mem[9][19] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net16),
    .DE(_0006_),
    .Q(\mem[9][1] ),
    .CLK(net85));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][20]$_DFFE_PP_  (.D(net17),
    .DE(_0006_),
    .Q(\mem[9][20] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][21]$_DFFE_PP_  (.D(net18),
    .DE(_0006_),
    .Q(\mem[9][21] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][22]$_DFFE_PP_  (.D(net19),
    .DE(_0006_),
    .Q(\mem[9][22] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][23]$_DFFE_PP_  (.D(net20),
    .DE(_0006_),
    .Q(\mem[9][23] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][24]$_DFFE_PP_  (.D(net21),
    .DE(_0006_),
    .Q(\mem[9][24] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][25]$_DFFE_PP_  (.D(net22),
    .DE(_0006_),
    .Q(\mem[9][25] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][26]$_DFFE_PP_  (.D(net23),
    .DE(_0006_),
    .Q(\mem[9][26] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][27]$_DFFE_PP_  (.D(net24),
    .DE(_0006_),
    .Q(\mem[9][27] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][28]$_DFFE_PP_  (.D(net25),
    .DE(_0006_),
    .Q(\mem[9][28] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][29]$_DFFE_PP_  (.D(net26),
    .DE(_0006_),
    .Q(\mem[9][29] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net27),
    .DE(_0006_),
    .Q(\mem[9][2] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][30]$_DFFE_PP_  (.D(net28),
    .DE(_0006_),
    .Q(\mem[9][30] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][31]$_DFFE_PP_  (.D(net29),
    .DE(_0006_),
    .Q(\mem[9][31] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net30),
    .DE(_0006_),
    .Q(\mem[9][3] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net31),
    .DE(_0006_),
    .Q(\mem[9][4] ),
    .CLK(net87));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net32),
    .DE(_0006_),
    .Q(\mem[9][5] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net33),
    .DE(_0006_),
    .Q(\mem[9][6] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net34),
    .DE(_0006_),
    .Q(\mem[9][7] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][8]$_DFFE_PP_  (.D(net35),
    .DE(_0006_),
    .Q(\mem[9][8] ),
    .CLK(net86));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][9]$_DFFE_PP_  (.D(net36),
    .DE(_0006_),
    .Q(\mem[9][9] ),
    .CLK(net86));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[0]$_DFFE_PN0P_  (.D(_0020_),
    .Q(net45),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[10]$_DFFE_PN0P_  (.D(_0021_),
    .Q(net46),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[11]$_DFFE_PN0P_  (.D(_0022_),
    .Q(net47),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[12]$_DFFE_PN0P_  (.D(_0023_),
    .Q(net48),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[13]$_DFFE_PN0P_  (.D(_0024_),
    .Q(net49),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[14]$_DFFE_PN0P_  (.D(_0025_),
    .Q(net50),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[15]$_DFFE_PN0P_  (.D(_0026_),
    .Q(net51),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[16]$_DFFE_PN0P_  (.D(_0027_),
    .Q(net52),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[17]$_DFFE_PN0P_  (.D(_0028_),
    .Q(net53),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[18]$_DFFE_PN0P_  (.D(_0029_),
    .Q(net54),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[19]$_DFFE_PN0P_  (.D(_0030_),
    .Q(net55),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[1]$_DFFE_PN0P_  (.D(_0031_),
    .Q(net56),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[20]$_DFFE_PN0P_  (.D(_0032_),
    .Q(net57),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[21]$_DFFE_PN0P_  (.D(_0033_),
    .Q(net58),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[22]$_DFFE_PN0P_  (.D(_0034_),
    .Q(net59),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[23]$_DFFE_PN0P_  (.D(_0035_),
    .Q(net60),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[24]$_DFFE_PN0P_  (.D(_0036_),
    .Q(net61),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[25]$_DFFE_PN0P_  (.D(_0037_),
    .Q(net62),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[26]$_DFFE_PN0P_  (.D(_0038_),
    .Q(net63),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[27]$_DFFE_PN0P_  (.D(_0039_),
    .Q(net64),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[28]$_DFFE_PN0P_  (.D(_0040_),
    .Q(net65),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[29]$_DFFE_PN0P_  (.D(_0041_),
    .Q(net66),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[2]$_DFFE_PN0P_  (.D(_0042_),
    .Q(net67),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[30]$_DFFE_PN0P_  (.D(_0043_),
    .Q(net68),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[31]$_DFFE_PN0P_  (.D(_0044_),
    .Q(net69),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[3]$_DFFE_PN0P_  (.D(_0045_),
    .Q(net70),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[4]$_DFFE_PN0P_  (.D(_0046_),
    .Q(net71),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[5]$_DFFE_PN0P_  (.D(_0047_),
    .Q(net72),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[6]$_DFFE_PN0P_  (.D(_0048_),
    .Q(net73),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[7]$_DFFE_PN0P_  (.D(_0049_),
    .Q(net74),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[8]$_DFFE_PN0P_  (.D(_0050_),
    .Q(net75),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data[9]$_DFFE_PN0P_  (.D(_0051_),
    .Q(net76),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_4 \rd_ptr_bin[0]$_DFFE_PN0P_  (.D(_0052_),
    .Q(\rd_ptr_bin[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr_bin[1]$_DFFE_PN0P_  (.D(_0053_),
    .Q(\rd_ptr_bin[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[2]$_DFFE_PN0P_  (.D(_0054_),
    .Q(\rd_ptr_bin[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[3]$_DFFE_PN0P_  (.D(_0055_),
    .Q(\rd_ptr_bin[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr_gray[0]$_DFFE_PN0P_  (.D(_0056_),
    .Q(\rd_ptr_gray[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[1]$_DFFE_PN0P_  (.D(_0057_),
    .Q(\rd_ptr_gray[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[2]$_DFFE_PN0P_  (.D(_0058_),
    .Q(\rd_ptr_gray[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[3]$_DFFE_PN0P_  (.D(_0059_),
    .Q(\rd_ptr_gray[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr_gray[4]$_DFFE_PN0P_  (.D(_0060_),
    .Q(\rd_ptr_bin[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\rd_ptr_gray[0] ),
    .Q(\rd_ptr_gray_sync1[0] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\rd_ptr_gray[1] ),
    .Q(\rd_ptr_gray_sync1[1] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\rd_ptr_gray[2] ),
    .Q(\rd_ptr_gray_sync1[2] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\rd_ptr_gray[3] ),
    .Q(\rd_ptr_gray_sync1[3] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\rd_ptr_bin[4] ),
    .Q(\rd_ptr_gray_sync1[4] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[0] ),
    .Q(\rd_ptr_gray_sync2[0] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[1] ),
    .Q(\rd_ptr_gray_sync2[1] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[2] ),
    .Q(\rd_ptr_gray_sync2[2] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[3] ),
    .Q(\rd_ptr_gray_sync2[3] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[4] ),
    .Q(\rd_ptr_gray_sync2[4] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_bin[0]$_DFFE_PN0P_  (.D(_0061_),
    .Q(\wr_ptr_bin[0] ),
    .RESET_B(net38),
    .CLK(net85));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr_bin[1]$_DFFE_PN0P_  (.D(_0062_),
    .Q(\wr_ptr_bin[1] ),
    .RESET_B(net38),
    .CLK(net85));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_bin[2]$_DFFE_PN0P_  (.D(_0063_),
    .Q(\wr_ptr_bin[2] ),
    .RESET_B(net38),
    .CLK(net85));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_bin[3]$_DFFE_PN0P_  (.D(_0064_),
    .Q(\wr_ptr_bin[3] ),
    .RESET_B(net38),
    .CLK(net85));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[0]$_DFFE_PN0P_  (.D(_0065_),
    .Q(\wr_ptr_gray[0] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[1]$_DFFE_PN0P_  (.D(_0066_),
    .Q(\wr_ptr_gray[1] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[2]$_DFFE_PN0P_  (.D(_0067_),
    .Q(\wr_ptr_gray[2] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[3]$_DFFE_PN0P_  (.D(_0068_),
    .Q(\wr_ptr_gray[3] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr_gray[4]$_DFFE_PN0P_  (.D(_0069_),
    .Q(\wr_ptr_bin[4] ),
    .RESET_B(net38),
    .CLK(net87));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\wr_ptr_gray[0] ),
    .Q(\wr_ptr_gray_sync1[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\wr_ptr_gray[1] ),
    .Q(\wr_ptr_gray_sync1[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\wr_ptr_gray[2] ),
    .Q(\wr_ptr_gray_sync1[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\wr_ptr_gray[3] ),
    .Q(\wr_ptr_gray_sync1[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\wr_ptr_bin[4] ),
    .Q(\wr_ptr_gray_sync1[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[0] ),
    .Q(\wr_ptr_gray_sync2[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[1] ),
    .Q(\wr_ptr_gray_sync2[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[2] ),
    .Q(\wr_ptr_gray_sync2[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[3] ),
    .Q(\wr_ptr_gray_sync2[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[4] ),
    .Q(\wr_ptr_gray_sync2[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_531 ();
 sky130_fd_sc_hd__buf_12 input1 (.A(rd_clk),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(rd_en),
    .X(net2));
 sky130_fd_sc_hd__buf_16 input3 (.A(rd_rst_n),
    .X(net3));
 sky130_fd_sc_hd__buf_16 input4 (.A(wr_clk),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(wr_data[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(wr_data[10]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(wr_data[11]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(wr_data[12]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(wr_data[13]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(wr_data[14]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(wr_data[15]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(wr_data[16]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(wr_data[17]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(wr_data[18]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(wr_data[19]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(wr_data[1]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(wr_data[20]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(wr_data[21]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(wr_data[22]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(wr_data[23]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(wr_data[24]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(wr_data[25]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(wr_data[26]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(wr_data[27]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(wr_data[28]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(wr_data[29]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(wr_data[2]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(wr_data[30]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(wr_data[31]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(wr_data[3]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(wr_data[4]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(wr_data[5]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(wr_data[6]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(wr_data[7]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(wr_data[8]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(wr_data[9]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(wr_en),
    .X(net37));
 sky130_fd_sc_hd__buf_12 input38 (.A(wr_rst_n),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net39),
    .X(rd_almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net40),
    .X(rd_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net41),
    .X(rd_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net42),
    .X(rd_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net43),
    .X(rd_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net44),
    .X(rd_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net45),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net46),
    .X(rd_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net47),
    .X(rd_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net48),
    .X(rd_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net49),
    .X(rd_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net50),
    .X(rd_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net51),
    .X(rd_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net52),
    .X(rd_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(rd_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(rd_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(rd_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(rd_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(rd_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(rd_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(rd_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(rd_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(rd_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(rd_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .X(rd_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .X(rd_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(rd_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(rd_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(rd_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(rd_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(rd_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(rd_empty));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(wr_almost_full));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(wr_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(wr_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(wr_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(wr_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(wr_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(wr_full));
 sky130_fd_sc_hd__buf_16 load_slew85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_16 load_slew86 (.A(net4),
    .X(net86));
 sky130_fd_sc_hd__buf_16 load_slew87 (.A(net4),
    .X(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net10));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_314 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_437 ();
endmodule
