module floating_point_adder (clk,
    inexact,
    invalid_op,
    overflow,
    rst_n,
    underflow,
    valid_in,
    valid_out,
    a,
    b,
    result);
 input clk;
 output inexact;
 output invalid_op;
 output overflow;
 input rst_n;
 output underflow;
 input valid_in;
 output valid_out;
 input [31:0] a;
 input [31:0] b;
 output [31:0] result;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire a_sign_stage1;
 wire \add_result[10] ;
 wire \add_result[11] ;
 wire \add_result[12] ;
 wire \add_result[13] ;
 wire \add_result[14] ;
 wire \add_result[15] ;
 wire \add_result[16] ;
 wire \add_result[17] ;
 wire \add_result[18] ;
 wire \add_result[19] ;
 wire \add_result[20] ;
 wire \add_result[21] ;
 wire \add_result[22] ;
 wire \add_result[23] ;
 wire \add_result[24] ;
 wire \add_result[25] ;
 wire \add_result[26] ;
 wire \add_result[2] ;
 wire \add_result[3] ;
 wire \add_result[4] ;
 wire \add_result[5] ;
 wire \add_result[6] ;
 wire \add_result[7] ;
 wire \add_result[8] ;
 wire \add_result[9] ;
 wire \aligned_a_mant[0] ;
 wire \aligned_a_mant[10] ;
 wire \aligned_a_mant[11] ;
 wire \aligned_a_mant[12] ;
 wire \aligned_a_mant[13] ;
 wire \aligned_a_mant[14] ;
 wire \aligned_a_mant[15] ;
 wire \aligned_a_mant[16] ;
 wire \aligned_a_mant[17] ;
 wire \aligned_a_mant[18] ;
 wire \aligned_a_mant[19] ;
 wire \aligned_a_mant[1] ;
 wire \aligned_a_mant[20] ;
 wire \aligned_a_mant[21] ;
 wire \aligned_a_mant[22] ;
 wire \aligned_a_mant[23] ;
 wire \aligned_a_mant[24] ;
 wire \aligned_a_mant[25] ;
 wire \aligned_a_mant[2] ;
 wire \aligned_a_mant[3] ;
 wire \aligned_a_mant[4] ;
 wire \aligned_a_mant[5] ;
 wire \aligned_a_mant[6] ;
 wire \aligned_a_mant[7] ;
 wire \aligned_a_mant[8] ;
 wire \aligned_a_mant[9] ;
 wire \aligned_b_mant[0] ;
 wire \aligned_b_mant[10] ;
 wire \aligned_b_mant[11] ;
 wire \aligned_b_mant[12] ;
 wire \aligned_b_mant[13] ;
 wire \aligned_b_mant[14] ;
 wire \aligned_b_mant[15] ;
 wire \aligned_b_mant[16] ;
 wire \aligned_b_mant[17] ;
 wire \aligned_b_mant[18] ;
 wire \aligned_b_mant[19] ;
 wire \aligned_b_mant[1] ;
 wire \aligned_b_mant[20] ;
 wire \aligned_b_mant[21] ;
 wire \aligned_b_mant[22] ;
 wire \aligned_b_mant[23] ;
 wire \aligned_b_mant[24] ;
 wire \aligned_b_mant[25] ;
 wire \aligned_b_mant[2] ;
 wire \aligned_b_mant[3] ;
 wire \aligned_b_mant[4] ;
 wire \aligned_b_mant[5] ;
 wire \aligned_b_mant[6] ;
 wire \aligned_b_mant[7] ;
 wire \aligned_b_mant[8] ;
 wire \aligned_b_mant[9] ;
 wire b_sign_stage1;
 wire \final_exp[0] ;
 wire \final_exp[1] ;
 wire \final_exp[2] ;
 wire \final_exp[3] ;
 wire \final_exp[4] ;
 wire \final_exp[5] ;
 wire \final_exp[6] ;
 wire \final_exp[7] ;
 wire \final_mant[0] ;
 wire \final_mant[10] ;
 wire \final_mant[11] ;
 wire \final_mant[12] ;
 wire \final_mant[13] ;
 wire \final_mant[14] ;
 wire \final_mant[15] ;
 wire \final_mant[16] ;
 wire \final_mant[17] ;
 wire \final_mant[18] ;
 wire \final_mant[19] ;
 wire \final_mant[1] ;
 wire \final_mant[20] ;
 wire \final_mant[21] ;
 wire \final_mant[22] ;
 wire \final_mant[2] ;
 wire \final_mant[3] ;
 wire \final_mant[4] ;
 wire \final_mant[5] ;
 wire \final_mant[6] ;
 wire \final_mant[7] ;
 wire \final_mant[8] ;
 wire \final_mant[9] ;
 wire inexact_stage2;
 wire invalid_op_stage2;
 wire is_a_larger_stage1;
 wire \larger_exp_stage1[0] ;
 wire \larger_exp_stage1[1] ;
 wire \larger_exp_stage1[2] ;
 wire \larger_exp_stage1[3] ;
 wire \larger_exp_stage1[4] ;
 wire \larger_exp_stage1[5] ;
 wire \larger_exp_stage1[6] ;
 wire \larger_exp_stage1[7] ;
 wire \result_exp_stage2[0] ;
 wire \result_exp_stage2[1] ;
 wire \result_exp_stage2[2] ;
 wire \result_exp_stage2[3] ;
 wire \result_exp_stage2[4] ;
 wire \result_exp_stage2[5] ;
 wire \result_exp_stage2[6] ;
 wire \result_exp_stage2[7] ;
 wire result_sign_stage2;
 wire valid_stage1;
 wire valid_stage2;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 BUF_X4 _2348_ (.A(\add_result[25] ),
    .Z(_1551_));
 INV_X2 _2349_ (.A(_1551_),
    .ZN(_1552_));
 NAND2_X2 _2350_ (.A1(_1552_),
    .A2(_0020_),
    .ZN(_1553_));
 INV_X1 _2351_ (.A(_0021_),
    .ZN(_1554_));
 BUF_X2 _2352_ (.A(_0023_),
    .Z(_1555_));
 INV_X1 _2353_ (.A(\add_result[20] ),
    .ZN(_1556_));
 OAI21_X1 _2354_ (.A(_1555_),
    .B1(\add_result[21] ),
    .B2(_1556_),
    .ZN(_1557_));
 CLKBUF_X2 _2355_ (.A(_0022_),
    .Z(_1558_));
 AOI21_X2 _2356_ (.A(_1554_),
    .B1(_1557_),
    .B2(_1558_),
    .ZN(_1559_));
 NOR2_X4 _2357_ (.A1(_1553_),
    .A2(_1559_),
    .ZN(_1560_));
 CLKBUF_X3 _2358_ (.A(_1560_),
    .Z(_1561_));
 BUF_X4 _2359_ (.A(_1561_),
    .Z(_2125_));
 INV_X1 _2360_ (.A(_1558_),
    .ZN(_1562_));
 NOR2_X1 _2361_ (.A1(\add_result[20] ),
    .A2(\add_result[21] ),
    .ZN(_1563_));
 NOR3_X1 _2362_ (.A1(\add_result[22] ),
    .A2(_1562_),
    .A3(_1563_),
    .ZN(_1564_));
 OR3_X1 _2363_ (.A1(\add_result[24] ),
    .A2(_1553_),
    .A3(_1564_),
    .ZN(_1565_));
 BUF_X2 _2364_ (.A(_1565_),
    .Z(_1566_));
 CLKBUF_X3 _2365_ (.A(_1566_),
    .Z(_1567_));
 CLKBUF_X3 _2366_ (.A(_1567_),
    .Z(_2132_));
 INV_X1 _2367_ (.A(_2132_),
    .ZN(_2004_));
 NOR4_X4 _2368_ (.A1(\add_result[22] ),
    .A2(\add_result[24] ),
    .A3(\add_result[23] ),
    .A4(_1551_),
    .ZN(_1568_));
 NAND2_X1 _2369_ (.A1(_0020_),
    .A2(_1568_),
    .ZN(_1569_));
 INV_X1 _2370_ (.A(_1569_),
    .ZN(_1570_));
 CLKBUF_X3 _2371_ (.A(_1570_),
    .Z(_2136_));
 INV_X1 _2372_ (.A(net38),
    .ZN(_2050_));
 INV_X1 _2373_ (.A(net47),
    .ZN(_2056_));
 INV_X1 _2374_ (.A(net50),
    .ZN(_2053_));
 INV_X1 _2375_ (.A(net51),
    .ZN(_2068_));
 INV_X1 _2376_ (.A(net52),
    .ZN(_2065_));
 BUF_X1 _2377_ (.A(b[6]),
    .Z(_1571_));
 INV_X1 _2378_ (.A(_1571_),
    .ZN(_2062_));
 BUF_X1 _2379_ (.A(b[7]),
    .Z(_1572_));
 INV_X1 _2380_ (.A(_1572_),
    .ZN(_2059_));
 BUF_X1 _2381_ (.A(b[8]),
    .Z(_1573_));
 INV_X1 _2382_ (.A(_1573_),
    .ZN(_2092_));
 BUF_X1 _2383_ (.A(b[9]),
    .Z(_1574_));
 INV_X1 _2384_ (.A(_1574_),
    .ZN(_2089_));
 INV_X1 _2385_ (.A(net34),
    .ZN(_2086_));
 INV_X2 _2386_ (.A(net35),
    .ZN(_2083_));
 INV_X1 _2387_ (.A(net36),
    .ZN(_2080_));
 BUF_X2 _2388_ (.A(b[13]),
    .Z(_1575_));
 INV_X1 _2389_ (.A(_1575_),
    .ZN(_2077_));
 CLKBUF_X2 _2390_ (.A(b[14]),
    .Z(_1576_));
 INV_X1 _2391_ (.A(_1576_),
    .ZN(_2074_));
 INV_X1 _2392_ (.A(net37),
    .ZN(_2071_));
 BUF_X2 _2393_ (.A(b[16]),
    .Z(_1577_));
 INV_X1 _2394_ (.A(_1577_),
    .ZN(_2104_));
 BUF_X2 _2395_ (.A(b[17]),
    .Z(_1578_));
 INV_X1 _2396_ (.A(_1578_),
    .ZN(_2101_));
 BUF_X2 _2397_ (.A(b[18]),
    .Z(_1579_));
 INV_X1 _2398_ (.A(_1579_),
    .ZN(_2098_));
 BUF_X2 _2399_ (.A(b[19]),
    .Z(_1580_));
 INV_X1 _2400_ (.A(_1580_),
    .ZN(_2095_));
 INV_X1 _2401_ (.A(net39),
    .ZN(_2110_));
 BUF_X2 _2402_ (.A(b[21]),
    .Z(_1581_));
 INV_X1 _2403_ (.A(_1581_),
    .ZN(_2107_));
 BUF_X2 _2404_ (.A(b[22]),
    .Z(_1582_));
 INV_X1 _2405_ (.A(_1582_),
    .ZN(_2113_));
 INV_X1 _2406_ (.A(net24),
    .ZN(_2007_));
 INV_X1 _2407_ (.A(net22),
    .ZN(_2013_));
 INV_X1 _2408_ (.A(net21),
    .ZN(_2019_));
 INV_X1 _2409_ (.A(net20),
    .ZN(_2025_));
 INV_X1 _2410_ (.A(net19),
    .ZN(_2031_));
 INV_X1 _2411_ (.A(net18),
    .ZN(_2037_));
 INV_X1 _2412_ (.A(net17),
    .ZN(_1994_));
 INV_X1 _2413_ (.A(net1),
    .ZN(_2047_));
 INV_X1 _2414_ (.A(_2120_),
    .ZN(_1995_));
 INV_X1 _2415_ (.A(_2117_),
    .ZN(_1999_));
 INV_X1 _2416_ (.A(net16),
    .ZN(_2116_));
 INV_X1 _2417_ (.A(net48),
    .ZN(_2010_));
 INV_X1 _2418_ (.A(net46),
    .ZN(_2016_));
 INV_X1 _2419_ (.A(net45),
    .ZN(_2022_));
 INV_X1 _2420_ (.A(net44),
    .ZN(_2028_));
 INV_X1 _2421_ (.A(net43),
    .ZN(_2034_));
 INV_X1 _2422_ (.A(net42),
    .ZN(_2040_));
 INV_X1 _2423_ (.A(net41),
    .ZN(_1998_));
 INV_X1 _2424_ (.A(net40),
    .ZN(_2119_));
 INV_X1 _2425_ (.A(_2125_),
    .ZN(_2127_));
 CLKBUF_X3 _2426_ (.A(_1569_),
    .Z(_1583_));
 CLKBUF_X3 _2427_ (.A(_1583_),
    .Z(_2139_));
 BUF_X1 _2428_ (.A(rst_n),
    .Z(_1584_));
 INV_X2 _2429_ (.A(_1584_),
    .ZN(_1585_));
 BUF_X4 _2430_ (.A(_1585_),
    .Z(_1586_));
 BUF_X4 _2431_ (.A(_1585_),
    .Z(_1587_));
 BUF_X4 _2432_ (.A(\add_result[26] ),
    .Z(_1588_));
 INV_X4 _2433_ (.A(_1588_),
    .ZN(_1589_));
 NOR4_X2 _2434_ (.A1(\add_result[3] ),
    .A2(\add_result[9] ),
    .A3(\add_result[12] ),
    .A4(\add_result[14] ),
    .ZN(_1590_));
 NOR4_X4 _2435_ (.A1(\add_result[13] ),
    .A2(\add_result[16] ),
    .A3(\add_result[15] ),
    .A4(\add_result[18] ),
    .ZN(_1591_));
 NOR3_X2 _2436_ (.A1(\add_result[4] ),
    .A2(\add_result[17] ),
    .A3(\add_result[19] ),
    .ZN(_1592_));
 NAND4_X4 _2437_ (.A1(_1568_),
    .A2(_1590_),
    .A3(_1591_),
    .A4(_1592_),
    .ZN(_1593_));
 NOR4_X2 _2438_ (.A1(\add_result[5] ),
    .A2(\add_result[8] ),
    .A3(\add_result[7] ),
    .A4(\add_result[10] ),
    .ZN(_1594_));
 NOR2_X1 _2439_ (.A1(\add_result[6] ),
    .A2(\add_result[11] ),
    .ZN(_1595_));
 NAND3_X2 _2440_ (.A1(_1563_),
    .A2(_1594_),
    .A3(_1595_),
    .ZN(_1596_));
 OAI21_X4 _2441_ (.A(_1589_),
    .B1(_1593_),
    .B2(_1596_),
    .ZN(_1597_));
 NOR2_X2 _2442_ (.A1(_1587_),
    .A2(_1597_),
    .ZN(_1598_));
 BUF_X4 _2443_ (.A(\result_exp_stage2[3] ),
    .Z(_1599_));
 INV_X2 _2444_ (.A(_2142_),
    .ZN(_1600_));
 NOR3_X4 _2445_ (.A1(_1599_),
    .A2(\result_exp_stage2[2] ),
    .A3(_1600_),
    .ZN(_1601_));
 BUF_X4 _2446_ (.A(\result_exp_stage2[7] ),
    .Z(_1602_));
 BUF_X4 _2447_ (.A(\result_exp_stage2[6] ),
    .Z(_1603_));
 BUF_X4 _2448_ (.A(\result_exp_stage2[5] ),
    .Z(_1604_));
 BUF_X4 _2449_ (.A(\result_exp_stage2[4] ),
    .Z(_1605_));
 NOR4_X4 _2450_ (.A1(_1602_),
    .A2(_1603_),
    .A3(_1604_),
    .A4(_1605_),
    .ZN(_1606_));
 INV_X2 _2451_ (.A(_1599_),
    .ZN(_1607_));
 NAND2_X1 _2452_ (.A1(_1607_),
    .A2(_2137_),
    .ZN(_1608_));
 INV_X1 _2453_ (.A(_2131_),
    .ZN(_1609_));
 INV_X1 _2454_ (.A(_2126_),
    .ZN(_1610_));
 AOI21_X1 _2455_ (.A(_1609_),
    .B1(_2128_),
    .B2(_1610_),
    .ZN(_1611_));
 NOR2_X1 _2456_ (.A1(_2130_),
    .A2(_1611_),
    .ZN(_1612_));
 BUF_X1 _2457_ (.A(_2138_),
    .Z(_1613_));
 NAND2_X1 _2458_ (.A1(_0024_),
    .A2(_1613_),
    .ZN(_1614_));
 OAI21_X2 _2459_ (.A(_1608_),
    .B1(_1612_),
    .B2(_1614_),
    .ZN(_1615_));
 AND2_X1 _2460_ (.A1(_1606_),
    .A2(_1615_),
    .ZN(_1616_));
 BUF_X4 _2461_ (.A(_1616_),
    .Z(_1617_));
 AOI21_X4 _2462_ (.A(_1551_),
    .B1(_1601_),
    .B2(_1617_),
    .ZN(_1618_));
 BUF_X4 _2463_ (.A(_1618_),
    .Z(_1619_));
 CLKBUF_X3 _2464_ (.A(\result_exp_stage2[0] ),
    .Z(_1620_));
 MUX2_X1 _2465_ (.A(_0006_),
    .B(_0007_),
    .S(_1620_),
    .Z(_1621_));
 CLKBUF_X3 _2466_ (.A(_1620_),
    .Z(_1622_));
 MUX2_X1 _2467_ (.A(_0004_),
    .B(_0005_),
    .S(_1622_),
    .Z(_1623_));
 CLKBUF_X3 _2468_ (.A(_2143_),
    .Z(_1624_));
 INV_X1 _2469_ (.A(_1624_),
    .ZN(_1625_));
 CLKBUF_X3 _2470_ (.A(_1625_),
    .Z(_1626_));
 MUX2_X1 _2471_ (.A(_1621_),
    .B(_1623_),
    .S(_1626_),
    .Z(_1627_));
 BUF_X4 _2472_ (.A(\result_exp_stage2[2] ),
    .Z(_1628_));
 XNOR2_X2 _2473_ (.A(_1628_),
    .B(_2142_),
    .ZN(_1629_));
 BUF_X4 _2474_ (.A(_1629_),
    .Z(_1630_));
 AND2_X1 _2475_ (.A1(_1627_),
    .A2(_1630_),
    .ZN(_1631_));
 BUF_X1 _2476_ (.A(_0002_),
    .Z(_1632_));
 CLKBUF_X2 _2477_ (.A(_0003_),
    .Z(_1633_));
 MUX2_X1 _2478_ (.A(_1632_),
    .B(_1633_),
    .S(_1622_),
    .Z(_1634_));
 BUF_X2 _2479_ (.A(_0000_),
    .Z(_1635_));
 BUF_X2 _2480_ (.A(_0001_),
    .Z(_1636_));
 MUX2_X1 _2481_ (.A(_1635_),
    .B(_1636_),
    .S(_1620_),
    .Z(_1637_));
 MUX2_X1 _2482_ (.A(_1634_),
    .B(_1637_),
    .S(_1625_),
    .Z(_1638_));
 XOR2_X2 _2483_ (.A(_1628_),
    .B(_2142_),
    .Z(_1639_));
 CLKBUF_X3 _2484_ (.A(_1639_),
    .Z(_1640_));
 INV_X2 _2485_ (.A(_1604_),
    .ZN(_1641_));
 INV_X2 _2486_ (.A(_1603_),
    .ZN(_1642_));
 OR4_X2 _2487_ (.A1(_1605_),
    .A2(_1599_),
    .A3(_1628_),
    .A4(_1600_),
    .ZN(_1643_));
 NOR3_X2 _2488_ (.A1(_1602_),
    .A2(_1642_),
    .A3(_1643_),
    .ZN(_1644_));
 NOR4_X4 _2489_ (.A1(_1605_),
    .A2(_1599_),
    .A3(_1628_),
    .A4(_1600_),
    .ZN(_1645_));
 NAND2_X1 _2490_ (.A1(_1602_),
    .A2(_1642_),
    .ZN(_1646_));
 NOR2_X2 _2491_ (.A1(_1605_),
    .A2(_1599_),
    .ZN(_1647_));
 NOR3_X4 _2492_ (.A1(\result_exp_stage2[2] ),
    .A2(\result_exp_stage2[1] ),
    .A3(_1620_),
    .ZN(_1648_));
 NAND2_X4 _2493_ (.A1(_1647_),
    .A2(_1648_),
    .ZN(_1649_));
 NOR3_X2 _2494_ (.A1(_1645_),
    .A2(_1646_),
    .A3(_1649_),
    .ZN(_1650_));
 OAI21_X4 _2495_ (.A(_1641_),
    .B1(_1644_),
    .B2(_1650_),
    .ZN(_1651_));
 AOI21_X4 _2496_ (.A(_1604_),
    .B1(_1643_),
    .B2(_1649_),
    .ZN(_1652_));
 OR3_X4 _2497_ (.A1(_1602_),
    .A2(_1603_),
    .A3(_1652_),
    .ZN(_1653_));
 AOI221_X2 _2498_ (.A(_1631_),
    .B1(_1638_),
    .B2(_1640_),
    .C1(_1651_),
    .C2(_1653_),
    .ZN(_1654_));
 XNOR2_X2 _2499_ (.A(_1607_),
    .B(_1648_),
    .ZN(_1655_));
 XNOR2_X2 _2500_ (.A(_1605_),
    .B(_1601_),
    .ZN(_1656_));
 XNOR2_X2 _2501_ (.A(_1641_),
    .B(_1649_),
    .ZN(_1657_));
 NAND2_X2 _2502_ (.A1(_1656_),
    .A2(_1657_),
    .ZN(_1658_));
 NOR2_X2 _2503_ (.A1(_1655_),
    .A2(_1658_),
    .ZN(_1659_));
 NAND2_X1 _2504_ (.A1(_1617_),
    .A2(_1659_),
    .ZN(_1660_));
 INV_X1 _2505_ (.A(_1660_),
    .ZN(_1661_));
 MUX2_X1 _2506_ (.A(_0005_),
    .B(_0007_),
    .S(_1567_),
    .Z(_1662_));
 MUX2_X1 _2507_ (.A(_0004_),
    .B(_0006_),
    .S(_1566_),
    .Z(_1663_));
 MUX2_X1 _2508_ (.A(_1662_),
    .B(_1663_),
    .S(_1561_),
    .Z(_1664_));
 OR2_X1 _2509_ (.A1(_2136_),
    .A2(_1664_),
    .ZN(_1665_));
 MUX2_X1 _2510_ (.A(_1636_),
    .B(_1633_),
    .S(_1566_),
    .Z(_1666_));
 MUX2_X1 _2511_ (.A(_1635_),
    .B(_1632_),
    .S(_1566_),
    .Z(_1667_));
 MUX2_X1 _2512_ (.A(_1666_),
    .B(_1667_),
    .S(_1560_),
    .Z(_1668_));
 OAI21_X1 _2513_ (.A(_1665_),
    .B1(_1668_),
    .B2(_2139_),
    .ZN(_1669_));
 NAND2_X4 _2514_ (.A1(_1606_),
    .A2(_1615_),
    .ZN(_1670_));
 BUF_X4 _2515_ (.A(_1670_),
    .Z(_1671_));
 AOI22_X2 _2516_ (.A1(_1654_),
    .A2(_1661_),
    .B1(_1669_),
    .B2(_1671_),
    .ZN(_1672_));
 BUF_X4 _2517_ (.A(_1551_),
    .Z(_1673_));
 CLKBUF_X3 _2518_ (.A(_1673_),
    .Z(_1674_));
 OAI22_X2 _2519_ (.A1(_0007_),
    .A2(_1619_),
    .B1(_1672_),
    .B2(_1674_),
    .ZN(_1675_));
 NOR2_X1 _2520_ (.A1(_1587_),
    .A2(_1589_),
    .ZN(_1676_));
 BUF_X4 _2521_ (.A(_1676_),
    .Z(_1677_));
 AOI222_X2 _2522_ (.A1(_1586_),
    .A2(\final_mant[7] ),
    .B1(_1598_),
    .B2(_1675_),
    .C1(_1677_),
    .C2(\add_result[10] ),
    .ZN(_1678_));
 INV_X1 _2523_ (.A(_1678_),
    .ZN(_0025_));
 BUF_X4 _2524_ (.A(_1588_),
    .Z(_1679_));
 NOR2_X2 _2525_ (.A1(_1593_),
    .A2(_1596_),
    .ZN(_1680_));
 NOR2_X4 _2526_ (.A1(_1588_),
    .A2(_1680_),
    .ZN(_1681_));
 NAND2_X4 _2527_ (.A1(_1651_),
    .A2(_1653_),
    .ZN(_1682_));
 XNOR2_X2 _2528_ (.A(_1599_),
    .B(_1648_),
    .ZN(_1683_));
 MUX2_X1 _2529_ (.A(_1633_),
    .B(_0004_),
    .S(_1622_),
    .Z(_1684_));
 OR2_X1 _2530_ (.A1(_1626_),
    .A2(_1684_),
    .ZN(_1685_));
 CLKBUF_X3 _2531_ (.A(_1620_),
    .Z(_1686_));
 MUX2_X1 _2532_ (.A(_1636_),
    .B(_1632_),
    .S(_1686_),
    .Z(_1687_));
 CLKBUF_X3 _2533_ (.A(_1624_),
    .Z(_1688_));
 OAI21_X2 _2534_ (.A(_1685_),
    .B1(_1687_),
    .B2(_1688_),
    .ZN(_1689_));
 NAND3_X1 _2535_ (.A1(_1640_),
    .A2(_1683_),
    .A3(_1689_),
    .ZN(_1690_));
 MUX2_X1 _2536_ (.A(_0007_),
    .B(_0008_),
    .S(_1622_),
    .Z(_1691_));
 MUX2_X1 _2537_ (.A(_0005_),
    .B(_0006_),
    .S(_1622_),
    .Z(_1692_));
 MUX2_X1 _2538_ (.A(_1691_),
    .B(_1692_),
    .S(_1626_),
    .Z(_1693_));
 NOR2_X1 _2539_ (.A1(_1655_),
    .A2(_1693_),
    .ZN(_1694_));
 OR2_X1 _2540_ (.A1(_2124_),
    .A2(_1626_),
    .ZN(_1695_));
 NOR2_X1 _2541_ (.A1(_1635_),
    .A2(_1695_),
    .ZN(_1696_));
 AOI21_X1 _2542_ (.A(_1694_),
    .B1(_1696_),
    .B2(_1655_),
    .ZN(_1697_));
 CLKBUF_X3 _2543_ (.A(_1640_),
    .Z(_1698_));
 OAI21_X1 _2544_ (.A(_1690_),
    .B1(_1697_),
    .B2(_1698_),
    .ZN(_1699_));
 NAND2_X1 _2545_ (.A1(_1682_),
    .A2(_1699_),
    .ZN(_1700_));
 AND2_X1 _2546_ (.A1(_1656_),
    .A2(_1657_),
    .ZN(_1701_));
 NAND2_X2 _2547_ (.A1(_1617_),
    .A2(_1701_),
    .ZN(_1702_));
 MUX2_X1 _2548_ (.A(_1632_),
    .B(_0004_),
    .S(_1567_),
    .Z(_1703_));
 MUX2_X1 _2549_ (.A(_1703_),
    .B(_1666_),
    .S(_1560_),
    .Z(_1704_));
 MUX2_X1 _2550_ (.A(_0006_),
    .B(_0008_),
    .S(_1567_),
    .Z(_1705_));
 MUX2_X1 _2551_ (.A(_1705_),
    .B(_1662_),
    .S(_1561_),
    .Z(_1706_));
 MUX2_X1 _2552_ (.A(_1704_),
    .B(_1706_),
    .S(_1569_),
    .Z(_1707_));
 CLKBUF_X3 _2553_ (.A(_1617_),
    .Z(_1708_));
 OAI22_X1 _2554_ (.A1(_1700_),
    .A2(_1702_),
    .B1(_1707_),
    .B2(_1708_),
    .ZN(_1709_));
 NAND2_X1 _2555_ (.A1(_1552_),
    .A2(_1709_),
    .ZN(_1710_));
 OAI21_X1 _2556_ (.A(_1710_),
    .B1(_1619_),
    .B2(_0008_),
    .ZN(_1711_));
 AOI221_X2 _2557_ (.A(_1586_),
    .B1(_1679_),
    .B2(\add_result[11] ),
    .C1(_1681_),
    .C2(_1711_),
    .ZN(_1712_));
 INV_X1 _2558_ (.A(\final_mant[8] ),
    .ZN(_1713_));
 CLKBUF_X3 _2559_ (.A(_1586_),
    .Z(_1714_));
 AOI21_X1 _2560_ (.A(_1712_),
    .B1(_1713_),
    .B2(_1714_),
    .ZN(_0026_));
 NAND2_X1 _2561_ (.A1(_1679_),
    .A2(\add_result[12] ),
    .ZN(_1715_));
 NOR2_X1 _2562_ (.A1(_0009_),
    .A2(_1619_),
    .ZN(_1716_));
 NOR2_X1 _2563_ (.A1(_1626_),
    .A2(_1637_),
    .ZN(_1717_));
 NOR3_X4 _2564_ (.A1(_1602_),
    .A2(_1603_),
    .A3(_1652_),
    .ZN(_1718_));
 INV_X1 _2565_ (.A(_1602_),
    .ZN(_1719_));
 NAND3_X2 _2566_ (.A1(_1719_),
    .A2(_1603_),
    .A3(_1645_),
    .ZN(_1720_));
 OR3_X2 _2567_ (.A1(_1645_),
    .A2(_1646_),
    .A3(_1649_),
    .ZN(_1721_));
 AOI21_X4 _2568_ (.A(_1604_),
    .B1(_1720_),
    .B2(_1721_),
    .ZN(_1722_));
 OAI21_X4 _2569_ (.A(_1717_),
    .B1(_1718_),
    .B2(_1722_),
    .ZN(_1723_));
 NOR3_X1 _2570_ (.A1(_1698_),
    .A2(_1683_),
    .A3(_1723_),
    .ZN(_1724_));
 MUX2_X1 _2571_ (.A(_0008_),
    .B(_0009_),
    .S(_1620_),
    .Z(_1725_));
 MUX2_X1 _2572_ (.A(_1621_),
    .B(_1725_),
    .S(_1624_),
    .Z(_1726_));
 AND2_X1 _2573_ (.A1(_1630_),
    .A2(_1726_),
    .ZN(_1727_));
 MUX2_X1 _2574_ (.A(_1623_),
    .B(_1634_),
    .S(_1626_),
    .Z(_1728_));
 AOI221_X2 _2575_ (.A(_1727_),
    .B1(_1728_),
    .B2(_1640_),
    .C1(_1651_),
    .C2(_1653_),
    .ZN(_1729_));
 AOI21_X1 _2576_ (.A(_1724_),
    .B1(_1729_),
    .B2(_1683_),
    .ZN(_1730_));
 MUX2_X1 _2577_ (.A(_1633_),
    .B(_0005_),
    .S(_1566_),
    .Z(_1731_));
 MUX2_X1 _2578_ (.A(_1731_),
    .B(_1703_),
    .S(_1560_),
    .Z(_1732_));
 MUX2_X1 _2579_ (.A(_0007_),
    .B(_0009_),
    .S(_1566_),
    .Z(_1733_));
 MUX2_X1 _2580_ (.A(_1733_),
    .B(_1705_),
    .S(_1561_),
    .Z(_1734_));
 MUX2_X1 _2581_ (.A(_1732_),
    .B(_1734_),
    .S(_1583_),
    .Z(_1735_));
 OAI22_X1 _2582_ (.A1(_1702_),
    .A2(_1730_),
    .B1(_1735_),
    .B2(_1708_),
    .ZN(_1736_));
 CLKBUF_X3 _2583_ (.A(_1552_),
    .Z(_1737_));
 AOI21_X1 _2584_ (.A(_1716_),
    .B1(_1736_),
    .B2(_1737_),
    .ZN(_1738_));
 OAI21_X1 _2585_ (.A(_1715_),
    .B1(_1738_),
    .B2(_1597_),
    .ZN(_1739_));
 BUF_X4 _2586_ (.A(_1584_),
    .Z(_1740_));
 BUF_X4 _2587_ (.A(_1740_),
    .Z(_1741_));
 MUX2_X1 _2588_ (.A(\final_mant[9] ),
    .B(_1739_),
    .S(_1741_),
    .Z(_0027_));
 INV_X2 _2589_ (.A(_1605_),
    .ZN(_1742_));
 NOR4_X4 _2590_ (.A1(_1642_),
    .A2(_1641_),
    .A3(_1742_),
    .A4(_1607_),
    .ZN(_1743_));
 NAND4_X4 _2591_ (.A1(_1602_),
    .A2(_1628_),
    .A3(_2144_),
    .A4(_1743_),
    .ZN(_1744_));
 NAND3_X1 _2592_ (.A1(_2124_),
    .A2(_1677_),
    .A3(_1744_),
    .ZN(_1745_));
 BUF_X4 _2593_ (.A(_1673_),
    .Z(_1746_));
 OAI21_X4 _2594_ (.A(_1598_),
    .B1(_1671_),
    .B2(_1746_),
    .ZN(_1747_));
 MUX2_X1 _2595_ (.A(_2126_),
    .B(_2124_),
    .S(_1674_),
    .Z(_1748_));
 INV_X1 _2596_ (.A(\final_exp[0] ),
    .ZN(_1749_));
 BUF_X2 _2597_ (.A(_1740_),
    .Z(_1750_));
 OAI221_X1 _2598_ (.A(_1745_),
    .B1(_1747_),
    .B2(_1748_),
    .C1(_1749_),
    .C2(_1750_),
    .ZN(_0166_));
 CLKBUF_X3 _2599_ (.A(_1586_),
    .Z(_1751_));
 AOI22_X1 _2600_ (.A1(_1751_),
    .A2(\final_exp[1] ),
    .B1(_1677_),
    .B2(_1688_),
    .ZN(_1752_));
 NAND2_X1 _2601_ (.A1(_1746_),
    .A2(_2002_),
    .ZN(_1753_));
 OAI21_X1 _2602_ (.A(_1753_),
    .B1(_2006_),
    .B2(_1746_),
    .ZN(_1754_));
 OAI21_X1 _2603_ (.A(_1752_),
    .B1(_1754_),
    .B2(_1747_),
    .ZN(_0167_));
 AND2_X1 _2604_ (.A1(_1628_),
    .A2(_2146_),
    .ZN(_1755_));
 NOR2_X1 _2605_ (.A1(_1628_),
    .A2(_2146_),
    .ZN(_1756_));
 OAI21_X1 _2606_ (.A(_1744_),
    .B1(_1755_),
    .B2(_1756_),
    .ZN(_1757_));
 NAND3_X1 _2607_ (.A1(_1741_),
    .A2(_1679_),
    .A3(_1757_),
    .ZN(_1758_));
 XOR2_X1 _2608_ (.A(_2005_),
    .B(_1613_),
    .Z(_1759_));
 MUX2_X1 _2609_ (.A(_2135_),
    .B(_1759_),
    .S(_1737_),
    .Z(_1760_));
 INV_X1 _2610_ (.A(\final_exp[2] ),
    .ZN(_1761_));
 OAI221_X1 _2611_ (.A(_1758_),
    .B1(_1760_),
    .B2(_1747_),
    .C1(_1761_),
    .C2(_1750_),
    .ZN(_0168_));
 NAND3_X1 _2612_ (.A1(_1628_),
    .A2(\result_exp_stage2[1] ),
    .A3(_1686_),
    .ZN(_1762_));
 XNOR2_X1 _2613_ (.A(_1607_),
    .B(_1762_),
    .ZN(_1763_));
 AOI21_X1 _2614_ (.A(_1589_),
    .B1(_1744_),
    .B2(_1763_),
    .ZN(_1764_));
 NAND2_X1 _2615_ (.A1(_1741_),
    .A2(_1764_),
    .ZN(_1765_));
 INV_X1 _2616_ (.A(_2133_),
    .ZN(_1766_));
 OAI21_X1 _2617_ (.A(_1766_),
    .B1(_1609_),
    .B2(_2003_),
    .ZN(_1767_));
 AOI21_X1 _2618_ (.A(_2140_),
    .B1(_1613_),
    .B2(_1767_),
    .ZN(_1768_));
 XNOR2_X1 _2619_ (.A(_1599_),
    .B(_1768_),
    .ZN(_1769_));
 MUX2_X1 _2620_ (.A(_0024_),
    .B(_1769_),
    .S(_1737_),
    .Z(_1770_));
 INV_X1 _2621_ (.A(\final_exp[3] ),
    .ZN(_1771_));
 OAI221_X1 _2622_ (.A(_1765_),
    .B1(_1770_),
    .B2(_1747_),
    .C1(_1771_),
    .C2(_1750_),
    .ZN(_0169_));
 NAND2_X1 _2623_ (.A1(_1599_),
    .A2(_1755_),
    .ZN(_1772_));
 XNOR2_X1 _2624_ (.A(_1742_),
    .B(_1772_),
    .ZN(_1773_));
 AOI21_X1 _2625_ (.A(_1589_),
    .B1(_1744_),
    .B2(_1773_),
    .ZN(_1774_));
 NAND2_X1 _2626_ (.A1(_1741_),
    .A2(_1774_),
    .ZN(_1775_));
 INV_X1 _2627_ (.A(_0024_),
    .ZN(_1776_));
 NOR3_X1 _2628_ (.A1(_1673_),
    .A2(_1776_),
    .A3(_2140_),
    .ZN(_1777_));
 INV_X1 _2629_ (.A(_1613_),
    .ZN(_1778_));
 OAI21_X1 _2630_ (.A(_1777_),
    .B1(_1778_),
    .B2(_2005_),
    .ZN(_1779_));
 XNOR2_X1 _2631_ (.A(_1742_),
    .B(_1779_),
    .ZN(_1780_));
 INV_X1 _2632_ (.A(\final_exp[4] ),
    .ZN(_1781_));
 OAI221_X1 _2633_ (.A(_1775_),
    .B1(_1780_),
    .B2(_1747_),
    .C1(_1750_),
    .C2(_1781_),
    .ZN(_0170_));
 NOR3_X1 _2634_ (.A1(_1742_),
    .A2(_1607_),
    .A3(_1762_),
    .ZN(_1782_));
 XNOR2_X1 _2635_ (.A(_1604_),
    .B(_1782_),
    .ZN(_1783_));
 AOI21_X1 _2636_ (.A(_1589_),
    .B1(_1744_),
    .B2(_1783_),
    .ZN(_1784_));
 NAND2_X1 _2637_ (.A1(_1741_),
    .A2(_1784_),
    .ZN(_1785_));
 AND3_X1 _2638_ (.A1(_1552_),
    .A2(_1647_),
    .A3(_1768_),
    .ZN(_1786_));
 XNOR2_X1 _2639_ (.A(_1604_),
    .B(_1786_),
    .ZN(_1787_));
 INV_X1 _2640_ (.A(\final_exp[5] ),
    .ZN(_1788_));
 OAI221_X1 _2641_ (.A(_1785_),
    .B1(_1787_),
    .B2(_1747_),
    .C1(_1750_),
    .C2(_1788_),
    .ZN(_0171_));
 NAND4_X1 _2642_ (.A1(_1604_),
    .A2(_1605_),
    .A3(_1599_),
    .A4(_1755_),
    .ZN(_1789_));
 XNOR2_X1 _2643_ (.A(_1642_),
    .B(_1789_),
    .ZN(_1790_));
 NAND2_X1 _2644_ (.A1(_1744_),
    .A2(_1790_),
    .ZN(_1791_));
 AOI22_X1 _2645_ (.A1(_1751_),
    .A2(\final_exp[6] ),
    .B1(_1677_),
    .B2(_1791_),
    .ZN(_1792_));
 NOR3_X1 _2646_ (.A1(_1604_),
    .A2(_1605_),
    .A3(_1779_),
    .ZN(_1793_));
 XNOR2_X1 _2647_ (.A(_1603_),
    .B(_1793_),
    .ZN(_1794_));
 OAI21_X1 _2648_ (.A(_1792_),
    .B1(_1794_),
    .B2(_1747_),
    .ZN(_0172_));
 NAND4_X1 _2649_ (.A1(_1628_),
    .A2(\result_exp_stage2[1] ),
    .A3(_1686_),
    .A4(_1743_),
    .ZN(_1795_));
 XNOR2_X1 _2650_ (.A(_1719_),
    .B(_1795_),
    .ZN(_1796_));
 NAND2_X1 _2651_ (.A1(_1744_),
    .A2(_1796_),
    .ZN(_1797_));
 AOI22_X1 _2652_ (.A1(_1751_),
    .A2(\final_exp[7] ),
    .B1(_1677_),
    .B2(_1797_),
    .ZN(_1798_));
 NAND3_X1 _2653_ (.A1(_1642_),
    .A2(_1641_),
    .A3(_1786_),
    .ZN(_1799_));
 XNOR2_X1 _2654_ (.A(_1719_),
    .B(_1799_),
    .ZN(_1800_));
 OAI21_X1 _2655_ (.A(_1798_),
    .B1(_1800_),
    .B2(_1747_),
    .ZN(_0173_));
 NAND2_X1 _2656_ (.A1(_1751_),
    .A2(\final_mant[0] ),
    .ZN(_1801_));
 NAND2_X2 _2657_ (.A1(_1601_),
    .A2(_1606_),
    .ZN(_1802_));
 NOR2_X1 _2658_ (.A1(_1722_),
    .A2(_1718_),
    .ZN(_1803_));
 BUF_X4 _2659_ (.A(_1803_),
    .Z(_1804_));
 NAND3_X2 _2660_ (.A1(_1629_),
    .A2(_1683_),
    .A3(_1701_),
    .ZN(_1805_));
 OR3_X1 _2661_ (.A1(_1804_),
    .A2(_1695_),
    .A3(_1805_),
    .ZN(_1806_));
 AOI21_X1 _2662_ (.A(_1671_),
    .B1(_1802_),
    .B2(_1806_),
    .ZN(_1807_));
 NAND2_X1 _2663_ (.A1(_2127_),
    .A2(_2132_),
    .ZN(_1808_));
 NOR3_X1 _2664_ (.A1(_2136_),
    .A2(_1708_),
    .A3(_1808_),
    .ZN(_1809_));
 NOR3_X1 _2665_ (.A1(_1674_),
    .A2(_1807_),
    .A3(_1809_),
    .ZN(_1810_));
 NOR3_X1 _2666_ (.A1(_1635_),
    .A2(_1597_),
    .A3(_1810_),
    .ZN(_1811_));
 AOI21_X1 _2667_ (.A(_1811_),
    .B1(\add_result[3] ),
    .B2(_1679_),
    .ZN(_1812_));
 BUF_X4 _2668_ (.A(_1586_),
    .Z(_1813_));
 OAI21_X1 _2669_ (.A(_1801_),
    .B1(_1812_),
    .B2(_1813_),
    .ZN(_0174_));
 NOR2_X2 _2670_ (.A1(_1670_),
    .A2(_1658_),
    .ZN(_1814_));
 CLKBUF_X3 _2671_ (.A(_1655_),
    .Z(_1815_));
 MUX2_X1 _2672_ (.A(_0009_),
    .B(_0010_),
    .S(_1622_),
    .Z(_1816_));
 MUX2_X1 _2673_ (.A(_1691_),
    .B(_1816_),
    .S(_1624_),
    .Z(_1817_));
 NAND2_X1 _2674_ (.A1(_1630_),
    .A2(_1817_),
    .ZN(_1818_));
 MUX2_X1 _2675_ (.A(_1692_),
    .B(_1684_),
    .S(_1626_),
    .Z(_1819_));
 NAND2_X1 _2676_ (.A1(_1640_),
    .A2(_1819_),
    .ZN(_1820_));
 NAND3_X1 _2677_ (.A1(_1682_),
    .A2(_1818_),
    .A3(_1820_),
    .ZN(_1821_));
 NOR2_X1 _2678_ (.A1(_1626_),
    .A2(_1687_),
    .ZN(_1822_));
 NOR3_X2 _2679_ (.A1(_2124_),
    .A2(_1624_),
    .A3(_1635_),
    .ZN(_1823_));
 OAI22_X4 _2680_ (.A1(_1722_),
    .A2(_1718_),
    .B1(_1822_),
    .B2(_1823_),
    .ZN(_1824_));
 BUF_X2 _2681_ (.A(_1630_),
    .Z(_1825_));
 NAND2_X1 _2682_ (.A1(_1825_),
    .A2(_1655_),
    .ZN(_1826_));
 OAI22_X2 _2683_ (.A1(_1815_),
    .A2(_1821_),
    .B1(_1824_),
    .B2(_1826_),
    .ZN(_1827_));
 MUX2_X1 _2684_ (.A(_0008_),
    .B(_0010_),
    .S(_1566_),
    .Z(_1828_));
 MUX2_X1 _2685_ (.A(_1828_),
    .B(_1733_),
    .S(_1560_),
    .Z(_1829_));
 OR2_X1 _2686_ (.A1(_2136_),
    .A2(_1829_),
    .ZN(_1830_));
 MUX2_X1 _2687_ (.A(_1663_),
    .B(_1731_),
    .S(_1560_),
    .Z(_1831_));
 OAI21_X1 _2688_ (.A(_1830_),
    .B1(_1831_),
    .B2(_1583_),
    .ZN(_1832_));
 AOI22_X2 _2689_ (.A1(_1814_),
    .A2(_1827_),
    .B1(_1832_),
    .B2(_1670_),
    .ZN(_1833_));
 OAI22_X2 _2690_ (.A1(_0010_),
    .A2(_1619_),
    .B1(_1833_),
    .B2(_1673_),
    .ZN(_1834_));
 AOI221_X2 _2691_ (.A(_1587_),
    .B1(_1679_),
    .B2(\add_result[13] ),
    .C1(_1681_),
    .C2(_1834_),
    .ZN(_1835_));
 INV_X1 _2692_ (.A(\final_mant[10] ),
    .ZN(_1836_));
 BUF_X4 _2693_ (.A(_1586_),
    .Z(_1837_));
 AOI21_X1 _2694_ (.A(_1835_),
    .B1(_1836_),
    .B2(_1837_),
    .ZN(_0175_));
 BUF_X1 _2695_ (.A(_0011_),
    .Z(_1838_));
 OR2_X1 _2696_ (.A1(_1552_),
    .A2(_1838_),
    .ZN(_1839_));
 MUX2_X1 _2697_ (.A(_0009_),
    .B(_1838_),
    .S(_1567_),
    .Z(_1840_));
 MUX2_X1 _2698_ (.A(_1840_),
    .B(_1828_),
    .S(_1561_),
    .Z(_1841_));
 MUX2_X1 _2699_ (.A(_1664_),
    .B(_1841_),
    .S(_1583_),
    .Z(_1842_));
 NAND2_X1 _2700_ (.A1(_1670_),
    .A2(_1842_),
    .ZN(_1843_));
 NOR2_X2 _2701_ (.A1(_1683_),
    .A2(_1658_),
    .ZN(_1844_));
 NOR2_X1 _2702_ (.A1(_1640_),
    .A2(_1638_),
    .ZN(_1845_));
 NAND3_X1 _2703_ (.A1(_1682_),
    .A2(_1844_),
    .A3(_1845_),
    .ZN(_1846_));
 NAND2_X1 _2704_ (.A1(_1627_),
    .A2(_1640_),
    .ZN(_1847_));
 MUX2_X1 _2705_ (.A(_0010_),
    .B(_1838_),
    .S(_1622_),
    .Z(_1848_));
 MUX2_X1 _2706_ (.A(_1725_),
    .B(_1848_),
    .S(_1688_),
    .Z(_1849_));
 NAND2_X1 _2707_ (.A1(_1630_),
    .A2(_1849_),
    .ZN(_1850_));
 NAND3_X1 _2708_ (.A1(_1682_),
    .A2(_1847_),
    .A3(_1850_),
    .ZN(_1851_));
 INV_X1 _2709_ (.A(_1659_),
    .ZN(_1852_));
 OR3_X2 _2710_ (.A1(_1599_),
    .A2(_1628_),
    .A3(_1600_),
    .ZN(_1853_));
 OAI221_X1 _2711_ (.A(_1846_),
    .B1(_1851_),
    .B2(_1852_),
    .C1(_1853_),
    .C2(_1838_),
    .ZN(_1854_));
 OAI21_X1 _2712_ (.A(_1843_),
    .B1(_1854_),
    .B2(_1670_),
    .ZN(_1855_));
 OAI21_X1 _2713_ (.A(_1839_),
    .B1(_1855_),
    .B2(_1673_),
    .ZN(_1856_));
 AOI221_X2 _2714_ (.A(_1587_),
    .B1(_1679_),
    .B2(\add_result[14] ),
    .C1(_1681_),
    .C2(_1856_),
    .ZN(_1857_));
 INV_X1 _2715_ (.A(\final_mant[11] ),
    .ZN(_1858_));
 AOI21_X1 _2716_ (.A(_1857_),
    .B1(_1858_),
    .B2(_1837_),
    .ZN(_0176_));
 NAND2_X1 _2717_ (.A1(_1679_),
    .A2(\add_result[15] ),
    .ZN(_1859_));
 NOR2_X1 _2718_ (.A1(_0012_),
    .A2(_1619_),
    .ZN(_1860_));
 MUX2_X1 _2719_ (.A(_1838_),
    .B(_0012_),
    .S(_1620_),
    .Z(_1861_));
 MUX2_X1 _2720_ (.A(_1816_),
    .B(_1861_),
    .S(_1688_),
    .Z(_1862_));
 MUX2_X1 _2721_ (.A(_1693_),
    .B(_1862_),
    .S(_1630_),
    .Z(_1863_));
 NOR3_X1 _2722_ (.A1(_1804_),
    .A2(_1815_),
    .A3(_1863_),
    .ZN(_1864_));
 NOR2_X1 _2723_ (.A1(_1825_),
    .A2(_1696_),
    .ZN(_1865_));
 NOR2_X1 _2724_ (.A1(_1698_),
    .A2(_1689_),
    .ZN(_1866_));
 NOR3_X2 _2725_ (.A1(_1804_),
    .A2(_1865_),
    .A3(_1866_),
    .ZN(_1867_));
 AOI21_X1 _2726_ (.A(_1864_),
    .B1(_1867_),
    .B2(_1815_),
    .ZN(_1868_));
 MUX2_X1 _2727_ (.A(_0010_),
    .B(_0012_),
    .S(_1567_),
    .Z(_1869_));
 MUX2_X1 _2728_ (.A(_1869_),
    .B(_1840_),
    .S(_1561_),
    .Z(_1870_));
 MUX2_X1 _2729_ (.A(_1706_),
    .B(_1870_),
    .S(_1583_),
    .Z(_1871_));
 OAI22_X1 _2730_ (.A1(_1702_),
    .A2(_1868_),
    .B1(_1871_),
    .B2(_1708_),
    .ZN(_1872_));
 AOI21_X1 _2731_ (.A(_1860_),
    .B1(_1872_),
    .B2(_1737_),
    .ZN(_1873_));
 OAI21_X1 _2732_ (.A(_1859_),
    .B1(_1873_),
    .B2(_1597_),
    .ZN(_1874_));
 MUX2_X1 _2733_ (.A(\final_mant[12] ),
    .B(_1874_),
    .S(_1741_),
    .Z(_0177_));
 NAND2_X1 _2734_ (.A1(_1679_),
    .A2(\add_result[16] ),
    .ZN(_1875_));
 CLKBUF_X2 _2735_ (.A(_0013_),
    .Z(_1876_));
 NAND2_X1 _2736_ (.A1(_1674_),
    .A2(_1876_),
    .ZN(_1877_));
 OAI21_X1 _2737_ (.A(_1617_),
    .B1(_1853_),
    .B2(_1876_),
    .ZN(_1878_));
 OR2_X1 _2738_ (.A1(_1640_),
    .A2(_1728_),
    .ZN(_1879_));
 OAI22_X4 _2739_ (.A1(_1630_),
    .A2(_1723_),
    .B1(_1879_),
    .B2(_1804_),
    .ZN(_1880_));
 AND2_X1 _2740_ (.A1(_1639_),
    .A2(_1726_),
    .ZN(_1881_));
 MUX2_X1 _2741_ (.A(_0012_),
    .B(_1876_),
    .S(_1686_),
    .Z(_1882_));
 MUX2_X1 _2742_ (.A(_1848_),
    .B(_1882_),
    .S(_1624_),
    .Z(_1883_));
 AOI221_X2 _2743_ (.A(_1881_),
    .B1(_1883_),
    .B2(_1629_),
    .C1(_1651_),
    .C2(_1653_),
    .ZN(_1884_));
 AOI221_X2 _2744_ (.A(_1878_),
    .B1(_1880_),
    .B2(_1844_),
    .C1(_1884_),
    .C2(_1659_),
    .ZN(_1885_));
 MUX2_X1 _2745_ (.A(_1838_),
    .B(_1876_),
    .S(_2132_),
    .Z(_1886_));
 MUX2_X1 _2746_ (.A(_1886_),
    .B(_1869_),
    .S(_2125_),
    .Z(_1887_));
 MUX2_X1 _2747_ (.A(_1734_),
    .B(_1887_),
    .S(_1583_),
    .Z(_1888_));
 AOI21_X1 _2748_ (.A(_1885_),
    .B1(_1888_),
    .B2(_1671_),
    .ZN(_1889_));
 OAI21_X1 _2749_ (.A(_1877_),
    .B1(_1889_),
    .B2(_1674_),
    .ZN(_1890_));
 OAI21_X1 _2750_ (.A(_1875_),
    .B1(_1890_),
    .B2(_1597_),
    .ZN(_1891_));
 MUX2_X1 _2751_ (.A(\final_mant[13] ),
    .B(_1891_),
    .S(_1741_),
    .Z(_0178_));
 NAND2_X1 _2752_ (.A1(_1679_),
    .A2(\add_result[17] ),
    .ZN(_1892_));
 CLKBUF_X2 _2753_ (.A(_0014_),
    .Z(_1893_));
 NAND2_X1 _2754_ (.A1(_1674_),
    .A2(_1893_),
    .ZN(_1894_));
 OAI21_X1 _2755_ (.A(_1617_),
    .B1(_1853_),
    .B2(_1893_),
    .ZN(_1895_));
 OR2_X1 _2756_ (.A1(_1639_),
    .A2(_1819_),
    .ZN(_1896_));
 OAI22_X4 _2757_ (.A1(_1630_),
    .A2(_1824_),
    .B1(_1896_),
    .B2(_1804_),
    .ZN(_1897_));
 MUX2_X1 _2758_ (.A(_1876_),
    .B(_1893_),
    .S(_1622_),
    .Z(_1898_));
 MUX2_X1 _2759_ (.A(_1861_),
    .B(_1898_),
    .S(_1624_),
    .Z(_1899_));
 AND2_X1 _2760_ (.A1(_1629_),
    .A2(_1899_),
    .ZN(_1900_));
 AOI221_X2 _2761_ (.A(_1900_),
    .B1(_1817_),
    .B2(_1640_),
    .C1(_1651_),
    .C2(_1653_),
    .ZN(_1901_));
 AOI221_X2 _2762_ (.A(_1895_),
    .B1(_1897_),
    .B2(_1844_),
    .C1(_1901_),
    .C2(_1659_),
    .ZN(_1902_));
 MUX2_X1 _2763_ (.A(_0012_),
    .B(_1893_),
    .S(_1567_),
    .Z(_0194_));
 MUX2_X1 _2764_ (.A(_0194_),
    .B(_1886_),
    .S(_2125_),
    .Z(_0195_));
 MUX2_X1 _2765_ (.A(_1829_),
    .B(_0195_),
    .S(_1583_),
    .Z(_0196_));
 AOI21_X1 _2766_ (.A(_1902_),
    .B1(_0196_),
    .B2(_1671_),
    .ZN(_0197_));
 OAI21_X1 _2767_ (.A(_1894_),
    .B1(_0197_),
    .B2(_1674_),
    .ZN(_0198_));
 OAI21_X1 _2768_ (.A(_1892_),
    .B1(_0198_),
    .B2(_1597_),
    .ZN(_0199_));
 MUX2_X1 _2769_ (.A(\final_mant[14] ),
    .B(_0199_),
    .S(_1741_),
    .Z(_0179_));
 NAND2_X1 _2770_ (.A1(_1679_),
    .A2(\add_result[18] ),
    .ZN(_0200_));
 NOR2_X1 _2771_ (.A1(_0015_),
    .A2(_1619_),
    .ZN(_0201_));
 MUX2_X1 _2772_ (.A(_1893_),
    .B(_0015_),
    .S(_1686_),
    .Z(_0202_));
 MUX2_X1 _2773_ (.A(_1882_),
    .B(_0202_),
    .S(_1624_),
    .Z(_0203_));
 MUX2_X1 _2774_ (.A(_1849_),
    .B(_0203_),
    .S(_1630_),
    .Z(_0204_));
 NOR3_X1 _2775_ (.A1(_1804_),
    .A2(_1815_),
    .A3(_0204_),
    .ZN(_0205_));
 AOI21_X1 _2776_ (.A(_0205_),
    .B1(_1815_),
    .B2(_1654_),
    .ZN(_0206_));
 MUX2_X1 _2777_ (.A(_1876_),
    .B(_0015_),
    .S(_1567_),
    .Z(_0207_));
 MUX2_X1 _2778_ (.A(_0207_),
    .B(_0194_),
    .S(_1561_),
    .Z(_0208_));
 MUX2_X1 _2779_ (.A(_1841_),
    .B(_0208_),
    .S(_1583_),
    .Z(_0209_));
 OAI22_X1 _2780_ (.A1(_1702_),
    .A2(_0206_),
    .B1(_0209_),
    .B2(_1708_),
    .ZN(_0210_));
 AOI21_X1 _2781_ (.A(_0201_),
    .B1(_0210_),
    .B2(_1737_),
    .ZN(_0211_));
 OAI21_X1 _2782_ (.A(_0200_),
    .B1(_0211_),
    .B2(_1597_),
    .ZN(_0212_));
 MUX2_X1 _2783_ (.A(\final_mant[15] ),
    .B(_0212_),
    .S(_1741_),
    .Z(_0180_));
 AOI22_X1 _2784_ (.A1(_1751_),
    .A2(\final_mant[16] ),
    .B1(_1677_),
    .B2(\add_result[19] ),
    .ZN(_0213_));
 NAND2_X1 _2785_ (.A1(_1657_),
    .A2(_1802_),
    .ZN(_0214_));
 XNOR2_X2 _2786_ (.A(_1742_),
    .B(_1601_),
    .ZN(_0215_));
 NOR3_X1 _2787_ (.A1(_1825_),
    .A2(_0215_),
    .A3(_1862_),
    .ZN(_0216_));
 AND3_X1 _2788_ (.A1(_1825_),
    .A2(_0215_),
    .A3(_1696_),
    .ZN(_0217_));
 OAI21_X1 _2789_ (.A(_1682_),
    .B1(_0216_),
    .B2(_0217_),
    .ZN(_0218_));
 CLKBUF_X3 _2790_ (.A(_1656_),
    .Z(_0219_));
 CLKBUF_X2 _2791_ (.A(_0016_),
    .Z(_0220_));
 MUX2_X1 _2792_ (.A(_0015_),
    .B(_0220_),
    .S(_1686_),
    .Z(_0221_));
 MUX2_X1 _2793_ (.A(_1898_),
    .B(_0221_),
    .S(_1688_),
    .Z(_0222_));
 AOI21_X2 _2794_ (.A(_0222_),
    .B1(_1653_),
    .B2(_1651_),
    .ZN(_0223_));
 NAND3_X1 _2795_ (.A1(_1825_),
    .A2(_0219_),
    .A3(_0223_),
    .ZN(_0224_));
 AOI21_X1 _2796_ (.A(_1815_),
    .B1(_0218_),
    .B2(_0224_),
    .ZN(_0225_));
 NAND2_X1 _2797_ (.A1(_1682_),
    .A2(_0219_),
    .ZN(_0226_));
 NOR2_X1 _2798_ (.A1(_1698_),
    .A2(_1693_),
    .ZN(_0227_));
 AOI21_X1 _2799_ (.A(_0227_),
    .B1(_1689_),
    .B2(_1698_),
    .ZN(_0228_));
 NOR2_X1 _2800_ (.A1(_0226_),
    .A2(_0228_),
    .ZN(_0229_));
 AOI21_X1 _2801_ (.A(_0225_),
    .B1(_0229_),
    .B2(_1815_),
    .ZN(_0230_));
 OAI221_X1 _2802_ (.A(_1708_),
    .B1(_0214_),
    .B2(_0230_),
    .C1(_1853_),
    .C2(_0220_),
    .ZN(_0231_));
 MUX2_X1 _2803_ (.A(_1893_),
    .B(_0220_),
    .S(_2132_),
    .Z(_0232_));
 MUX2_X1 _2804_ (.A(_0232_),
    .B(_0207_),
    .S(_2125_),
    .Z(_0233_));
 MUX2_X1 _2805_ (.A(_1870_),
    .B(_0233_),
    .S(_2139_),
    .Z(_0234_));
 NAND2_X1 _2806_ (.A1(_1671_),
    .A2(_0234_),
    .ZN(_0235_));
 AOI21_X1 _2807_ (.A(_1746_),
    .B1(_0231_),
    .B2(_0235_),
    .ZN(_0236_));
 NAND2_X2 _2808_ (.A1(_1740_),
    .A2(_1681_),
    .ZN(_0237_));
 AOI21_X1 _2809_ (.A(_0237_),
    .B1(_0220_),
    .B2(_1746_),
    .ZN(_0238_));
 INV_X1 _2810_ (.A(_0238_),
    .ZN(_0239_));
 OAI21_X1 _2811_ (.A(_0213_),
    .B1(_0236_),
    .B2(_0239_),
    .ZN(_0181_));
 CLKBUF_X2 _2812_ (.A(_0017_),
    .Z(_0240_));
 MUX2_X1 _2813_ (.A(_0015_),
    .B(_0240_),
    .S(_2132_),
    .Z(_0241_));
 MUX2_X1 _2814_ (.A(_0241_),
    .B(_0232_),
    .S(_2125_),
    .Z(_0242_));
 MUX2_X1 _2815_ (.A(_1887_),
    .B(_0242_),
    .S(_2139_),
    .Z(_0243_));
 NAND2_X1 _2816_ (.A1(_1671_),
    .A2(_0243_),
    .ZN(_0244_));
 AND2_X1 _2817_ (.A1(_1698_),
    .A2(_1883_),
    .ZN(_0245_));
 MUX2_X1 _2818_ (.A(_0220_),
    .B(_0240_),
    .S(_1622_),
    .Z(_0246_));
 MUX2_X1 _2819_ (.A(_0202_),
    .B(_0246_),
    .S(_1688_),
    .Z(_0247_));
 AND2_X1 _2820_ (.A1(_1825_),
    .A2(_0247_),
    .ZN(_0248_));
 OAI33_X1 _2821_ (.A1(_1698_),
    .A2(_0219_),
    .A3(_1723_),
    .B1(_0226_),
    .B2(_0245_),
    .B3(_0248_),
    .ZN(_0249_));
 NOR2_X2 _2822_ (.A1(_1683_),
    .A2(_0215_),
    .ZN(_0250_));
 AOI22_X2 _2823_ (.A1(_1683_),
    .A2(_0249_),
    .B1(_0250_),
    .B2(_1729_),
    .ZN(_0251_));
 OAI221_X2 _2824_ (.A(_1708_),
    .B1(_0214_),
    .B2(_0251_),
    .C1(_1853_),
    .C2(_0240_),
    .ZN(_0252_));
 NAND4_X1 _2825_ (.A1(_1737_),
    .A2(_1598_),
    .A3(_0244_),
    .A4(_0252_),
    .ZN(_0253_));
 NOR3_X1 _2826_ (.A1(_1737_),
    .A2(_0240_),
    .A3(_0237_),
    .ZN(_0254_));
 AOI221_X1 _2827_ (.A(_0254_),
    .B1(_1676_),
    .B2(\add_result[20] ),
    .C1(_1586_),
    .C2(\final_mant[17] ),
    .ZN(_0255_));
 NAND2_X1 _2828_ (.A1(_0253_),
    .A2(_0255_),
    .ZN(_0182_));
 AOI22_X1 _2829_ (.A1(_1751_),
    .A2(\final_mant[18] ),
    .B1(_1677_),
    .B2(\add_result[21] ),
    .ZN(_0256_));
 BUF_X1 _2830_ (.A(_0018_),
    .Z(_0257_));
 NOR2_X1 _2831_ (.A1(_0257_),
    .A2(_1619_),
    .ZN(_0258_));
 OR3_X1 _2832_ (.A1(_1804_),
    .A2(_1825_),
    .A3(_1899_),
    .ZN(_0259_));
 AOI21_X1 _2833_ (.A(_0215_),
    .B1(_0259_),
    .B2(_1683_),
    .ZN(_0260_));
 MUX2_X1 _2834_ (.A(_0240_),
    .B(_0257_),
    .S(_1686_),
    .Z(_0261_));
 NOR2_X1 _2835_ (.A1(_1626_),
    .A2(_0261_),
    .ZN(_0262_));
 NOR2_X1 _2836_ (.A1(_1688_),
    .A2(_0221_),
    .ZN(_0263_));
 OAI22_X1 _2837_ (.A1(_1722_),
    .A2(_1718_),
    .B1(_0262_),
    .B2(_0263_),
    .ZN(_0264_));
 MUX2_X1 _2838_ (.A(_1824_),
    .B(_0264_),
    .S(_0219_),
    .Z(_0265_));
 NOR2_X1 _2839_ (.A1(_1698_),
    .A2(_0265_),
    .ZN(_0266_));
 NOR3_X1 _2840_ (.A1(_1605_),
    .A2(_1601_),
    .A3(_1821_),
    .ZN(_0267_));
 OAI221_X2 _2841_ (.A(_1814_),
    .B1(_0260_),
    .B2(_0266_),
    .C1(_0267_),
    .C2(_1683_),
    .ZN(_0268_));
 MUX2_X1 _2842_ (.A(_0220_),
    .B(_0257_),
    .S(_1567_),
    .Z(_0269_));
 MUX2_X1 _2843_ (.A(_0269_),
    .B(_0241_),
    .S(_2125_),
    .Z(_0270_));
 MUX2_X1 _2844_ (.A(_0195_),
    .B(_0270_),
    .S(_2139_),
    .Z(_0271_));
 OAI21_X1 _2845_ (.A(_0268_),
    .B1(_0271_),
    .B2(_1708_),
    .ZN(_0272_));
 AOI21_X1 _2846_ (.A(_0258_),
    .B1(_0272_),
    .B2(_1737_),
    .ZN(_0273_));
 OAI21_X1 _2847_ (.A(_0256_),
    .B1(_0273_),
    .B2(_0237_),
    .ZN(_0183_));
 CLKBUF_X2 _2848_ (.A(_0019_),
    .Z(_0274_));
 MUX2_X1 _2849_ (.A(_0240_),
    .B(_0274_),
    .S(_1567_),
    .Z(_0275_));
 MUX2_X1 _2850_ (.A(_0275_),
    .B(_0269_),
    .S(_1561_),
    .Z(_0276_));
 OR2_X1 _2851_ (.A1(_2136_),
    .A2(_0276_),
    .ZN(_0277_));
 OAI21_X1 _2852_ (.A(_0277_),
    .B1(_0208_),
    .B2(_1583_),
    .ZN(_0278_));
 NAND2_X1 _2853_ (.A1(_1655_),
    .A2(_0219_),
    .ZN(_0279_));
 MUX2_X1 _2854_ (.A(_0257_),
    .B(_0274_),
    .S(_1622_),
    .Z(_0280_));
 MUX2_X1 _2855_ (.A(_0246_),
    .B(_0280_),
    .S(_1624_),
    .Z(_0281_));
 MUX2_X1 _2856_ (.A(_1638_),
    .B(_0281_),
    .S(_1656_),
    .Z(_0282_));
 NOR2_X1 _2857_ (.A1(_1640_),
    .A2(_0282_),
    .ZN(_0283_));
 NOR3_X1 _2858_ (.A1(_1630_),
    .A2(_0215_),
    .A3(_0203_),
    .ZN(_0284_));
 OAI21_X1 _2859_ (.A(_1682_),
    .B1(_0283_),
    .B2(_0284_),
    .ZN(_0285_));
 OAI22_X2 _2860_ (.A1(_1851_),
    .A2(_0279_),
    .B1(_0285_),
    .B2(_1655_),
    .ZN(_0286_));
 AOI22_X2 _2861_ (.A1(_1670_),
    .A2(_0278_),
    .B1(_0286_),
    .B2(_1814_),
    .ZN(_0287_));
 OAI22_X2 _2862_ (.A1(_0274_),
    .A2(_1619_),
    .B1(_0287_),
    .B2(_1673_),
    .ZN(_0288_));
 AOI221_X2 _2863_ (.A(_1587_),
    .B1(_1588_),
    .B2(\add_result[22] ),
    .C1(_1681_),
    .C2(_0288_),
    .ZN(_0289_));
 INV_X1 _2864_ (.A(\final_mant[19] ),
    .ZN(_0290_));
 AOI21_X1 _2865_ (.A(_0289_),
    .B1(_0290_),
    .B2(_1837_),
    .ZN(_0184_));
 OAI22_X2 _2866_ (.A1(_1636_),
    .A2(_1802_),
    .B1(_1723_),
    .B2(_1805_),
    .ZN(_0291_));
 MUX2_X1 _2867_ (.A(_1636_),
    .B(_1635_),
    .S(_1560_),
    .Z(_0292_));
 NOR2_X1 _2868_ (.A1(_2004_),
    .A2(_0292_),
    .ZN(_0293_));
 NOR2_X1 _2869_ (.A1(_1570_),
    .A2(_1617_),
    .ZN(_0294_));
 AOI221_X2 _2870_ (.A(_1673_),
    .B1(_1617_),
    .B2(_0291_),
    .C1(_0293_),
    .C2(_0294_),
    .ZN(_0295_));
 AOI21_X1 _2871_ (.A(_0295_),
    .B1(_1636_),
    .B2(_1674_),
    .ZN(_0296_));
 AOI221_X2 _2872_ (.A(_1587_),
    .B1(_1588_),
    .B2(\add_result[4] ),
    .C1(_1681_),
    .C2(_0296_),
    .ZN(_0297_));
 INV_X1 _2873_ (.A(\final_mant[1] ),
    .ZN(_0298_));
 AOI21_X1 _2874_ (.A(_0297_),
    .B1(_0298_),
    .B2(_1837_),
    .ZN(_0185_));
 AOI22_X1 _2875_ (.A1(_1751_),
    .A2(\final_mant[20] ),
    .B1(_1677_),
    .B2(\add_result[23] ),
    .ZN(_0299_));
 NAND2_X1 _2876_ (.A1(_1737_),
    .A2(_1671_),
    .ZN(_0300_));
 MUX2_X1 _2877_ (.A(_0257_),
    .B(_1555_),
    .S(_2132_),
    .Z(_0301_));
 MUX2_X1 _2878_ (.A(_0301_),
    .B(_0275_),
    .S(_2125_),
    .Z(_0302_));
 MUX2_X1 _2879_ (.A(_0233_),
    .B(_0302_),
    .S(_2139_),
    .Z(_0303_));
 OAI22_X1 _2880_ (.A1(_1555_),
    .A2(_1619_),
    .B1(_0300_),
    .B2(_0303_),
    .ZN(_0304_));
 NOR2_X1 _2881_ (.A1(_1746_),
    .A2(_1702_),
    .ZN(_0305_));
 NOR2_X1 _2882_ (.A1(_0219_),
    .A2(_1867_),
    .ZN(_0306_));
 MUX2_X1 _2883_ (.A(_0274_),
    .B(_1555_),
    .S(_1686_),
    .Z(_0307_));
 MUX2_X1 _2884_ (.A(_0261_),
    .B(_0307_),
    .S(_1688_),
    .Z(_0308_));
 NOR2_X1 _2885_ (.A1(_1698_),
    .A2(_0308_),
    .ZN(_0309_));
 AOI221_X2 _2886_ (.A(_0215_),
    .B1(_0223_),
    .B2(_1698_),
    .C1(_0309_),
    .C2(_1682_),
    .ZN(_0310_));
 OAI33_X1 _2887_ (.A1(_1804_),
    .A2(_1863_),
    .A3(_0279_),
    .B1(_0306_),
    .B2(_0310_),
    .B3(_1815_),
    .ZN(_0311_));
 AOI21_X1 _2888_ (.A(_0304_),
    .B1(_0305_),
    .B2(_0311_),
    .ZN(_0312_));
 OAI21_X1 _2889_ (.A(_0299_),
    .B1(_0312_),
    .B2(_0237_),
    .ZN(_0186_));
 AOI22_X1 _2890_ (.A1(_1751_),
    .A2(\final_mant[21] ),
    .B1(_1677_),
    .B2(\add_result[24] ),
    .ZN(_0313_));
 NOR2_X1 _2891_ (.A1(_2139_),
    .A2(_0242_),
    .ZN(_0314_));
 OAI21_X1 _2892_ (.A(_1562_),
    .B1(_0021_),
    .B2(_1553_),
    .ZN(_0315_));
 OAI21_X1 _2893_ (.A(_0315_),
    .B1(_1553_),
    .B2(_1555_),
    .ZN(_0316_));
 NAND2_X1 _2894_ (.A1(_2132_),
    .A2(_0316_),
    .ZN(_0317_));
 MUX2_X1 _2895_ (.A(_0274_),
    .B(_0257_),
    .S(_2125_),
    .Z(_0318_));
 OAI21_X1 _2896_ (.A(_0317_),
    .B1(_0318_),
    .B2(_2132_),
    .ZN(_0319_));
 AOI21_X1 _2897_ (.A(_0314_),
    .B1(_0319_),
    .B2(_2139_),
    .ZN(_0320_));
 OAI22_X1 _2898_ (.A1(_1558_),
    .A2(_1619_),
    .B1(_0300_),
    .B2(_0320_),
    .ZN(_0321_));
 NAND2_X1 _2899_ (.A1(_1884_),
    .A2(_0250_),
    .ZN(_0322_));
 MUX2_X1 _2900_ (.A(_1555_),
    .B(_1558_),
    .S(_1686_),
    .Z(_0323_));
 MUX2_X1 _2901_ (.A(_0280_),
    .B(_0323_),
    .S(_1688_),
    .Z(_0324_));
 MUX2_X1 _2902_ (.A(_0247_),
    .B(_0324_),
    .S(_1825_),
    .Z(_0325_));
 OAI21_X1 _2903_ (.A(_0219_),
    .B1(_0325_),
    .B2(_1804_),
    .ZN(_0326_));
 OAI21_X1 _2904_ (.A(_0326_),
    .B1(_1880_),
    .B2(_0219_),
    .ZN(_0327_));
 OAI21_X1 _2905_ (.A(_0322_),
    .B1(_0327_),
    .B2(_1815_),
    .ZN(_0328_));
 AOI21_X1 _2906_ (.A(_0321_),
    .B1(_0328_),
    .B2(_0305_),
    .ZN(_0329_));
 OAI21_X1 _2907_ (.A(_0313_),
    .B1(_0329_),
    .B2(_0237_),
    .ZN(_0187_));
 NAND2_X1 _2908_ (.A1(_1751_),
    .A2(\final_mant[22] ),
    .ZN(_0330_));
 AOI221_X2 _2909_ (.A(_1670_),
    .B1(_1901_),
    .B2(_0250_),
    .C1(_1601_),
    .C2(_1554_),
    .ZN(_0331_));
 NOR2_X1 _2910_ (.A1(_1688_),
    .A2(_0307_),
    .ZN(_0332_));
 MUX2_X1 _2911_ (.A(_1558_),
    .B(_0021_),
    .S(_1686_),
    .Z(_0333_));
 NOR2_X1 _2912_ (.A1(_1626_),
    .A2(_0333_),
    .ZN(_0334_));
 OAI21_X1 _2913_ (.A(_1825_),
    .B1(_0332_),
    .B2(_0334_),
    .ZN(_0335_));
 OAI221_X1 _2914_ (.A(_0219_),
    .B1(_0264_),
    .B2(_1825_),
    .C1(_0335_),
    .C2(_1804_),
    .ZN(_0336_));
 OAI21_X1 _2915_ (.A(_0336_),
    .B1(_1897_),
    .B2(_0219_),
    .ZN(_0337_));
 OAI21_X1 _2916_ (.A(_0331_),
    .B1(_0337_),
    .B2(_1815_),
    .ZN(_0338_));
 NAND2_X1 _2917_ (.A1(_2136_),
    .A2(_0270_),
    .ZN(_0339_));
 MUX2_X1 _2918_ (.A(_1555_),
    .B(_0274_),
    .S(_1561_),
    .Z(_0340_));
 OAI21_X1 _2919_ (.A(_1554_),
    .B1(_1553_),
    .B2(_1562_),
    .ZN(_0341_));
 MUX2_X1 _2920_ (.A(_0340_),
    .B(_0341_),
    .S(_2132_),
    .Z(_0342_));
 NAND2_X1 _2921_ (.A1(_2139_),
    .A2(_0342_),
    .ZN(_0343_));
 AOI21_X1 _2922_ (.A(_1708_),
    .B1(_0339_),
    .B2(_0343_),
    .ZN(_0344_));
 NOR3_X1 _2923_ (.A1(_1746_),
    .A2(_1597_),
    .A3(_0344_),
    .ZN(_0345_));
 OAI21_X1 _2924_ (.A(_1589_),
    .B1(_0021_),
    .B2(_1680_),
    .ZN(_0346_));
 AOI22_X1 _2925_ (.A1(_0338_),
    .A2(_0345_),
    .B1(_0346_),
    .B2(_1746_),
    .ZN(_0347_));
 OAI21_X1 _2926_ (.A(_0330_),
    .B1(_0347_),
    .B2(_1813_),
    .ZN(_0188_));
 OAI221_X1 _2927_ (.A(_1617_),
    .B1(_1805_),
    .B2(_1824_),
    .C1(_1802_),
    .C2(_1632_),
    .ZN(_0348_));
 NOR2_X1 _2928_ (.A1(_1561_),
    .A2(_1667_),
    .ZN(_0349_));
 NOR2_X1 _2929_ (.A1(_1636_),
    .A2(_2004_),
    .ZN(_0350_));
 AOI21_X1 _2930_ (.A(_0349_),
    .B1(_0350_),
    .B2(_2125_),
    .ZN(_0351_));
 OAI21_X1 _2931_ (.A(_1670_),
    .B1(_0351_),
    .B2(_2136_),
    .ZN(_0352_));
 AOI21_X1 _2932_ (.A(_1673_),
    .B1(_0348_),
    .B2(_0352_),
    .ZN(_0353_));
 AOI21_X1 _2933_ (.A(_0353_),
    .B1(_1632_),
    .B2(_1674_),
    .ZN(_0354_));
 AOI221_X2 _2934_ (.A(_1587_),
    .B1(_1588_),
    .B2(\add_result[5] ),
    .C1(_1681_),
    .C2(_0354_),
    .ZN(_0355_));
 INV_X1 _2935_ (.A(\final_mant[2] ),
    .ZN(_0356_));
 AOI21_X1 _2936_ (.A(_0355_),
    .B1(_0356_),
    .B2(_1837_),
    .ZN(_0189_));
 INV_X1 _2937_ (.A(_1668_),
    .ZN(_0357_));
 OR3_X1 _2938_ (.A1(_1803_),
    .A2(_1638_),
    .A3(_1805_),
    .ZN(_0358_));
 OAI21_X1 _2939_ (.A(_0358_),
    .B1(_1802_),
    .B2(_1633_),
    .ZN(_0359_));
 AOI221_X2 _2940_ (.A(_1551_),
    .B1(_0357_),
    .B2(_0294_),
    .C1(_0359_),
    .C2(_1617_),
    .ZN(_0360_));
 AOI21_X1 _2941_ (.A(_0360_),
    .B1(_1633_),
    .B2(_1674_),
    .ZN(_0361_));
 AOI221_X2 _2942_ (.A(_1587_),
    .B1(_1588_),
    .B2(\add_result[6] ),
    .C1(_1681_),
    .C2(_0361_),
    .ZN(_0362_));
 INV_X1 _2943_ (.A(\final_mant[3] ),
    .ZN(_0363_));
 AOI21_X1 _2944_ (.A(_0362_),
    .B1(_0363_),
    .B2(_1837_),
    .ZN(_0190_));
 AOI22_X1 _2945_ (.A1(_1751_),
    .A2(\final_mant[4] ),
    .B1(_1677_),
    .B2(\add_result[7] ),
    .ZN(_0364_));
 AOI21_X1 _2946_ (.A(_1671_),
    .B1(_1659_),
    .B2(_1867_),
    .ZN(_0365_));
 NOR2_X1 _2947_ (.A1(_2136_),
    .A2(_1704_),
    .ZN(_0366_));
 NOR3_X1 _2948_ (.A1(_1635_),
    .A2(_2139_),
    .A3(_1808_),
    .ZN(_0367_));
 NOR3_X1 _2949_ (.A1(_1708_),
    .A2(_0366_),
    .A3(_0367_),
    .ZN(_0368_));
 NOR3_X1 _2950_ (.A1(_1746_),
    .A2(_0365_),
    .A3(_0368_),
    .ZN(_0369_));
 OAI21_X1 _2951_ (.A(_1737_),
    .B1(_1853_),
    .B2(_0368_),
    .ZN(_0370_));
 INV_X1 _2952_ (.A(_0004_),
    .ZN(_0371_));
 AOI21_X1 _2953_ (.A(_0369_),
    .B1(_0370_),
    .B2(_0371_),
    .ZN(_0372_));
 OAI21_X1 _2954_ (.A(_0364_),
    .B1(_0372_),
    .B2(_0237_),
    .ZN(_0191_));
 INV_X1 _2955_ (.A(_1732_),
    .ZN(_0373_));
 MUX2_X1 _2956_ (.A(_0373_),
    .B(_0293_),
    .S(_2136_),
    .Z(_0374_));
 AOI22_X1 _2957_ (.A1(_1661_),
    .A2(_1880_),
    .B1(_0374_),
    .B2(_1670_),
    .ZN(_0375_));
 OAI22_X2 _2958_ (.A1(_0005_),
    .A2(_1618_),
    .B1(_0375_),
    .B2(_1673_),
    .ZN(_0376_));
 AOI221_X2 _2959_ (.A(_1587_),
    .B1(_1588_),
    .B2(\add_result[8] ),
    .C1(_1681_),
    .C2(_0376_),
    .ZN(_0377_));
 INV_X1 _2960_ (.A(\final_mant[5] ),
    .ZN(_0378_));
 AOI21_X1 _2961_ (.A(_0377_),
    .B1(_0378_),
    .B2(_1837_),
    .ZN(_0192_));
 OR2_X1 _2962_ (.A1(_2136_),
    .A2(_1831_),
    .ZN(_0379_));
 OAI21_X1 _2963_ (.A(_0379_),
    .B1(_0351_),
    .B2(_1583_),
    .ZN(_0380_));
 AOI22_X1 _2964_ (.A1(_1661_),
    .A2(_1897_),
    .B1(_0380_),
    .B2(_1670_),
    .ZN(_0381_));
 OAI22_X2 _2965_ (.A1(_0006_),
    .A2(_1618_),
    .B1(_0381_),
    .B2(_1673_),
    .ZN(_0382_));
 AOI221_X2 _2966_ (.A(_1587_),
    .B1(_1588_),
    .B2(\add_result[9] ),
    .C1(_1681_),
    .C2(_0382_),
    .ZN(_0383_));
 INV_X1 _2967_ (.A(\final_mant[6] ),
    .ZN(_0384_));
 AOI21_X1 _2968_ (.A(_0383_),
    .B1(_0384_),
    .B2(_1837_),
    .ZN(_0193_));
 NAND4_X2 _2969_ (.A1(net21),
    .A2(net20),
    .A3(net24),
    .A4(net22),
    .ZN(_0385_));
 NAND4_X2 _2970_ (.A1(net17),
    .A2(net16),
    .A3(net19),
    .A4(net18),
    .ZN(_0386_));
 NOR2_X4 _2971_ (.A1(_0385_),
    .A2(_0386_),
    .ZN(_0387_));
 NOR4_X1 _2972_ (.A1(net12),
    .A2(net1),
    .A3(net26),
    .A4(net15),
    .ZN(_0388_));
 CLKBUF_X2 _2973_ (.A(net8),
    .Z(_0389_));
 CLKBUF_X2 _2974_ (.A(net13),
    .Z(_0390_));
 NOR4_X1 _2975_ (.A1(_0389_),
    .A2(net10),
    .A3(net14),
    .A4(_0390_),
    .ZN(_0391_));
 BUF_X2 _2976_ (.A(net2),
    .Z(_0392_));
 BUF_X2 _2977_ (.A(net6),
    .Z(_0393_));
 NOR4_X1 _2978_ (.A1(_0392_),
    .A2(_0393_),
    .A3(net9),
    .A4(net11),
    .ZN(_0394_));
 CLKBUF_X2 _2979_ (.A(net5),
    .Z(_0395_));
 CLKBUF_X2 _2980_ (.A(net4),
    .Z(_0396_));
 CLKBUF_X2 _2981_ (.A(net7),
    .Z(_0397_));
 NOR3_X1 _2982_ (.A1(_0395_),
    .A2(_0396_),
    .A3(_0397_),
    .ZN(_0398_));
 NAND4_X1 _2983_ (.A1(_0388_),
    .A2(_0391_),
    .A3(_0394_),
    .A4(_0398_),
    .ZN(_0399_));
 BUF_X2 _2984_ (.A(net27),
    .Z(_0400_));
 BUF_X1 _2985_ (.A(net32),
    .Z(_0401_));
 BUF_X1 _2986_ (.A(net31),
    .Z(_0402_));
 NOR4_X1 _2987_ (.A1(_0400_),
    .A2(net29),
    .A3(_0401_),
    .A4(_0402_),
    .ZN(_0403_));
 CLKBUF_X2 _2988_ (.A(net30),
    .Z(_0404_));
 CLKBUF_X2 _2989_ (.A(net3),
    .Z(_0405_));
 NOR4_X1 _2990_ (.A1(net23),
    .A2(net28),
    .A3(_0404_),
    .A4(_0405_),
    .ZN(_0406_));
 NAND2_X1 _2991_ (.A1(_0403_),
    .A2(_0406_),
    .ZN(_0407_));
 NOR2_X1 _2992_ (.A1(_0399_),
    .A2(_0407_),
    .ZN(_0408_));
 INV_X1 _2993_ (.A(_0408_),
    .ZN(_0409_));
 BUF_X1 _2994_ (.A(is_a_larger_stage1),
    .Z(_0410_));
 CLKBUF_X3 _2995_ (.A(_0410_),
    .Z(_0411_));
 BUF_X4 _2996_ (.A(_0411_),
    .Z(_0412_));
 MUX2_X1 _2997_ (.A(b_sign_stage1),
    .B(a_sign_stage1),
    .S(_0412_),
    .Z(_0413_));
 AND2_X1 _2998_ (.A1(_0387_),
    .A2(_0408_),
    .ZN(_0414_));
 MUX2_X1 _2999_ (.A(_0413_),
    .B(net25),
    .S(_0414_),
    .Z(_0415_));
 NAND4_X2 _3000_ (.A1(net41),
    .A2(net40),
    .A3(net42),
    .A4(net43),
    .ZN(_0416_));
 NAND4_X2 _3001_ (.A1(net45),
    .A2(net44),
    .A3(net48),
    .A4(net46),
    .ZN(_0417_));
 OAI21_X1 _3002_ (.A(_0415_),
    .B1(_0416_),
    .B2(_0417_),
    .ZN(_0418_));
 NOR2_X2 _3003_ (.A1(_0417_),
    .A2(_0416_),
    .ZN(_0419_));
 MUX2_X1 _3004_ (.A(net49),
    .B(_2122_),
    .S(_0414_),
    .Z(_0420_));
 NOR4_X4 _3005_ (.A1(net38),
    .A2(net33),
    .A3(net50),
    .A4(_1582_),
    .ZN(_0421_));
 NOR4_X2 _3006_ (.A1(_1577_),
    .A2(_1579_),
    .A3(_1581_),
    .A4(net39),
    .ZN(_0422_));
 NOR4_X2 _3007_ (.A1(net34),
    .A2(_1576_),
    .A3(_1578_),
    .A4(_1580_),
    .ZN(_0423_));
 NOR3_X2 _3008_ (.A1(_1575_),
    .A2(net36),
    .A3(net37),
    .ZN(_0424_));
 NAND4_X4 _3009_ (.A1(_0421_),
    .A2(_0422_),
    .A3(_0423_),
    .A4(_0424_),
    .ZN(_0425_));
 NOR4_X1 _3010_ (.A1(net51),
    .A2(_1571_),
    .A3(_1574_),
    .A4(_1573_),
    .ZN(_0426_));
 NOR4_X2 _3011_ (.A1(net47),
    .A2(net52),
    .A3(_1572_),
    .A4(net35),
    .ZN(_0427_));
 NAND2_X2 _3012_ (.A1(_0426_),
    .A2(_0427_),
    .ZN(_0428_));
 NOR2_X1 _3013_ (.A1(_0425_),
    .A2(_0428_),
    .ZN(_0429_));
 NAND3_X1 _3014_ (.A1(_0419_),
    .A2(_0420_),
    .A3(_0429_),
    .ZN(_0430_));
 AOI221_X1 _3015_ (.A(_1586_),
    .B1(_0387_),
    .B2(_0409_),
    .C1(_0418_),
    .C2(_0430_),
    .ZN(_0082_));
 NOR3_X1 _3016_ (.A1(_1746_),
    .A2(_0237_),
    .A3(_1671_),
    .ZN(_0083_));
 NOR2_X1 _3017_ (.A1(_0419_),
    .A2(_0387_),
    .ZN(_0431_));
 NAND2_X2 _3018_ (.A1(_1740_),
    .A2(_0431_),
    .ZN(_0432_));
 CLKBUF_X3 _3019_ (.A(_0432_),
    .Z(_0433_));
 CLKBUF_X3 _3020_ (.A(_2222_),
    .Z(_0434_));
 INV_X1 _3021_ (.A(_0434_),
    .ZN(_0435_));
 INV_X1 _3022_ (.A(_2218_),
    .ZN(_0436_));
 CLKBUF_X3 _3023_ (.A(_2214_),
    .Z(_0437_));
 INV_X1 _3024_ (.A(_0437_),
    .ZN(_0438_));
 BUF_X2 _3025_ (.A(_2206_),
    .Z(_0439_));
 INV_X1 _3026_ (.A(_2202_),
    .ZN(_0440_));
 BUF_X1 _3027_ (.A(_2190_),
    .Z(_0441_));
 INV_X1 _3028_ (.A(_0441_),
    .ZN(_0442_));
 NOR2_X1 _3029_ (.A1(_0442_),
    .A2(_2194_),
    .ZN(_0443_));
 BUF_X2 _3030_ (.A(_2198_),
    .Z(_0444_));
 OAI21_X2 _3031_ (.A(_0440_),
    .B1(_0443_),
    .B2(_0444_),
    .ZN(_0445_));
 INV_X1 _3032_ (.A(_0445_),
    .ZN(_0446_));
 CLKBUF_X3 _3033_ (.A(_2166_),
    .Z(_0447_));
 CLKBUF_X3 _3034_ (.A(_2174_),
    .Z(_0448_));
 CLKBUF_X3 _3035_ (.A(_2182_),
    .Z(_0449_));
 INV_X1 _3036_ (.A(_2162_),
    .ZN(_0450_));
 BUF_X1 _3037_ (.A(\aligned_a_mant[0] ),
    .Z(_0451_));
 CLKBUF_X2 _3038_ (.A(\aligned_b_mant[0] ),
    .Z(_0452_));
 NAND2_X1 _3039_ (.A1(_0451_),
    .A2(_0452_),
    .ZN(_0453_));
 OAI21_X2 _3040_ (.A(_0450_),
    .B1(_0453_),
    .B2(_2158_),
    .ZN(_0454_));
 INV_X2 _3041_ (.A(_2150_),
    .ZN(_0455_));
 AOI21_X4 _3042_ (.A(_2154_),
    .B1(_0454_),
    .B2(_0455_),
    .ZN(_0456_));
 OR4_X1 _3043_ (.A1(_0447_),
    .A2(_0448_),
    .A3(_0449_),
    .A4(_0456_),
    .ZN(_0457_));
 INV_X1 _3044_ (.A(_2186_),
    .ZN(_0458_));
 INV_X1 _3045_ (.A(_0448_),
    .ZN(_0459_));
 AOI21_X1 _3046_ (.A(_2178_),
    .B1(_0459_),
    .B2(_2170_),
    .ZN(_0460_));
 OAI21_X1 _3047_ (.A(_0458_),
    .B1(_0460_),
    .B2(_0449_),
    .ZN(_0461_));
 NOR3_X1 _3048_ (.A1(_2194_),
    .A2(_2202_),
    .A3(_0461_),
    .ZN(_0462_));
 AOI211_X2 _3049_ (.A(_0439_),
    .B(_0446_),
    .C1(_0457_),
    .C2(_0462_),
    .ZN(_0463_));
 OAI21_X1 _3050_ (.A(_0438_),
    .B1(_0463_),
    .B2(_2210_),
    .ZN(_0464_));
 XNOR2_X2 _3051_ (.A(b_sign_stage1),
    .B(a_sign_stage1),
    .ZN(_0465_));
 AND3_X1 _3052_ (.A1(_0436_),
    .A2(_0464_),
    .A3(_0465_),
    .ZN(_0466_));
 AOI21_X1 _3053_ (.A(_2216_),
    .B1(_2208_),
    .B2(_0437_),
    .ZN(_0467_));
 AOI21_X2 _3054_ (.A(_2200_),
    .B1(_2192_),
    .B2(_0444_),
    .ZN(_0468_));
 NAND2_X1 _3055_ (.A1(_0439_),
    .A2(_0437_),
    .ZN(_0469_));
 OAI21_X1 _3056_ (.A(_0467_),
    .B1(_0468_),
    .B2(_0469_),
    .ZN(_0470_));
 AND2_X1 _3057_ (.A1(_0411_),
    .A2(_0470_),
    .ZN(_0471_));
 AOI21_X1 _3058_ (.A(_2213_),
    .B1(_2205_),
    .B2(_0437_),
    .ZN(_0472_));
 AOI21_X2 _3059_ (.A(_2197_),
    .B1(_2189_),
    .B2(_0444_),
    .ZN(_0473_));
 OAI21_X1 _3060_ (.A(_0472_),
    .B1(_0469_),
    .B2(_0473_),
    .ZN(_0474_));
 INV_X1 _3061_ (.A(_0410_),
    .ZN(_0475_));
 AOI21_X1 _3062_ (.A(_0471_),
    .B1(_0474_),
    .B2(_0475_),
    .ZN(_0476_));
 AND2_X1 _3063_ (.A1(_0441_),
    .A2(_0444_),
    .ZN(_0477_));
 AND3_X1 _3064_ (.A1(_0439_),
    .A2(_0437_),
    .A3(_0477_),
    .ZN(_0478_));
 INV_X1 _3065_ (.A(_2158_),
    .ZN(_0479_));
 INV_X1 _3066_ (.A(_0451_),
    .ZN(_0480_));
 AOI21_X1 _3067_ (.A(_0479_),
    .B1(_0452_),
    .B2(_0480_),
    .ZN(_0481_));
 NOR3_X1 _3068_ (.A1(_0475_),
    .A2(_2160_),
    .A3(_0481_),
    .ZN(_0482_));
 INV_X1 _3069_ (.A(_0452_),
    .ZN(_0483_));
 AOI21_X1 _3070_ (.A(_0479_),
    .B1(_0483_),
    .B2(_0451_),
    .ZN(_0484_));
 NOR3_X1 _3071_ (.A1(_0410_),
    .A2(_2157_),
    .A3(_0484_),
    .ZN(_0485_));
 AND2_X1 _3072_ (.A1(_2150_),
    .A2(_0447_),
    .ZN(_0486_));
 NAND3_X1 _3073_ (.A1(_0448_),
    .A2(_0449_),
    .A3(_0486_),
    .ZN(_0487_));
 NOR3_X1 _3074_ (.A1(_0482_),
    .A2(_0485_),
    .A3(_0487_),
    .ZN(_0488_));
 AOI21_X1 _3075_ (.A(_2181_),
    .B1(_2173_),
    .B2(_0449_),
    .ZN(_0489_));
 NAND2_X1 _3076_ (.A1(_0448_),
    .A2(_0449_),
    .ZN(_0490_));
 AOI21_X2 _3077_ (.A(_2165_),
    .B1(_2149_),
    .B2(_0447_),
    .ZN(_0491_));
 OAI21_X1 _3078_ (.A(_0489_),
    .B1(_0490_),
    .B2(_0491_),
    .ZN(_0492_));
 AOI21_X1 _3079_ (.A(_2184_),
    .B1(_2176_),
    .B2(_0449_),
    .ZN(_0493_));
 AOI21_X2 _3080_ (.A(_2168_),
    .B1(_2152_),
    .B2(_0447_),
    .ZN(_0494_));
 OAI21_X1 _3081_ (.A(_0493_),
    .B1(_0494_),
    .B2(_0490_),
    .ZN(_0495_));
 MUX2_X1 _3082_ (.A(_0492_),
    .B(_0495_),
    .S(_0410_),
    .Z(_0496_));
 OAI21_X1 _3083_ (.A(_0478_),
    .B1(_0488_),
    .B2(_0496_),
    .ZN(_0497_));
 NAND2_X1 _3084_ (.A1(_0476_),
    .A2(_0497_),
    .ZN(_0498_));
 XOR2_X2 _3085_ (.A(b_sign_stage1),
    .B(a_sign_stage1),
    .Z(_0499_));
 CLKBUF_X3 _3086_ (.A(_0499_),
    .Z(_0500_));
 CLKBUF_X3 _3087_ (.A(_0500_),
    .Z(_0501_));
 AOI21_X1 _3088_ (.A(_0466_),
    .B1(_0498_),
    .B2(_0501_),
    .ZN(_0502_));
 XNOR2_X1 _3089_ (.A(_0435_),
    .B(_0502_),
    .ZN(_0503_));
 NOR2_X1 _3090_ (.A1(_0433_),
    .A2(_0503_),
    .ZN(_0088_));
 INV_X1 _3091_ (.A(_2230_),
    .ZN(_0504_));
 AOI21_X1 _3092_ (.A(_2189_),
    .B1(_2181_),
    .B2(_0441_),
    .ZN(_0505_));
 AOI21_X1 _3093_ (.A(_2192_),
    .B1(_2184_),
    .B2(_0441_),
    .ZN(_0506_));
 MUX2_X1 _3094_ (.A(_0505_),
    .B(_0506_),
    .S(_0411_),
    .Z(_0507_));
 NOR2_X1 _3095_ (.A1(_0411_),
    .A2(_2173_),
    .ZN(_0508_));
 INV_X1 _3096_ (.A(_2165_),
    .ZN(_0509_));
 OAI21_X1 _3097_ (.A(_0508_),
    .B1(_0509_),
    .B2(_0459_),
    .ZN(_0510_));
 INV_X1 _3098_ (.A(_2176_),
    .ZN(_0511_));
 NAND2_X1 _3099_ (.A1(_0448_),
    .A2(_2168_),
    .ZN(_0512_));
 NAND3_X1 _3100_ (.A1(_0411_),
    .A2(_0511_),
    .A3(_0512_),
    .ZN(_0513_));
 AND2_X1 _3101_ (.A1(_0510_),
    .A2(_0513_),
    .ZN(_0514_));
 AND2_X1 _3102_ (.A1(_0447_),
    .A2(_0448_),
    .ZN(_0515_));
 INV_X1 _3103_ (.A(_2157_),
    .ZN(_0516_));
 OAI21_X2 _3104_ (.A(_2158_),
    .B1(_0452_),
    .B2(_0480_),
    .ZN(_0517_));
 AOI21_X4 _3105_ (.A(_0455_),
    .B1(_0516_),
    .B2(_0517_),
    .ZN(_0518_));
 OR2_X1 _3106_ (.A1(_2149_),
    .A2(_0510_),
    .ZN(_0519_));
 OAI22_X4 _3107_ (.A1(_0514_),
    .A2(_0515_),
    .B1(_0518_),
    .B2(_0519_),
    .ZN(_0520_));
 AND2_X1 _3108_ (.A1(_0449_),
    .A2(_0441_),
    .ZN(_0521_));
 INV_X1 _3109_ (.A(_2160_),
    .ZN(_0522_));
 OAI21_X1 _3110_ (.A(_2158_),
    .B1(_0483_),
    .B2(_0451_),
    .ZN(_0523_));
 AOI21_X2 _3111_ (.A(_0455_),
    .B1(_0522_),
    .B2(_0523_),
    .ZN(_0524_));
 OR2_X1 _3112_ (.A1(_2152_),
    .A2(_0513_),
    .ZN(_0525_));
 OAI21_X1 _3113_ (.A(_0521_),
    .B1(_0524_),
    .B2(_0525_),
    .ZN(_0526_));
 OAI21_X2 _3114_ (.A(_0507_),
    .B1(_0520_),
    .B2(_0526_),
    .ZN(_0527_));
 AND2_X1 _3115_ (.A1(_0444_),
    .A2(_0439_),
    .ZN(_0528_));
 NAND4_X2 _3116_ (.A1(_0437_),
    .A2(_0434_),
    .A3(_0527_),
    .A4(_0528_),
    .ZN(_0529_));
 INV_X1 _3117_ (.A(_2216_),
    .ZN(_0530_));
 AOI21_X1 _3118_ (.A(_2208_),
    .B1(_2200_),
    .B2(_0439_),
    .ZN(_0531_));
 OAI21_X1 _3119_ (.A(_0530_),
    .B1(_0531_),
    .B2(_0438_),
    .ZN(_0532_));
 AOI21_X1 _3120_ (.A(_2224_),
    .B1(_0532_),
    .B2(_0434_),
    .ZN(_0533_));
 INV_X1 _3121_ (.A(_2213_),
    .ZN(_0534_));
 AOI21_X1 _3122_ (.A(_2205_),
    .B1(_2197_),
    .B2(_0439_),
    .ZN(_0535_));
 OAI21_X1 _3123_ (.A(_0534_),
    .B1(_0535_),
    .B2(_0438_),
    .ZN(_0536_));
 AOI21_X1 _3124_ (.A(_2221_),
    .B1(_0536_),
    .B2(_0434_),
    .ZN(_0537_));
 CLKBUF_X3 _3125_ (.A(_0475_),
    .Z(_0538_));
 MUX2_X1 _3126_ (.A(_0533_),
    .B(_0537_),
    .S(_0538_),
    .Z(_0539_));
 AND2_X1 _3127_ (.A1(_0529_),
    .A2(_0539_),
    .ZN(_0540_));
 NAND2_X1 _3128_ (.A1(_0501_),
    .A2(_0540_),
    .ZN(_0541_));
 CLKBUF_X3 _3129_ (.A(_0465_),
    .Z(_0542_));
 AOI21_X1 _3130_ (.A(_0434_),
    .B1(_0464_),
    .B2(_0436_),
    .ZN(_0543_));
 OAI21_X1 _3131_ (.A(_0542_),
    .B1(_0543_),
    .B2(_2226_),
    .ZN(_0544_));
 NAND2_X1 _3132_ (.A1(_0541_),
    .A2(_0544_),
    .ZN(_0545_));
 XNOR2_X1 _3133_ (.A(_0504_),
    .B(_0545_),
    .ZN(_0546_));
 NOR2_X1 _3134_ (.A1(_0433_),
    .A2(_0546_),
    .ZN(_0089_));
 BUF_X4 _3135_ (.A(_2238_),
    .Z(_0547_));
 INV_X2 _3136_ (.A(_0547_),
    .ZN(_0548_));
 INV_X1 _3137_ (.A(_2232_),
    .ZN(_0549_));
 BUF_X4 _3138_ (.A(_2230_),
    .Z(_0550_));
 NOR2_X1 _3139_ (.A1(_0435_),
    .A2(_0467_),
    .ZN(_0551_));
 OAI21_X1 _3140_ (.A(_0550_),
    .B1(_2224_),
    .B2(_0551_),
    .ZN(_0552_));
 NAND3_X1 _3141_ (.A1(_0411_),
    .A2(_0549_),
    .A3(_0552_),
    .ZN(_0553_));
 NAND4_X1 _3142_ (.A1(_0439_),
    .A2(_0437_),
    .A3(_0434_),
    .A4(_0550_),
    .ZN(_0554_));
 OAI21_X1 _3143_ (.A(_0486_),
    .B1(_0481_),
    .B2(_2160_),
    .ZN(_0555_));
 AOI21_X1 _3144_ (.A(_0490_),
    .B1(_0494_),
    .B2(_0555_),
    .ZN(_0556_));
 INV_X1 _3145_ (.A(_0493_),
    .ZN(_0557_));
 OAI21_X1 _3146_ (.A(_0477_),
    .B1(_0556_),
    .B2(_0557_),
    .ZN(_0558_));
 AOI21_X1 _3147_ (.A(_0554_),
    .B1(_0558_),
    .B2(_0468_),
    .ZN(_0559_));
 OAI21_X1 _3148_ (.A(_0486_),
    .B1(_0484_),
    .B2(_2157_),
    .ZN(_0560_));
 AOI21_X1 _3149_ (.A(_0490_),
    .B1(_0491_),
    .B2(_0560_),
    .ZN(_0561_));
 INV_X1 _3150_ (.A(_0489_),
    .ZN(_0562_));
 OAI21_X1 _3151_ (.A(_0477_),
    .B1(_0561_),
    .B2(_0562_),
    .ZN(_0563_));
 AOI21_X1 _3152_ (.A(_0554_),
    .B1(_0563_),
    .B2(_0473_),
    .ZN(_0564_));
 INV_X1 _3153_ (.A(_2229_),
    .ZN(_0565_));
 NOR2_X1 _3154_ (.A1(_0435_),
    .A2(_0472_),
    .ZN(_0566_));
 OAI21_X1 _3155_ (.A(_0550_),
    .B1(_2221_),
    .B2(_0566_),
    .ZN(_0567_));
 NAND3_X1 _3156_ (.A1(_0538_),
    .A2(_0565_),
    .A3(_0567_),
    .ZN(_0568_));
 OAI22_X2 _3157_ (.A1(_0553_),
    .A2(_0559_),
    .B1(_0564_),
    .B2(_0568_),
    .ZN(_0569_));
 NOR2_X1 _3158_ (.A1(_0542_),
    .A2(_0569_),
    .ZN(_0570_));
 CLKBUF_X3 _3159_ (.A(_0500_),
    .Z(_0571_));
 NOR2_X1 _3160_ (.A1(_2234_),
    .A2(_0571_),
    .ZN(_0572_));
 OAI21_X1 _3161_ (.A(_0504_),
    .B1(_0543_),
    .B2(_2226_),
    .ZN(_0573_));
 AOI21_X1 _3162_ (.A(_0570_),
    .B1(_0572_),
    .B2(_0573_),
    .ZN(_0574_));
 XNOR2_X1 _3163_ (.A(_0548_),
    .B(_0574_),
    .ZN(_0575_));
 NOR2_X1 _3164_ (.A1(_0433_),
    .A2(_0575_),
    .ZN(_0090_));
 CLKBUF_X3 _3165_ (.A(_2246_),
    .Z(_0576_));
 INV_X1 _3166_ (.A(_0576_),
    .ZN(_0577_));
 AOI21_X1 _3167_ (.A(_2224_),
    .B1(_2216_),
    .B2(_2222_),
    .ZN(_0578_));
 OAI21_X1 _3168_ (.A(_0549_),
    .B1(_0578_),
    .B2(_0504_),
    .ZN(_0579_));
 AOI21_X1 _3169_ (.A(_2240_),
    .B1(_0579_),
    .B2(_0547_),
    .ZN(_0580_));
 AOI21_X1 _3170_ (.A(_2221_),
    .B1(_2213_),
    .B2(_0434_),
    .ZN(_0581_));
 OAI21_X1 _3171_ (.A(_0565_),
    .B1(_0581_),
    .B2(_0504_),
    .ZN(_0582_));
 AOI21_X1 _3172_ (.A(_2237_),
    .B1(_0582_),
    .B2(_0547_),
    .ZN(_0583_));
 MUX2_X1 _3173_ (.A(_0580_),
    .B(_0583_),
    .S(_0538_),
    .Z(_0584_));
 NAND4_X1 _3174_ (.A1(_0437_),
    .A2(_0434_),
    .A3(_0550_),
    .A4(_0547_),
    .ZN(_0585_));
 MUX2_X1 _3175_ (.A(_0531_),
    .B(_0535_),
    .S(_0475_),
    .Z(_0586_));
 INV_X1 _3176_ (.A(_0586_),
    .ZN(_0587_));
 NOR2_X1 _3177_ (.A1(_0528_),
    .A2(_0587_),
    .ZN(_0588_));
 OAI21_X1 _3178_ (.A(_0584_),
    .B1(_0585_),
    .B2(_0588_),
    .ZN(_0589_));
 NAND3_X1 _3179_ (.A1(_0507_),
    .A2(_0584_),
    .A3(_0586_),
    .ZN(_0590_));
 NOR2_X1 _3180_ (.A1(_0520_),
    .A2(_0526_),
    .ZN(_0591_));
 OAI21_X2 _3181_ (.A(_0589_),
    .B1(_0590_),
    .B2(_0591_),
    .ZN(_0592_));
 NOR2_X1 _3182_ (.A1(_0542_),
    .A2(_0592_),
    .ZN(_0593_));
 NOR4_X4 _3183_ (.A1(_0437_),
    .A2(_0434_),
    .A3(_0550_),
    .A4(_0547_),
    .ZN(_0594_));
 INV_X1 _3184_ (.A(_2234_),
    .ZN(_0595_));
 INV_X1 _3185_ (.A(_2210_),
    .ZN(_0596_));
 OAI21_X1 _3186_ (.A(_0436_),
    .B1(_0437_),
    .B2(_0596_),
    .ZN(_0597_));
 AOI21_X1 _3187_ (.A(_2226_),
    .B1(_0597_),
    .B2(_0435_),
    .ZN(_0598_));
 OAI21_X2 _3188_ (.A(_0595_),
    .B1(_0598_),
    .B2(_0550_),
    .ZN(_0599_));
 AOI221_X2 _3189_ (.A(_2242_),
    .B1(_0463_),
    .B2(_0594_),
    .C1(_0599_),
    .C2(_0548_),
    .ZN(_0600_));
 AOI21_X1 _3190_ (.A(_0593_),
    .B1(_0600_),
    .B2(_0542_),
    .ZN(_0601_));
 XNOR2_X1 _3191_ (.A(_0577_),
    .B(_0601_),
    .ZN(_0602_));
 NOR2_X1 _3192_ (.A1(_0433_),
    .A2(_0602_),
    .ZN(_0091_));
 CLKBUF_X3 _3193_ (.A(_2254_),
    .Z(_0603_));
 INV_X1 _3194_ (.A(_0603_),
    .ZN(_0604_));
 INV_X1 _3195_ (.A(_2250_),
    .ZN(_0605_));
 OAI21_X1 _3196_ (.A(_0605_),
    .B1(_0600_),
    .B2(_0576_),
    .ZN(_0606_));
 INV_X1 _3197_ (.A(_2245_),
    .ZN(_0607_));
 AOI21_X1 _3198_ (.A(_2229_),
    .B1(_2221_),
    .B2(_0550_),
    .ZN(_0608_));
 NOR2_X1 _3199_ (.A1(_0548_),
    .A2(_0608_),
    .ZN(_0609_));
 OAI21_X1 _3200_ (.A(_0576_),
    .B1(_2237_),
    .B2(_0609_),
    .ZN(_0610_));
 AOI21_X1 _3201_ (.A(_0411_),
    .B1(_0607_),
    .B2(_0610_),
    .ZN(_0611_));
 INV_X1 _3202_ (.A(_2248_),
    .ZN(_0612_));
 AOI21_X1 _3203_ (.A(_2232_),
    .B1(_2224_),
    .B2(_0550_),
    .ZN(_0613_));
 NOR2_X1 _3204_ (.A1(_0548_),
    .A2(_0613_),
    .ZN(_0614_));
 OAI21_X1 _3205_ (.A(_0576_),
    .B1(_2240_),
    .B2(_0614_),
    .ZN(_0615_));
 AOI21_X1 _3206_ (.A(_0538_),
    .B1(_0612_),
    .B2(_0615_),
    .ZN(_0616_));
 NAND4_X1 _3207_ (.A1(_0434_),
    .A2(_0550_),
    .A3(_0547_),
    .A4(_0576_),
    .ZN(_0617_));
 AOI21_X1 _3208_ (.A(_0617_),
    .B1(_0497_),
    .B2(_0476_),
    .ZN(_0618_));
 NOR3_X1 _3209_ (.A1(_0611_),
    .A2(_0616_),
    .A3(_0618_),
    .ZN(_0619_));
 MUX2_X1 _3210_ (.A(_0606_),
    .B(_0619_),
    .S(_0571_),
    .Z(_0620_));
 XNOR2_X1 _3211_ (.A(_0604_),
    .B(_0620_),
    .ZN(_0621_));
 NOR2_X1 _3212_ (.A1(_0433_),
    .A2(_0621_),
    .ZN(_0092_));
 CLKBUF_X3 _3213_ (.A(_2262_),
    .Z(_0622_));
 INV_X1 _3214_ (.A(_0622_),
    .ZN(_0623_));
 AOI21_X2 _3215_ (.A(_2242_),
    .B1(_0599_),
    .B2(_0548_),
    .ZN(_0624_));
 NOR2_X2 _3216_ (.A1(_2250_),
    .A2(_2258_),
    .ZN(_0625_));
 INV_X1 _3217_ (.A(_0439_),
    .ZN(_0626_));
 NAND3_X2 _3218_ (.A1(_0626_),
    .A2(_0445_),
    .A3(_0594_),
    .ZN(_0627_));
 NOR4_X4 _3219_ (.A1(_0447_),
    .A2(_0448_),
    .A3(_0449_),
    .A4(_0456_),
    .ZN(_0628_));
 OR3_X1 _3220_ (.A1(_2194_),
    .A2(_2202_),
    .A3(_0461_),
    .ZN(_0629_));
 NOR2_X2 _3221_ (.A1(_0628_),
    .A2(_0629_),
    .ZN(_0630_));
 OAI211_X4 _3222_ (.A(_0624_),
    .B(_0625_),
    .C1(_0627_),
    .C2(_0630_),
    .ZN(_0631_));
 AOI21_X1 _3223_ (.A(_0603_),
    .B1(_0605_),
    .B2(_2246_),
    .ZN(_0632_));
 NOR2_X1 _3224_ (.A1(_2258_),
    .A2(_0632_),
    .ZN(_0633_));
 NOR2_X1 _3225_ (.A1(_0500_),
    .A2(_0633_),
    .ZN(_0634_));
 NAND2_X1 _3226_ (.A1(_0631_),
    .A2(_0634_),
    .ZN(_0635_));
 AOI21_X1 _3227_ (.A(_2240_),
    .B1(_2232_),
    .B2(_0547_),
    .ZN(_0636_));
 OAI21_X1 _3228_ (.A(_0612_),
    .B1(_0636_),
    .B2(_0577_),
    .ZN(_0637_));
 AOI21_X1 _3229_ (.A(_2256_),
    .B1(_0637_),
    .B2(_0603_),
    .ZN(_0638_));
 AOI21_X1 _3230_ (.A(_2237_),
    .B1(_2229_),
    .B2(_0547_),
    .ZN(_0639_));
 OAI21_X1 _3231_ (.A(_0607_),
    .B1(_0639_),
    .B2(_0577_),
    .ZN(_0640_));
 AOI21_X1 _3232_ (.A(_2253_),
    .B1(_0640_),
    .B2(_0603_),
    .ZN(_0641_));
 MUX2_X1 _3233_ (.A(_0638_),
    .B(_0641_),
    .S(_0538_),
    .Z(_0642_));
 NAND4_X1 _3234_ (.A1(_0550_),
    .A2(_0547_),
    .A3(_0576_),
    .A4(_0603_),
    .ZN(_0643_));
 OAI21_X1 _3235_ (.A(_0642_),
    .B1(_0643_),
    .B2(_0540_),
    .ZN(_0644_));
 OAI21_X1 _3236_ (.A(_0635_),
    .B1(_0644_),
    .B2(_0542_),
    .ZN(_0645_));
 XNOR2_X1 _3237_ (.A(_0623_),
    .B(_0645_),
    .ZN(_0646_));
 NOR2_X1 _3238_ (.A1(_0433_),
    .A2(_0646_),
    .ZN(_0093_));
 CLKBUF_X3 _3239_ (.A(_2270_),
    .Z(_0647_));
 NOR2_X1 _3240_ (.A1(_0622_),
    .A2(_0633_),
    .ZN(_0648_));
 AOI21_X1 _3241_ (.A(_2266_),
    .B1(_0631_),
    .B2(_0648_),
    .ZN(_0649_));
 INV_X1 _3242_ (.A(_2264_),
    .ZN(_0650_));
 AOI21_X1 _3243_ (.A(_2248_),
    .B1(_2240_),
    .B2(_0576_),
    .ZN(_0651_));
 NOR2_X1 _3244_ (.A1(_0604_),
    .A2(_0651_),
    .ZN(_0652_));
 OAI21_X1 _3245_ (.A(_0622_),
    .B1(_2256_),
    .B2(_0652_),
    .ZN(_0653_));
 NAND3_X1 _3246_ (.A1(_0412_),
    .A2(_0650_),
    .A3(_0653_),
    .ZN(_0654_));
 AOI21_X1 _3247_ (.A(_2261_),
    .B1(_2253_),
    .B2(_0622_),
    .ZN(_0655_));
 NAND2_X1 _3248_ (.A1(_0603_),
    .A2(_0622_),
    .ZN(_0656_));
 AOI21_X1 _3249_ (.A(_2245_),
    .B1(_2237_),
    .B2(_0576_),
    .ZN(_0657_));
 OAI21_X1 _3250_ (.A(_0655_),
    .B1(_0656_),
    .B2(_0657_),
    .ZN(_0658_));
 OAI21_X1 _3251_ (.A(_0654_),
    .B1(_0658_),
    .B2(_0412_),
    .ZN(_0659_));
 NAND4_X1 _3252_ (.A1(_0547_),
    .A2(_0576_),
    .A3(_0603_),
    .A4(_0622_),
    .ZN(_0660_));
 OAI21_X1 _3253_ (.A(_0659_),
    .B1(_0660_),
    .B2(_0569_),
    .ZN(_0661_));
 MUX2_X1 _3254_ (.A(_0649_),
    .B(_0661_),
    .S(_0571_),
    .Z(_0662_));
 XNOR2_X1 _3255_ (.A(_0647_),
    .B(_0662_),
    .ZN(_0663_));
 NOR2_X1 _3256_ (.A1(_0433_),
    .A2(_0663_),
    .ZN(_0094_));
 CLKBUF_X3 _3257_ (.A(_2278_),
    .Z(_0664_));
 INV_X1 _3258_ (.A(_0664_),
    .ZN(_0665_));
 INV_X1 _3259_ (.A(_2274_),
    .ZN(_0666_));
 OAI21_X1 _3260_ (.A(_0666_),
    .B1(_0649_),
    .B2(_0647_),
    .ZN(_0667_));
 AOI21_X1 _3261_ (.A(_2256_),
    .B1(_2248_),
    .B2(_0603_),
    .ZN(_0668_));
 OAI21_X1 _3262_ (.A(_0650_),
    .B1(_0668_),
    .B2(_0623_),
    .ZN(_0669_));
 AOI21_X1 _3263_ (.A(_2272_),
    .B1(_0669_),
    .B2(_0647_),
    .ZN(_0670_));
 INV_X1 _3264_ (.A(_2261_),
    .ZN(_0671_));
 AOI21_X1 _3265_ (.A(_2253_),
    .B1(_2245_),
    .B2(_0603_),
    .ZN(_0672_));
 OAI21_X1 _3266_ (.A(_0671_),
    .B1(_0672_),
    .B2(_0623_),
    .ZN(_0673_));
 AOI21_X1 _3267_ (.A(_2269_),
    .B1(_0673_),
    .B2(_0647_),
    .ZN(_0674_));
 MUX2_X1 _3268_ (.A(_0670_),
    .B(_0674_),
    .S(_0538_),
    .Z(_0675_));
 NAND4_X1 _3269_ (.A1(_0576_),
    .A2(_0603_),
    .A3(_0622_),
    .A4(_0647_),
    .ZN(_0676_));
 OR2_X1 _3270_ (.A1(_0592_),
    .A2(_0676_),
    .ZN(_0677_));
 AND2_X1 _3271_ (.A1(_0675_),
    .A2(_0677_),
    .ZN(_0678_));
 MUX2_X1 _3272_ (.A(_0667_),
    .B(_0678_),
    .S(_0571_),
    .Z(_0679_));
 XNOR2_X1 _3273_ (.A(_0665_),
    .B(_0679_),
    .ZN(_0680_));
 NOR2_X1 _3274_ (.A1(_0433_),
    .A2(_0680_),
    .ZN(_0095_));
 CLKBUF_X3 _3275_ (.A(_2286_),
    .Z(_0681_));
 INV_X1 _3276_ (.A(_2282_),
    .ZN(_0682_));
 NOR2_X1 _3277_ (.A1(_0682_),
    .A2(_0500_),
    .ZN(_0683_));
 NOR2_X1 _3278_ (.A1(_0664_),
    .A2(_0499_),
    .ZN(_0684_));
 AOI21_X1 _3279_ (.A(_2280_),
    .B1(_2272_),
    .B2(_0664_),
    .ZN(_0685_));
 NAND2_X1 _3280_ (.A1(_0647_),
    .A2(_0664_),
    .ZN(_0686_));
 AOI21_X1 _3281_ (.A(_2264_),
    .B1(_2256_),
    .B2(_0622_),
    .ZN(_0687_));
 OAI21_X1 _3282_ (.A(_0685_),
    .B1(_0686_),
    .B2(_0687_),
    .ZN(_0688_));
 AND2_X1 _3283_ (.A1(_0411_),
    .A2(_0688_),
    .ZN(_0689_));
 NOR2_X1 _3284_ (.A1(_0656_),
    .A2(_0686_),
    .ZN(_0690_));
 OR3_X1 _3285_ (.A1(_0611_),
    .A2(_0616_),
    .A3(_0618_),
    .ZN(_0691_));
 AOI21_X1 _3286_ (.A(_2277_),
    .B1(_2269_),
    .B2(_0664_),
    .ZN(_0692_));
 OAI21_X1 _3287_ (.A(_0692_),
    .B1(_0686_),
    .B2(_0655_),
    .ZN(_0693_));
 AOI221_X2 _3288_ (.A(_0689_),
    .B1(_0690_),
    .B2(_0691_),
    .C1(_0693_),
    .C2(_0538_),
    .ZN(_0694_));
 AOI221_X2 _3289_ (.A(_0683_),
    .B1(_0684_),
    .B2(_0667_),
    .C1(_0500_),
    .C2(_0694_),
    .ZN(_0695_));
 XNOR2_X1 _3290_ (.A(_0681_),
    .B(_0695_),
    .ZN(_0696_));
 NOR2_X1 _3291_ (.A1(_0433_),
    .A2(_0696_),
    .ZN(_0096_));
 BUF_X2 _3292_ (.A(_2294_),
    .Z(_0697_));
 INV_X1 _3293_ (.A(_2280_),
    .ZN(_0698_));
 AOI21_X1 _3294_ (.A(_2272_),
    .B1(_2264_),
    .B2(_2270_),
    .ZN(_0699_));
 OAI21_X1 _3295_ (.A(_0698_),
    .B1(_0699_),
    .B2(_0665_),
    .ZN(_0700_));
 AOI21_X1 _3296_ (.A(_2288_),
    .B1(_0700_),
    .B2(_0681_),
    .ZN(_0701_));
 INV_X1 _3297_ (.A(_2277_),
    .ZN(_0702_));
 AOI21_X1 _3298_ (.A(_2269_),
    .B1(_2261_),
    .B2(_0647_),
    .ZN(_0703_));
 OAI21_X1 _3299_ (.A(_0702_),
    .B1(_0703_),
    .B2(_0665_),
    .ZN(_0704_));
 AOI21_X1 _3300_ (.A(_2285_),
    .B1(_0704_),
    .B2(_0681_),
    .ZN(_0705_));
 MUX2_X1 _3301_ (.A(_0701_),
    .B(_0705_),
    .S(_0538_),
    .Z(_0706_));
 AND3_X1 _3302_ (.A1(_0642_),
    .A2(_0643_),
    .A3(_0706_),
    .ZN(_0707_));
 NAND4_X1 _3303_ (.A1(_0622_),
    .A2(_0647_),
    .A3(_0664_),
    .A4(_0681_),
    .ZN(_0708_));
 AND3_X1 _3304_ (.A1(_0539_),
    .A2(_0642_),
    .A3(_0706_),
    .ZN(_0709_));
 AOI221_X2 _3305_ (.A(_0707_),
    .B1(_0708_),
    .B2(_0706_),
    .C1(_0529_),
    .C2(_0709_),
    .ZN(_0710_));
 NAND2_X1 _3306_ (.A1(_0501_),
    .A2(_0710_),
    .ZN(_0711_));
 INV_X1 _3307_ (.A(_0647_),
    .ZN(_0712_));
 AOI21_X1 _3308_ (.A(_2274_),
    .B1(_0712_),
    .B2(_2266_),
    .ZN(_0713_));
 OAI21_X1 _3309_ (.A(_0682_),
    .B1(_0713_),
    .B2(_0664_),
    .ZN(_0714_));
 INV_X1 _3310_ (.A(_0681_),
    .ZN(_0715_));
 AOI21_X1 _3311_ (.A(_2290_),
    .B1(_0714_),
    .B2(_0715_),
    .ZN(_0716_));
 NAND3_X1 _3312_ (.A1(_0712_),
    .A2(_0665_),
    .A3(_0715_),
    .ZN(_0717_));
 NAND2_X1 _3313_ (.A1(_0631_),
    .A2(_0648_),
    .ZN(_0718_));
 OAI21_X1 _3314_ (.A(_0716_),
    .B1(_0717_),
    .B2(_0718_),
    .ZN(_0719_));
 OAI21_X1 _3315_ (.A(_0711_),
    .B1(_0719_),
    .B2(_0501_),
    .ZN(_0720_));
 XNOR2_X1 _3316_ (.A(_0697_),
    .B(_0720_),
    .ZN(_0721_));
 NOR2_X1 _3317_ (.A1(_0433_),
    .A2(_0721_),
    .ZN(_0097_));
 BUF_X2 _3318_ (.A(_2302_),
    .Z(_0722_));
 NOR2_X1 _3319_ (.A1(_0722_),
    .A2(_0432_),
    .ZN(_0723_));
 INV_X1 _3320_ (.A(_0722_),
    .ZN(_0724_));
 BUF_X2 _3321_ (.A(_0724_),
    .Z(_0725_));
 NOR2_X1 _3322_ (.A1(_0725_),
    .A2(_0432_),
    .ZN(_0726_));
 INV_X1 _3323_ (.A(_0697_),
    .ZN(_0727_));
 AOI21_X1 _3324_ (.A(_2298_),
    .B1(_0719_),
    .B2(_0727_),
    .ZN(_0728_));
 NAND4_X1 _3325_ (.A1(_0647_),
    .A2(_0664_),
    .A3(_0681_),
    .A4(_0697_),
    .ZN(_0729_));
 INV_X1 _3326_ (.A(_0729_),
    .ZN(_0730_));
 AND2_X1 _3327_ (.A1(_0661_),
    .A2(_0730_),
    .ZN(_0731_));
 INV_X1 _3328_ (.A(_2288_),
    .ZN(_0732_));
 OAI21_X1 _3329_ (.A(_0732_),
    .B1(_0685_),
    .B2(_0715_),
    .ZN(_0733_));
 AOI21_X1 _3330_ (.A(_2296_),
    .B1(_0733_),
    .B2(_0697_),
    .ZN(_0734_));
 INV_X1 _3331_ (.A(_2285_),
    .ZN(_0735_));
 OAI21_X1 _3332_ (.A(_0735_),
    .B1(_0692_),
    .B2(_0715_),
    .ZN(_0736_));
 AOI21_X1 _3333_ (.A(_2293_),
    .B1(_0736_),
    .B2(_0697_),
    .ZN(_0737_));
 CLKBUF_X3 _3334_ (.A(_0538_),
    .Z(_0738_));
 MUX2_X1 _3335_ (.A(_0734_),
    .B(_0737_),
    .S(_0738_),
    .Z(_0739_));
 NAND2_X1 _3336_ (.A1(_0571_),
    .A2(_0739_),
    .ZN(_0740_));
 OAI22_X1 _3337_ (.A1(_0501_),
    .A2(_0728_),
    .B1(_0731_),
    .B2(_0740_),
    .ZN(_0741_));
 MUX2_X1 _3338_ (.A(_0723_),
    .B(_0726_),
    .S(_0741_),
    .Z(_0098_));
 CLKBUF_X3 _3339_ (.A(_0432_),
    .Z(_0742_));
 CLKBUF_X3 _3340_ (.A(_2310_),
    .Z(_0743_));
 NAND2_X1 _3341_ (.A1(_2298_),
    .A2(_0725_),
    .ZN(_0744_));
 NAND2_X1 _3342_ (.A1(_0727_),
    .A2(_0724_),
    .ZN(_0745_));
 OAI21_X1 _3343_ (.A(_0744_),
    .B1(_0745_),
    .B2(_0716_),
    .ZN(_0746_));
 OR4_X1 _3344_ (.A1(_0622_),
    .A2(_0633_),
    .A3(_0717_),
    .A4(_0745_),
    .ZN(_0747_));
 INV_X1 _3345_ (.A(_0747_),
    .ZN(_0748_));
 AOI211_X2 _3346_ (.A(_2306_),
    .B(_0746_),
    .C1(_0748_),
    .C2(_0631_),
    .ZN(_0749_));
 INV_X1 _3347_ (.A(_2296_),
    .ZN(_0750_));
 AOI21_X1 _3348_ (.A(_2288_),
    .B1(_2280_),
    .B2(_0681_),
    .ZN(_0751_));
 OAI21_X1 _3349_ (.A(_0750_),
    .B1(_0751_),
    .B2(_0727_),
    .ZN(_0752_));
 AOI21_X1 _3350_ (.A(_2304_),
    .B1(_0752_),
    .B2(_0722_),
    .ZN(_0753_));
 INV_X1 _3351_ (.A(_2293_),
    .ZN(_0754_));
 AOI21_X1 _3352_ (.A(_2285_),
    .B1(_2277_),
    .B2(_0681_),
    .ZN(_0755_));
 OAI21_X1 _3353_ (.A(_0754_),
    .B1(_0755_),
    .B2(_0727_),
    .ZN(_0756_));
 AOI21_X1 _3354_ (.A(_2301_),
    .B1(_0756_),
    .B2(_0722_),
    .ZN(_0757_));
 MUX2_X1 _3355_ (.A(_0753_),
    .B(_0757_),
    .S(_0538_),
    .Z(_0758_));
 NAND4_X2 _3356_ (.A1(_0664_),
    .A2(_0681_),
    .A3(_0697_),
    .A4(_0722_),
    .ZN(_0759_));
 OR2_X1 _3357_ (.A1(_0676_),
    .A2(_0759_),
    .ZN(_0760_));
 OAI221_X2 _3358_ (.A(_0758_),
    .B1(_0759_),
    .B2(_0675_),
    .C1(_0760_),
    .C2(_0592_),
    .ZN(_0761_));
 MUX2_X1 _3359_ (.A(_0749_),
    .B(_0761_),
    .S(_0500_),
    .Z(_0762_));
 XNOR2_X1 _3360_ (.A(_0743_),
    .B(_0762_),
    .ZN(_0763_));
 NOR2_X1 _3361_ (.A1(_0742_),
    .A2(_0763_),
    .ZN(_0099_));
 BUF_X2 _3362_ (.A(_2318_),
    .Z(_0764_));
 NOR2_X1 _3363_ (.A1(_0764_),
    .A2(_0432_),
    .ZN(_0765_));
 INV_X2 _3364_ (.A(_0764_),
    .ZN(_0766_));
 NOR2_X1 _3365_ (.A1(_0766_),
    .A2(_0432_),
    .ZN(_0767_));
 INV_X1 _3366_ (.A(_2314_),
    .ZN(_0768_));
 OAI21_X1 _3367_ (.A(_0768_),
    .B1(_0749_),
    .B2(_0743_),
    .ZN(_0769_));
 INV_X1 _3368_ (.A(_2304_),
    .ZN(_0770_));
 AOI21_X1 _3369_ (.A(_2296_),
    .B1(_2288_),
    .B2(_0697_),
    .ZN(_0771_));
 OAI21_X1 _3370_ (.A(_0770_),
    .B1(_0771_),
    .B2(_0725_),
    .ZN(_0772_));
 AOI21_X1 _3371_ (.A(_2312_),
    .B1(_0772_),
    .B2(_0743_),
    .ZN(_0773_));
 NAND2_X1 _3372_ (.A1(_0412_),
    .A2(_0773_),
    .ZN(_0774_));
 INV_X1 _3373_ (.A(_2301_),
    .ZN(_0775_));
 AOI21_X1 _3374_ (.A(_2293_),
    .B1(_2285_),
    .B2(_0697_),
    .ZN(_0776_));
 OAI21_X1 _3375_ (.A(_0775_),
    .B1(_0776_),
    .B2(_0725_),
    .ZN(_0777_));
 AOI21_X1 _3376_ (.A(_2309_),
    .B1(_0777_),
    .B2(_0743_),
    .ZN(_0778_));
 NAND2_X1 _3377_ (.A1(_0738_),
    .A2(_0778_),
    .ZN(_0779_));
 INV_X1 _3378_ (.A(_0743_),
    .ZN(_0780_));
 NOR4_X1 _3379_ (.A1(_0715_),
    .A2(_0727_),
    .A3(_0725_),
    .A4(_0780_),
    .ZN(_0781_));
 AOI21_X1 _3380_ (.A(_0689_),
    .B1(_0693_),
    .B2(_0738_),
    .ZN(_0782_));
 OR2_X1 _3381_ (.A1(_0656_),
    .A2(_0686_),
    .ZN(_0783_));
 OAI21_X1 _3382_ (.A(_0782_),
    .B1(_0783_),
    .B2(_0619_),
    .ZN(_0784_));
 AOI22_X2 _3383_ (.A1(_0774_),
    .A2(_0779_),
    .B1(_0781_),
    .B2(_0784_),
    .ZN(_0785_));
 MUX2_X1 _3384_ (.A(_0769_),
    .B(_0785_),
    .S(_0571_),
    .Z(_0786_));
 MUX2_X1 _3385_ (.A(_0765_),
    .B(_0767_),
    .S(_0786_),
    .Z(_0100_));
 BUF_X2 _3386_ (.A(_2326_),
    .Z(_0787_));
 AOI21_X1 _3387_ (.A(_2322_),
    .B1(_0766_),
    .B2(_2314_),
    .ZN(_0788_));
 AND2_X1 _3388_ (.A1(_0465_),
    .A2(_0788_),
    .ZN(_0789_));
 NAND2_X1 _3389_ (.A1(_0780_),
    .A2(_0766_),
    .ZN(_0790_));
 OAI21_X1 _3390_ (.A(_0789_),
    .B1(_0790_),
    .B2(_0749_),
    .ZN(_0791_));
 INV_X1 _3391_ (.A(_2320_),
    .ZN(_0792_));
 OAI21_X1 _3392_ (.A(_0770_),
    .B1(_0750_),
    .B2(_0725_),
    .ZN(_0793_));
 AOI21_X1 _3393_ (.A(_2312_),
    .B1(_0793_),
    .B2(_0743_),
    .ZN(_0794_));
 OAI21_X1 _3394_ (.A(_0792_),
    .B1(_0794_),
    .B2(_0766_),
    .ZN(_0795_));
 INV_X1 _3395_ (.A(_2317_),
    .ZN(_0796_));
 OAI21_X1 _3396_ (.A(_0775_),
    .B1(_0754_),
    .B2(_0725_),
    .ZN(_0797_));
 AOI21_X1 _3397_ (.A(_2309_),
    .B1(_0797_),
    .B2(_0743_),
    .ZN(_0798_));
 OAI21_X1 _3398_ (.A(_0796_),
    .B1(_0798_),
    .B2(_0766_),
    .ZN(_0799_));
 MUX2_X1 _3399_ (.A(_0795_),
    .B(_0799_),
    .S(_0738_),
    .Z(_0800_));
 NOR4_X1 _3400_ (.A1(_0727_),
    .A2(_0725_),
    .A3(_0780_),
    .A4(_0766_),
    .ZN(_0801_));
 AOI21_X1 _3401_ (.A(_0800_),
    .B1(_0801_),
    .B2(_0710_),
    .ZN(_0802_));
 OAI21_X1 _3402_ (.A(_0791_),
    .B1(_0802_),
    .B2(_0542_),
    .ZN(_0803_));
 XNOR2_X1 _3403_ (.A(_0787_),
    .B(_0803_),
    .ZN(_0804_));
 NOR2_X1 _3404_ (.A1(_0742_),
    .A2(_0804_),
    .ZN(_0101_));
 BUF_X2 _3405_ (.A(_2334_),
    .Z(_0805_));
 INV_X1 _3406_ (.A(_0805_),
    .ZN(_0806_));
 NOR3_X1 _3407_ (.A1(_0738_),
    .A2(_2320_),
    .A3(_2328_),
    .ZN(_0807_));
 OAI21_X1 _3408_ (.A(_0770_),
    .B1(_0734_),
    .B2(_0725_),
    .ZN(_0808_));
 AOI21_X1 _3409_ (.A(_2312_),
    .B1(_0808_),
    .B2(_0743_),
    .ZN(_0809_));
 OAI21_X1 _3410_ (.A(_0807_),
    .B1(_0809_),
    .B2(_0766_),
    .ZN(_0810_));
 NOR3_X1 _3411_ (.A1(_0411_),
    .A2(_2317_),
    .A3(_2325_),
    .ZN(_0811_));
 OAI21_X1 _3412_ (.A(_0775_),
    .B1(_0737_),
    .B2(_0725_),
    .ZN(_0812_));
 AOI21_X1 _3413_ (.A(_2309_),
    .B1(_0812_),
    .B2(_0743_),
    .ZN(_0813_));
 OAI21_X1 _3414_ (.A(_0811_),
    .B1(_0813_),
    .B2(_0766_),
    .ZN(_0814_));
 INV_X2 _3415_ (.A(_0787_),
    .ZN(_0815_));
 INV_X1 _3416_ (.A(_2325_),
    .ZN(_0816_));
 NAND3_X1 _3417_ (.A1(_0738_),
    .A2(_0815_),
    .A3(_0816_),
    .ZN(_0817_));
 INV_X1 _3418_ (.A(_2328_),
    .ZN(_0818_));
 NAND3_X1 _3419_ (.A1(_0412_),
    .A2(_0815_),
    .A3(_0818_),
    .ZN(_0819_));
 AND4_X1 _3420_ (.A1(_0810_),
    .A2(_0814_),
    .A3(_0817_),
    .A4(_0819_),
    .ZN(_0820_));
 NAND4_X1 _3421_ (.A1(_0722_),
    .A2(_0743_),
    .A3(_0764_),
    .A4(_0787_),
    .ZN(_0821_));
 NOR3_X1 _3422_ (.A1(_0465_),
    .A2(_0729_),
    .A3(_0821_),
    .ZN(_0822_));
 AOI22_X1 _3423_ (.A1(_0571_),
    .A2(_0820_),
    .B1(_0822_),
    .B2(_0661_),
    .ZN(_0823_));
 NOR2_X1 _3424_ (.A1(_2330_),
    .A2(_0499_),
    .ZN(_0824_));
 NAND2_X1 _3425_ (.A1(_0788_),
    .A2(_0824_),
    .ZN(_0825_));
 INV_X1 _3426_ (.A(_0825_),
    .ZN(_0826_));
 OR2_X1 _3427_ (.A1(_0749_),
    .A2(_0790_),
    .ZN(_0827_));
 AOI22_X1 _3428_ (.A1(_0787_),
    .A2(_0824_),
    .B1(_0826_),
    .B2(_0827_),
    .ZN(_0828_));
 AND3_X1 _3429_ (.A1(_0806_),
    .A2(_0823_),
    .A3(_0828_),
    .ZN(_0829_));
 AOI21_X1 _3430_ (.A(_0806_),
    .B1(_0823_),
    .B2(_0828_),
    .ZN(_0830_));
 NOR3_X1 _3431_ (.A1(_0742_),
    .A2(_0829_),
    .A3(_0830_),
    .ZN(_0102_));
 CLKBUF_X2 _3432_ (.A(_2342_),
    .Z(_0831_));
 NOR4_X1 _3433_ (.A1(_0764_),
    .A2(_0787_),
    .A3(_0805_),
    .A4(_0831_),
    .ZN(_0832_));
 NAND2_X1 _3434_ (.A1(_0769_),
    .A2(_0832_),
    .ZN(_0833_));
 OR2_X1 _3435_ (.A1(_2346_),
    .A2(_0500_),
    .ZN(_0834_));
 INV_X1 _3436_ (.A(_2338_),
    .ZN(_0835_));
 AOI21_X1 _3437_ (.A(_2330_),
    .B1(_0815_),
    .B2(_2322_),
    .ZN(_0836_));
 OAI21_X1 _3438_ (.A(_0835_),
    .B1(_0836_),
    .B2(_0805_),
    .ZN(_0837_));
 INV_X1 _3439_ (.A(_0831_),
    .ZN(_0838_));
 AOI21_X1 _3440_ (.A(_0834_),
    .B1(_0837_),
    .B2(_0838_),
    .ZN(_0839_));
 OAI21_X1 _3441_ (.A(_0818_),
    .B1(_0792_),
    .B2(_0815_),
    .ZN(_0840_));
 AOI21_X1 _3442_ (.A(_2336_),
    .B1(_0840_),
    .B2(_0805_),
    .ZN(_0841_));
 NOR2_X1 _3443_ (.A1(_0838_),
    .A2(_0841_),
    .ZN(_0842_));
 OAI21_X1 _3444_ (.A(_0412_),
    .B1(_2344_),
    .B2(_0842_),
    .ZN(_0843_));
 NAND4_X1 _3445_ (.A1(_0764_),
    .A2(_0787_),
    .A3(_0805_),
    .A4(_0831_),
    .ZN(_0844_));
 INV_X1 _3446_ (.A(_2333_),
    .ZN(_0845_));
 AOI21_X1 _3447_ (.A(_2325_),
    .B1(_2317_),
    .B2(_0787_),
    .ZN(_0846_));
 OAI21_X1 _3448_ (.A(_0845_),
    .B1(_0846_),
    .B2(_0806_),
    .ZN(_0847_));
 AOI21_X1 _3449_ (.A(_2341_),
    .B1(_0847_),
    .B2(_0831_),
    .ZN(_0848_));
 OAI221_X2 _3450_ (.A(_0843_),
    .B1(_0844_),
    .B2(_0785_),
    .C1(_0848_),
    .C2(_0412_),
    .ZN(_0849_));
 AOI221_X2 _3451_ (.A(_0432_),
    .B1(_0833_),
    .B2(_0839_),
    .C1(_0849_),
    .C2(_0501_),
    .ZN(_0104_));
 OR2_X1 _3452_ (.A1(_0482_),
    .A2(_0485_),
    .ZN(_0850_));
 MUX2_X1 _3453_ (.A(_0454_),
    .B(_0850_),
    .S(_0500_),
    .Z(_0851_));
 XNOR2_X1 _3454_ (.A(_0455_),
    .B(_0851_),
    .ZN(_0852_));
 NOR2_X1 _3455_ (.A1(_0742_),
    .A2(_0852_),
    .ZN(_0105_));
 NOR3_X1 _3456_ (.A1(_1586_),
    .A2(_0419_),
    .A3(_0387_),
    .ZN(_0853_));
 NOR3_X1 _3457_ (.A1(_0738_),
    .A2(_2152_),
    .A3(_0524_),
    .ZN(_0854_));
 NOR3_X1 _3458_ (.A1(_0412_),
    .A2(_2149_),
    .A3(_0518_),
    .ZN(_0855_));
 OAI21_X1 _3459_ (.A(_0571_),
    .B1(_0854_),
    .B2(_0855_),
    .ZN(_0856_));
 OAI21_X1 _3460_ (.A(_0856_),
    .B1(_0501_),
    .B2(_0456_),
    .ZN(_0857_));
 XNOR2_X1 _3461_ (.A(_0447_),
    .B(_0857_),
    .ZN(_0858_));
 AND2_X1 _3462_ (.A1(_0853_),
    .A2(_0858_),
    .ZN(_0106_));
 NOR2_X1 _3463_ (.A1(_0447_),
    .A2(_0456_),
    .ZN(_0859_));
 NOR2_X1 _3464_ (.A1(_2170_),
    .A2(_0859_),
    .ZN(_0860_));
 NAND3_X1 _3465_ (.A1(_0412_),
    .A2(_0494_),
    .A3(_0555_),
    .ZN(_0861_));
 NAND3_X1 _3466_ (.A1(_0738_),
    .A2(_0491_),
    .A3(_0560_),
    .ZN(_0862_));
 AND2_X1 _3467_ (.A1(_0861_),
    .A2(_0862_),
    .ZN(_0863_));
 MUX2_X1 _3468_ (.A(_0860_),
    .B(_0863_),
    .S(_0500_),
    .Z(_0864_));
 XNOR2_X1 _3469_ (.A(_0448_),
    .B(_0864_),
    .ZN(_0865_));
 NOR2_X1 _3470_ (.A1(_0742_),
    .A2(_0865_),
    .ZN(_0107_));
 NOR2_X1 _3471_ (.A1(_0524_),
    .A2(_0525_),
    .ZN(_0866_));
 OR3_X1 _3472_ (.A1(_0542_),
    .A2(_0520_),
    .A3(_0866_),
    .ZN(_0867_));
 INV_X1 _3473_ (.A(_2178_),
    .ZN(_0868_));
 OAI21_X1 _3474_ (.A(_0868_),
    .B1(_0860_),
    .B2(_0448_),
    .ZN(_0869_));
 OAI21_X1 _3475_ (.A(_0867_),
    .B1(_0869_),
    .B2(_0501_),
    .ZN(_0870_));
 XNOR2_X1 _3476_ (.A(_0449_),
    .B(_0870_),
    .ZN(_0871_));
 NOR2_X1 _3477_ (.A1(_0742_),
    .A2(_0871_),
    .ZN(_0108_));
 OR2_X1 _3478_ (.A1(_0628_),
    .A2(_0461_),
    .ZN(_0872_));
 NOR2_X1 _3479_ (.A1(_0872_),
    .A2(_0571_),
    .ZN(_0873_));
 OR2_X1 _3480_ (.A1(_0496_),
    .A2(_0488_),
    .ZN(_0874_));
 AOI21_X1 _3481_ (.A(_0873_),
    .B1(_0874_),
    .B2(_0501_),
    .ZN(_0875_));
 XNOR2_X1 _3482_ (.A(_0442_),
    .B(_0875_),
    .ZN(_0876_));
 NOR2_X1 _3483_ (.A1(_0742_),
    .A2(_0876_),
    .ZN(_0109_));
 AOI21_X1 _3484_ (.A(_2194_),
    .B1(_0872_),
    .B2(_0442_),
    .ZN(_0877_));
 MUX2_X1 _3485_ (.A(_0527_),
    .B(_0877_),
    .S(_0542_),
    .Z(_0878_));
 XNOR2_X1 _3486_ (.A(_0444_),
    .B(_0878_),
    .ZN(_0879_));
 NOR2_X1 _3487_ (.A1(_0742_),
    .A2(_0879_),
    .ZN(_0110_));
 OAI21_X1 _3488_ (.A(_0445_),
    .B1(_0628_),
    .B2(_0629_),
    .ZN(_0880_));
 NAND2_X1 _3489_ (.A1(_0880_),
    .A2(_0542_),
    .ZN(_0881_));
 NAND3_X1 _3490_ (.A1(_0412_),
    .A2(_0468_),
    .A3(_0558_),
    .ZN(_0882_));
 NAND3_X1 _3491_ (.A1(_0738_),
    .A2(_0473_),
    .A3(_0563_),
    .ZN(_0883_));
 NAND2_X1 _3492_ (.A1(_0882_),
    .A2(_0883_),
    .ZN(_0884_));
 OAI21_X1 _3493_ (.A(_0881_),
    .B1(_0884_),
    .B2(_0542_),
    .ZN(_0885_));
 XNOR2_X1 _3494_ (.A(_0439_),
    .B(_0885_),
    .ZN(_0886_));
 NOR2_X1 _3495_ (.A1(_0742_),
    .A2(_0886_),
    .ZN(_0111_));
 NOR2_X1 _3496_ (.A1(_2210_),
    .A2(_0463_),
    .ZN(_0887_));
 AND2_X1 _3497_ (.A1(_0527_),
    .A2(_0528_),
    .ZN(_0888_));
 NAND2_X1 _3498_ (.A1(_0571_),
    .A2(_0586_),
    .ZN(_0889_));
 OAI22_X1 _3499_ (.A1(_0887_),
    .A2(_0501_),
    .B1(_0888_),
    .B2(_0889_),
    .ZN(_0890_));
 XNOR2_X1 _3500_ (.A(_0438_),
    .B(_0890_),
    .ZN(_0891_));
 NOR2_X1 _3501_ (.A1(_0742_),
    .A2(_0891_),
    .ZN(_0112_));
 CLKBUF_X3 _3502_ (.A(_2033_),
    .Z(_0892_));
 INV_X1 _3503_ (.A(_0892_),
    .ZN(_0893_));
 CLKBUF_X3 _3504_ (.A(_2039_),
    .Z(_0894_));
 NAND3_X2 _3505_ (.A1(_0894_),
    .A2(_1999_),
    .A3(_2044_),
    .ZN(_0895_));
 AOI21_X4 _3506_ (.A(_2041_),
    .B1(_2045_),
    .B2(_0894_),
    .ZN(_0896_));
 NAND2_X1 _3507_ (.A1(_0895_),
    .A2(_0896_),
    .ZN(_0897_));
 AND3_X1 _3508_ (.A1(_0894_),
    .A2(_1995_),
    .A3(_2044_),
    .ZN(_0898_));
 AOI21_X1 _3509_ (.A(_2038_),
    .B1(_2043_),
    .B2(_0894_),
    .ZN(_0899_));
 INV_X1 _3510_ (.A(_0899_),
    .ZN(_0900_));
 OR2_X1 _3511_ (.A1(_0898_),
    .A2(_0900_),
    .ZN(_0901_));
 BUF_X2 _3512_ (.A(_2015_),
    .Z(_0902_));
 BUF_X4 _3513_ (.A(_2027_),
    .Z(_0903_));
 CLKBUF_X3 _3514_ (.A(_2021_),
    .Z(_0904_));
 NAND4_X4 _3515_ (.A1(_0902_),
    .A2(_0903_),
    .A3(_0892_),
    .A4(_0904_),
    .ZN(_0905_));
 BUF_X2 _3516_ (.A(_2009_),
    .Z(_0906_));
 NAND4_X4 _3517_ (.A1(_0894_),
    .A2(_2118_),
    .A3(_0906_),
    .A4(_2044_),
    .ZN(_0907_));
 NOR2_X2 _3518_ (.A1(_0905_),
    .A2(_0907_),
    .ZN(_0908_));
 INV_X1 _3519_ (.A(_2017_),
    .ZN(_0909_));
 AND2_X1 _3520_ (.A1(_0903_),
    .A2(_2035_),
    .ZN(_0910_));
 NOR3_X2 _3521_ (.A1(_2023_),
    .A2(_2029_),
    .A3(_0910_),
    .ZN(_0911_));
 OAI21_X2 _3522_ (.A(_0902_),
    .B1(_0904_),
    .B2(_2023_),
    .ZN(_0912_));
 OAI21_X4 _3523_ (.A(_0909_),
    .B1(_0911_),
    .B2(_0912_),
    .ZN(_0913_));
 AOI21_X4 _3524_ (.A(_0905_),
    .B1(_0896_),
    .B2(_0895_),
    .ZN(_0914_));
 OR4_X4 _3525_ (.A1(_2011_),
    .A2(_0908_),
    .A3(_0913_),
    .A4(_0914_),
    .ZN(_0915_));
 NOR2_X2 _3526_ (.A1(_2011_),
    .A2(_0906_),
    .ZN(_0916_));
 INV_X1 _3527_ (.A(_2097_),
    .ZN(_0917_));
 NAND3_X2 _3528_ (.A1(_2112_),
    .A2(_2109_),
    .A3(_2115_),
    .ZN(_0918_));
 NOR2_X2 _3529_ (.A1(_0917_),
    .A2(_0918_),
    .ZN(_0919_));
 INV_X1 _3530_ (.A(_2114_),
    .ZN(_0920_));
 INV_X1 _3531_ (.A(_2096_),
    .ZN(_0921_));
 AOI21_X1 _3532_ (.A(_2108_),
    .B1(_2111_),
    .B2(_2109_),
    .ZN(_0922_));
 INV_X1 _3533_ (.A(_2115_),
    .ZN(_0923_));
 OAI221_X2 _3534_ (.A(_0920_),
    .B1(_0921_),
    .B2(_0918_),
    .C1(_0922_),
    .C2(_0923_),
    .ZN(_0924_));
 NOR4_X4 _3535_ (.A1(_0919_),
    .A2(_0905_),
    .A3(_0907_),
    .A4(_0924_),
    .ZN(_0925_));
 NOR2_X4 _3536_ (.A1(_0916_),
    .A2(_0925_),
    .ZN(_0926_));
 NAND4_X4 _3537_ (.A1(_2073_),
    .A2(_2100_),
    .A3(_2103_),
    .A4(_2106_),
    .ZN(_0927_));
 INV_X1 _3538_ (.A(_0927_),
    .ZN(_0928_));
 INV_X1 _3539_ (.A(_2084_),
    .ZN(_0929_));
 NAND3_X2 _3540_ (.A1(_2076_),
    .A2(_2079_),
    .A3(_2082_),
    .ZN(_0930_));
 AOI21_X1 _3541_ (.A(_2078_),
    .B1(_2081_),
    .B2(_2079_),
    .ZN(_0931_));
 INV_X1 _3542_ (.A(_2076_),
    .ZN(_0932_));
 OAI22_X1 _3543_ (.A1(_0929_),
    .A2(_0930_),
    .B1(_0931_),
    .B2(_0932_),
    .ZN(_0933_));
 OAI21_X2 _3544_ (.A(_0928_),
    .B1(_0933_),
    .B2(_2075_),
    .ZN(_0934_));
 INV_X1 _3545_ (.A(_2085_),
    .ZN(_0935_));
 NAND4_X2 _3546_ (.A1(_2061_),
    .A2(_2088_),
    .A3(_2091_),
    .A4(_2094_),
    .ZN(_0936_));
 NOR4_X4 _3547_ (.A1(_0935_),
    .A2(_0927_),
    .A3(_0930_),
    .A4(_0936_),
    .ZN(_0937_));
 AND4_X1 _3548_ (.A1(_2064_),
    .A2(_2055_),
    .A3(_2067_),
    .A4(_2070_),
    .ZN(_0938_));
 NAND2_X1 _3549_ (.A1(_2052_),
    .A2(_2058_),
    .ZN(_0939_));
 INV_X1 _3550_ (.A(_2049_),
    .ZN(_0940_));
 AOI21_X1 _3551_ (.A(_0939_),
    .B1(_0940_),
    .B2(_2048_),
    .ZN(_0941_));
 AOI21_X1 _3552_ (.A(_2057_),
    .B1(_2058_),
    .B2(_2051_),
    .ZN(_0942_));
 INV_X1 _3553_ (.A(_0942_),
    .ZN(_0943_));
 OAI211_X2 _3554_ (.A(_0937_),
    .B(_0938_),
    .C1(_0941_),
    .C2(_0943_),
    .ZN(_0944_));
 AOI21_X1 _3555_ (.A(_2099_),
    .B1(_2100_),
    .B2(_2102_),
    .ZN(_0945_));
 AOI21_X1 _3556_ (.A(_2105_),
    .B1(_2106_),
    .B2(_2072_),
    .ZN(_0946_));
 NAND2_X1 _3557_ (.A1(_2100_),
    .A2(_2103_),
    .ZN(_0947_));
 OAI21_X2 _3558_ (.A(_0945_),
    .B1(_0946_),
    .B2(_0947_),
    .ZN(_0948_));
 NOR4_X4 _3559_ (.A1(_0905_),
    .A2(_0907_),
    .A3(_0924_),
    .A4(_0948_),
    .ZN(_0949_));
 AOI21_X1 _3560_ (.A(_2087_),
    .B1(_2088_),
    .B2(_2090_),
    .ZN(_0950_));
 AOI21_X1 _3561_ (.A(_2093_),
    .B1(_2094_),
    .B2(_2060_),
    .ZN(_0951_));
 NAND2_X1 _3562_ (.A1(_2088_),
    .A2(_2091_),
    .ZN(_0952_));
 OAI21_X2 _3563_ (.A(_0950_),
    .B1(_0951_),
    .B2(_0952_),
    .ZN(_0953_));
 NOR3_X2 _3564_ (.A1(_0935_),
    .A2(_0927_),
    .A3(_0930_),
    .ZN(_0954_));
 AOI21_X1 _3565_ (.A(_2063_),
    .B1(_2066_),
    .B2(_2064_),
    .ZN(_0955_));
 AOI21_X1 _3566_ (.A(_2069_),
    .B1(_2070_),
    .B2(_2054_),
    .ZN(_0956_));
 NAND2_X1 _3567_ (.A1(_2064_),
    .A2(_2067_),
    .ZN(_0957_));
 OAI21_X2 _3568_ (.A(_0955_),
    .B1(_0956_),
    .B2(_0957_),
    .ZN(_0958_));
 AOI22_X4 _3569_ (.A1(_0953_),
    .A2(_0954_),
    .B1(_0958_),
    .B2(_0937_),
    .ZN(_0959_));
 NAND4_X4 _3570_ (.A1(_0934_),
    .A2(_0944_),
    .A3(_0949_),
    .A4(_0959_),
    .ZN(_0960_));
 NAND3_X4 _3571_ (.A1(_0915_),
    .A2(_0926_),
    .A3(_0960_),
    .ZN(_0961_));
 MUX2_X2 _3572_ (.A(_0897_),
    .B(_0901_),
    .S(_0961_),
    .Z(_0962_));
 XNOR2_X2 _3573_ (.A(_0893_),
    .B(_0962_),
    .ZN(_0963_));
 BUF_X4 _3574_ (.A(_0963_),
    .Z(_0964_));
 AOI21_X1 _3575_ (.A(_2041_),
    .B1(_2000_),
    .B2(_0894_),
    .ZN(_0965_));
 INV_X1 _3576_ (.A(_0965_),
    .ZN(_0966_));
 AOI21_X1 _3577_ (.A(_2035_),
    .B1(_0966_),
    .B2(_0892_),
    .ZN(_0967_));
 AOI21_X1 _3578_ (.A(_2038_),
    .B1(_1996_),
    .B2(_0894_),
    .ZN(_0968_));
 INV_X1 _3579_ (.A(_0968_),
    .ZN(_0969_));
 AOI21_X1 _3580_ (.A(_2032_),
    .B1(_0969_),
    .B2(_0892_),
    .ZN(_0970_));
 BUF_X8 _3581_ (.A(_0961_),
    .Z(_0971_));
 MUX2_X2 _3582_ (.A(_0967_),
    .B(_0970_),
    .S(_0971_),
    .Z(_0972_));
 XNOR2_X2 _3583_ (.A(_0903_),
    .B(_0972_),
    .ZN(_0973_));
 INV_X1 _3584_ (.A(_0894_),
    .ZN(_0974_));
 NOR2_X2 _3585_ (.A1(_0974_),
    .A2(_1996_),
    .ZN(_0975_));
 AND2_X1 _3586_ (.A1(_0974_),
    .A2(_1996_),
    .ZN(_0976_));
 OAI21_X4 _3587_ (.A(_0971_),
    .B1(_0975_),
    .B2(_0976_),
    .ZN(_0977_));
 NOR4_X4 _3588_ (.A1(_2011_),
    .A2(_0908_),
    .A3(_0913_),
    .A4(_0914_),
    .ZN(_0978_));
 OR2_X2 _3589_ (.A1(_0916_),
    .A2(_0925_),
    .ZN(_0979_));
 AND4_X2 _3590_ (.A1(_0934_),
    .A2(_0944_),
    .A3(_0949_),
    .A4(_0959_),
    .ZN(_0980_));
 NOR3_X4 _3591_ (.A1(_0978_),
    .A2(_0979_),
    .A3(_0980_),
    .ZN(_0981_));
 NOR2_X2 _3592_ (.A1(_0974_),
    .A2(_2000_),
    .ZN(_0982_));
 AND2_X1 _3593_ (.A1(_0974_),
    .A2(_2000_),
    .ZN(_0983_));
 OAI21_X4 _3594_ (.A(_0981_),
    .B1(_0982_),
    .B2(_0983_),
    .ZN(_0984_));
 NAND2_X4 _3595_ (.A1(_0977_),
    .A2(_0984_),
    .ZN(_0985_));
 BUF_X4 _3596_ (.A(_2118_),
    .Z(_0986_));
 BUF_X4 _3597_ (.A(_0986_),
    .Z(_0987_));
 BUF_X4 _3598_ (.A(_0987_),
    .Z(_0988_));
 INV_X1 _3599_ (.A(_2001_),
    .ZN(_0989_));
 NOR4_X4 _3600_ (.A1(_0989_),
    .A2(_0978_),
    .A3(_0979_),
    .A4(_0980_),
    .ZN(_0990_));
 BUF_X4 _3601_ (.A(_1997_),
    .Z(_0991_));
 AOI21_X4 _3602_ (.A(_0990_),
    .B1(_0971_),
    .B2(_0991_),
    .ZN(_0992_));
 NOR2_X1 _3603_ (.A1(_0988_),
    .A2(_0992_),
    .ZN(_0993_));
 OAI211_X4 _3604_ (.A(_0964_),
    .B(_0973_),
    .C1(_0985_),
    .C2(_0993_),
    .ZN(_0994_));
 BUF_X4 _3605_ (.A(_0971_),
    .Z(_0995_));
 NOR4_X1 _3606_ (.A1(net21),
    .A2(net20),
    .A3(net24),
    .A4(net22),
    .ZN(_0996_));
 NOR4_X2 _3607_ (.A1(net17),
    .A2(net16),
    .A3(net19),
    .A4(net18),
    .ZN(_0997_));
 NAND2_X2 _3608_ (.A1(_0996_),
    .A2(_0997_),
    .ZN(_0998_));
 NOR2_X4 _3609_ (.A1(_0409_),
    .A2(_0998_),
    .ZN(_0999_));
 NOR2_X2 _3610_ (.A1(_1585_),
    .A2(_0999_),
    .ZN(_1000_));
 NOR4_X2 _3611_ (.A1(net45),
    .A2(net44),
    .A3(net48),
    .A4(net46),
    .ZN(_1001_));
 NOR4_X2 _3612_ (.A1(net41),
    .A2(net40),
    .A3(net42),
    .A4(net43),
    .ZN(_1002_));
 NAND2_X2 _3613_ (.A1(_1001_),
    .A2(_1002_),
    .ZN(_1003_));
 NOR3_X4 _3614_ (.A1(_0425_),
    .A2(_0428_),
    .A3(_1003_),
    .ZN(_1004_));
 INV_X1 _3615_ (.A(_1004_),
    .ZN(_1005_));
 AOI21_X1 _3616_ (.A(_2020_),
    .B1(_2026_),
    .B2(_0904_),
    .ZN(_1006_));
 NAND2_X1 _3617_ (.A1(_0903_),
    .A2(_0904_),
    .ZN(_1007_));
 OAI21_X1 _3618_ (.A(_1006_),
    .B1(_1007_),
    .B2(_0970_),
    .ZN(_1008_));
 INV_X1 _3619_ (.A(_2020_),
    .ZN(_1009_));
 AOI21_X2 _3620_ (.A(_2026_),
    .B1(_2032_),
    .B2(_0903_),
    .ZN(_1010_));
 INV_X1 _3621_ (.A(_0904_),
    .ZN(_1011_));
 OAI21_X1 _3622_ (.A(_1009_),
    .B1(_1010_),
    .B2(_1011_),
    .ZN(_1012_));
 AOI21_X1 _3623_ (.A(_2014_),
    .B1(_1012_),
    .B2(_0902_),
    .ZN(_1013_));
 INV_X1 _3624_ (.A(_0902_),
    .ZN(_1014_));
 NAND2_X1 _3625_ (.A1(_0903_),
    .A2(_0892_),
    .ZN(_1015_));
 NOR3_X1 _3626_ (.A1(_1014_),
    .A2(_1011_),
    .A3(_1015_),
    .ZN(_1016_));
 OAI21_X1 _3627_ (.A(_1016_),
    .B1(_0898_),
    .B2(_0900_),
    .ZN(_1017_));
 NOR2_X1 _3628_ (.A1(_2008_),
    .A2(_2014_),
    .ZN(_1018_));
 NOR2_X1 _3629_ (.A1(_0906_),
    .A2(_1018_),
    .ZN(_1019_));
 AND3_X1 _3630_ (.A1(_1013_),
    .A2(_1017_),
    .A3(_1019_),
    .ZN(_1020_));
 INV_X1 _3631_ (.A(_0906_),
    .ZN(_1021_));
 AOI21_X1 _3632_ (.A(_1021_),
    .B1(_1013_),
    .B2(_1017_),
    .ZN(_1022_));
 OAI211_X2 _3633_ (.A(_0902_),
    .B(_1008_),
    .C1(_1020_),
    .C2(_1022_),
    .ZN(_1023_));
 OR3_X1 _3634_ (.A1(_0902_),
    .A2(_1018_),
    .A3(_1008_),
    .ZN(_1024_));
 NAND2_X1 _3635_ (.A1(_1013_),
    .A2(_1017_),
    .ZN(_1025_));
 XNOR2_X2 _3636_ (.A(_1021_),
    .B(_1025_),
    .ZN(_1026_));
 OAI211_X4 _3637_ (.A(_0971_),
    .B(_1023_),
    .C1(_1024_),
    .C2(_1026_),
    .ZN(_1027_));
 NAND4_X2 _3638_ (.A1(_0995_),
    .A2(_1000_),
    .A3(_1005_),
    .A4(_1027_),
    .ZN(_1028_));
 AND2_X1 _3639_ (.A1(_0895_),
    .A2(_0896_),
    .ZN(_1029_));
 INV_X1 _3640_ (.A(_0901_),
    .ZN(_1030_));
 MUX2_X1 _3641_ (.A(_1029_),
    .B(_1030_),
    .S(_0971_),
    .Z(_1031_));
 NOR2_X1 _3642_ (.A1(_2029_),
    .A2(_0910_),
    .ZN(_1032_));
 AND4_X1 _3643_ (.A1(_1032_),
    .A2(_0915_),
    .A3(_0926_),
    .A4(_0960_),
    .ZN(_1033_));
 AND2_X1 _3644_ (.A1(_0995_),
    .A2(_1010_),
    .ZN(_1034_));
 OAI221_X2 _3645_ (.A(_1011_),
    .B1(_1015_),
    .B2(_1031_),
    .C1(_1033_),
    .C2(_1034_),
    .ZN(_1035_));
 AOI21_X2 _3646_ (.A(_1033_),
    .B1(_1010_),
    .B2(_0995_),
    .ZN(_1036_));
 NOR2_X1 _3647_ (.A1(_1011_),
    .A2(_1015_),
    .ZN(_1037_));
 AOI22_X4 _3648_ (.A1(_0904_),
    .A2(_1036_),
    .B1(_1037_),
    .B2(_0962_),
    .ZN(_1038_));
 AOI21_X4 _3649_ (.A(_1028_),
    .B1(_1035_),
    .B2(_1038_),
    .ZN(_1039_));
 NAND2_X2 _3650_ (.A1(_0994_),
    .A2(_1039_),
    .ZN(_1040_));
 XNOR2_X2 _3651_ (.A(_0892_),
    .B(_0962_),
    .ZN(_1041_));
 NOR2_X1 _3652_ (.A1(_2029_),
    .A2(_2035_),
    .ZN(_1042_));
 OAI21_X1 _3653_ (.A(_1042_),
    .B1(_0965_),
    .B2(_0893_),
    .ZN(_1043_));
 OAI21_X1 _3654_ (.A(_0904_),
    .B1(_2029_),
    .B2(_0903_),
    .ZN(_1044_));
 INV_X1 _3655_ (.A(_1044_),
    .ZN(_1045_));
 AOI21_X2 _3656_ (.A(_2023_),
    .B1(_1043_),
    .B2(_1045_),
    .ZN(_1046_));
 OAI21_X1 _3657_ (.A(_0909_),
    .B1(_1046_),
    .B2(_1014_),
    .ZN(_1047_));
 AOI21_X2 _3658_ (.A(_2011_),
    .B1(_0906_),
    .B2(_1047_),
    .ZN(_1048_));
 XNOR2_X1 _3659_ (.A(_1014_),
    .B(_1046_),
    .ZN(_1049_));
 OAI21_X1 _3660_ (.A(_1021_),
    .B1(_0913_),
    .B2(_0914_),
    .ZN(_1050_));
 OR3_X1 _3661_ (.A1(_1021_),
    .A2(_0913_),
    .A3(_0914_),
    .ZN(_1051_));
 NAND3_X2 _3662_ (.A1(_1049_),
    .A2(_1050_),
    .A3(_1051_),
    .ZN(_1052_));
 OAI21_X4 _3663_ (.A(_0981_),
    .B1(_1048_),
    .B2(_1052_),
    .ZN(_1053_));
 NAND2_X2 _3664_ (.A1(_1027_),
    .A2(_1053_),
    .ZN(_1054_));
 BUF_X4 _3665_ (.A(_1054_),
    .Z(_1055_));
 NOR2_X2 _3666_ (.A1(_1041_),
    .A2(_1055_),
    .ZN(_1056_));
 INV_X4 _3667_ (.A(_0986_),
    .ZN(_1057_));
 BUF_X4 _3668_ (.A(_1057_),
    .Z(_1058_));
 CLKBUF_X3 _3669_ (.A(_1058_),
    .Z(_1059_));
 CLKBUF_X3 _3670_ (.A(_1059_),
    .Z(_1060_));
 INV_X1 _3671_ (.A(_0975_),
    .ZN(_1061_));
 INV_X1 _3672_ (.A(_0976_),
    .ZN(_1062_));
 AOI21_X4 _3673_ (.A(_0981_),
    .B1(_1061_),
    .B2(_1062_),
    .ZN(_1063_));
 INV_X1 _3674_ (.A(_0982_),
    .ZN(_1064_));
 INV_X1 _3675_ (.A(_0983_),
    .ZN(_1065_));
 AOI21_X4 _3676_ (.A(_0971_),
    .B1(_1064_),
    .B2(_1065_),
    .ZN(_1066_));
 NOR2_X4 _3677_ (.A1(_1063_),
    .A2(_1066_),
    .ZN(_1067_));
 NAND4_X4 _3678_ (.A1(_2001_),
    .A2(_0915_),
    .A3(_0926_),
    .A4(_0960_),
    .ZN(_1068_));
 INV_X2 _3679_ (.A(_0991_),
    .ZN(_1069_));
 OAI21_X4 _3680_ (.A(_1068_),
    .B1(_0981_),
    .B2(_1069_),
    .ZN(_1070_));
 BUF_X8 _3681_ (.A(_1070_),
    .Z(_1071_));
 MUX2_X1 _3682_ (.A(_0392_),
    .B(_0396_),
    .S(_1071_),
    .Z(_1072_));
 NOR3_X1 _3683_ (.A1(_1060_),
    .A2(_1067_),
    .A3(_1072_),
    .ZN(_1073_));
 BUF_X4 _3684_ (.A(_0987_),
    .Z(_1074_));
 BUF_X4 _3685_ (.A(_1074_),
    .Z(_1075_));
 BUF_X4 _3686_ (.A(_1070_),
    .Z(_1076_));
 MUX2_X1 _3687_ (.A(_0405_),
    .B(_0395_),
    .S(_1076_),
    .Z(_1077_));
 NOR3_X1 _3688_ (.A1(_1075_),
    .A2(_1067_),
    .A3(_1077_),
    .ZN(_1078_));
 BUF_X4 _3689_ (.A(_1058_),
    .Z(_1079_));
 BUF_X4 _3690_ (.A(_1070_),
    .Z(_1080_));
 MUX2_X1 _3691_ (.A(net29),
    .B(_0402_),
    .S(_1080_),
    .Z(_1081_));
 NOR3_X1 _3692_ (.A1(_1079_),
    .A2(_0985_),
    .A3(_1081_),
    .ZN(_1082_));
 MUX2_X1 _3693_ (.A(_0404_),
    .B(_0401_),
    .S(_1080_),
    .Z(_1083_));
 NOR3_X1 _3694_ (.A1(_1075_),
    .A2(_0985_),
    .A3(_1083_),
    .ZN(_1084_));
 NOR4_X2 _3695_ (.A1(_1073_),
    .A2(_1078_),
    .A3(_1082_),
    .A4(_1084_),
    .ZN(_1085_));
 NAND2_X1 _3696_ (.A1(_1056_),
    .A2(_1085_),
    .ZN(_1086_));
 BUF_X4 _3697_ (.A(_0973_),
    .Z(_1087_));
 NOR2_X4 _3698_ (.A1(_0963_),
    .A2(_1055_),
    .ZN(_1088_));
 MUX2_X1 _3699_ (.A(net23),
    .B(_0400_),
    .S(_1071_),
    .Z(_1089_));
 MUX2_X1 _3700_ (.A(net26),
    .B(net28),
    .S(_1071_),
    .Z(_1090_));
 MUX2_X1 _3701_ (.A(_1089_),
    .B(_1090_),
    .S(_1058_),
    .Z(_1091_));
 CLKBUF_X3 _3702_ (.A(_0992_),
    .Z(_1092_));
 CLKBUF_X3 _3703_ (.A(_1092_),
    .Z(_1093_));
 INV_X1 _3704_ (.A(net12),
    .ZN(_1094_));
 MUX2_X1 _3705_ (.A(_1094_),
    .B(_2047_),
    .S(_1074_),
    .Z(_1095_));
 NOR2_X1 _3706_ (.A1(_1093_),
    .A2(_1095_),
    .ZN(_1096_));
 BUF_X4 _3707_ (.A(_1067_),
    .Z(_1097_));
 MUX2_X1 _3708_ (.A(_1091_),
    .B(_1096_),
    .S(_1097_),
    .Z(_1098_));
 AOI21_X1 _3709_ (.A(_1087_),
    .B1(_1088_),
    .B2(_1098_),
    .ZN(_1099_));
 AND2_X2 _3710_ (.A1(_1027_),
    .A2(_1053_),
    .ZN(_1100_));
 MUX2_X1 _3711_ (.A(net11),
    .B(net10),
    .S(_0986_),
    .Z(_1101_));
 MUX2_X1 _3712_ (.A(net14),
    .B(_0390_),
    .S(_0986_),
    .Z(_1102_));
 MUX2_X1 _3713_ (.A(_1101_),
    .B(_1102_),
    .S(_1080_),
    .Z(_1103_));
 AND4_X1 _3714_ (.A1(_1041_),
    .A2(_0985_),
    .A3(_1100_),
    .A4(_1103_),
    .ZN(_1104_));
 BUF_X4 _3715_ (.A(_0985_),
    .Z(_1105_));
 NOR2_X1 _3716_ (.A1(_0964_),
    .A2(_1105_),
    .ZN(_1106_));
 MUX2_X1 _3717_ (.A(net9),
    .B(_0389_),
    .S(_0986_),
    .Z(_1107_));
 NAND2_X1 _3718_ (.A1(_0393_),
    .A2(_0987_),
    .ZN(_1108_));
 NAND2_X1 _3719_ (.A1(_0397_),
    .A2(_1057_),
    .ZN(_1109_));
 NAND2_X1 _3720_ (.A1(_1108_),
    .A2(_1109_),
    .ZN(_1110_));
 MUX2_X1 _3721_ (.A(_1107_),
    .B(_1110_),
    .S(_0992_),
    .Z(_1111_));
 AND2_X1 _3722_ (.A1(_1100_),
    .A2(_1111_),
    .ZN(_1112_));
 MUX2_X1 _3723_ (.A(net15),
    .B(_0998_),
    .S(_1057_),
    .Z(_1113_));
 NAND2_X1 _3724_ (.A1(_1092_),
    .A2(_1113_),
    .ZN(_1114_));
 NOR3_X4 _3725_ (.A1(_1105_),
    .A2(_1055_),
    .A3(_1114_),
    .ZN(_1115_));
 AOI221_X2 _3726_ (.A(_1104_),
    .B1(_1106_),
    .B2(_1112_),
    .C1(_1115_),
    .C2(_0964_),
    .ZN(_1116_));
 AOI221_X2 _3727_ (.A(_1040_),
    .B1(_1086_),
    .B2(_1099_),
    .C1(_1116_),
    .C2(_1087_),
    .ZN(_0113_));
 INV_X1 _3728_ (.A(_0999_),
    .ZN(_1117_));
 NAND2_X4 _3729_ (.A1(_1740_),
    .A2(_1117_),
    .ZN(_1118_));
 NOR2_X1 _3730_ (.A1(_0981_),
    .A2(_1004_),
    .ZN(_1119_));
 NOR2_X1 _3731_ (.A1(_1118_),
    .A2(_1119_),
    .ZN(_1120_));
 CLKBUF_X3 _3732_ (.A(_1120_),
    .Z(_1121_));
 NAND2_X1 _3733_ (.A1(_0402_),
    .A2(_1121_),
    .ZN(_1122_));
 XOR2_X2 _3734_ (.A(_0903_),
    .B(_0972_),
    .Z(_1123_));
 BUF_X4 _3735_ (.A(_1123_),
    .Z(_1124_));
 NAND2_X2 _3736_ (.A1(_1124_),
    .A2(_1039_),
    .ZN(_1125_));
 AND4_X1 _3737_ (.A1(_0977_),
    .A2(_0984_),
    .A3(_1027_),
    .A4(_1053_),
    .ZN(_1126_));
 BUF_X4 _3738_ (.A(_1126_),
    .Z(_1127_));
 NAND2_X1 _3739_ (.A1(_0405_),
    .A2(_1059_),
    .ZN(_1128_));
 NAND2_X1 _3740_ (.A1(_0392_),
    .A2(_0988_),
    .ZN(_1129_));
 AOI21_X1 _3741_ (.A(_1092_),
    .B1(_1128_),
    .B2(_1129_),
    .ZN(_1130_));
 BUF_X8 _3742_ (.A(_1071_),
    .Z(_1131_));
 BUF_X4 _3743_ (.A(_1131_),
    .Z(_1132_));
 NAND2_X1 _3744_ (.A1(_0401_),
    .A2(_1059_),
    .ZN(_1133_));
 NAND2_X1 _3745_ (.A1(_0402_),
    .A2(_0988_),
    .ZN(_1134_));
 AOI21_X1 _3746_ (.A(_1132_),
    .B1(_1133_),
    .B2(_1134_),
    .ZN(_1135_));
 OAI21_X1 _3747_ (.A(_1127_),
    .B1(_1130_),
    .B2(_1135_),
    .ZN(_1136_));
 CLKBUF_X3 _3748_ (.A(_1100_),
    .Z(_1137_));
 AOI21_X2 _3749_ (.A(_1092_),
    .B1(_1108_),
    .B2(_1109_),
    .ZN(_1138_));
 BUF_X4 _3750_ (.A(_1076_),
    .Z(_1139_));
 NAND2_X1 _3751_ (.A1(_0395_),
    .A2(_1058_),
    .ZN(_1140_));
 NAND2_X1 _3752_ (.A1(_0396_),
    .A2(_0988_),
    .ZN(_1141_));
 AOI21_X2 _3753_ (.A(_1139_),
    .B1(_1140_),
    .B2(_1141_),
    .ZN(_1142_));
 OAI221_X2 _3754_ (.A(_1137_),
    .B1(_1138_),
    .B2(_1142_),
    .C1(_1066_),
    .C2(_1063_),
    .ZN(_1143_));
 AND2_X1 _3755_ (.A1(_1136_),
    .A2(_1143_),
    .ZN(_1144_));
 MUX2_X1 _3756_ (.A(_1113_),
    .B(_1102_),
    .S(_0992_),
    .Z(_1145_));
 MUX2_X1 _3757_ (.A(_1101_),
    .B(_1107_),
    .S(_0992_),
    .Z(_1146_));
 MUX2_X1 _3758_ (.A(_1145_),
    .B(_1146_),
    .S(_1097_),
    .Z(_1147_));
 NAND2_X1 _3759_ (.A1(_1137_),
    .A2(_1147_),
    .ZN(_1148_));
 BUF_X4 _3760_ (.A(_0964_),
    .Z(_1149_));
 MUX2_X1 _3761_ (.A(_1144_),
    .B(_1148_),
    .S(_1149_),
    .Z(_1150_));
 OAI21_X1 _3762_ (.A(_1122_),
    .B1(_1125_),
    .B2(_1150_),
    .ZN(_0114_));
 INV_X1 _3763_ (.A(_0401_),
    .ZN(_1151_));
 CLKBUF_X3 _3764_ (.A(_1119_),
    .Z(_1152_));
 CLKBUF_X3 _3765_ (.A(_1041_),
    .Z(_1153_));
 BUF_X4 _3766_ (.A(_1127_),
    .Z(_1154_));
 MUX2_X1 _3767_ (.A(_0401_),
    .B(_0405_),
    .S(_1071_),
    .Z(_1155_));
 MUX2_X1 _3768_ (.A(_1072_),
    .B(_1155_),
    .S(_1074_),
    .Z(_1156_));
 MUX2_X1 _3769_ (.A(_0395_),
    .B(_0397_),
    .S(_1131_),
    .Z(_1157_));
 MUX2_X1 _3770_ (.A(_0393_),
    .B(_0389_),
    .S(_1131_),
    .Z(_1158_));
 MUX2_X1 _3771_ (.A(_1157_),
    .B(_1158_),
    .S(_1059_),
    .Z(_1159_));
 NOR2_X4 _3772_ (.A1(_1067_),
    .A2(_1054_),
    .ZN(_1160_));
 AOI22_X2 _3773_ (.A1(_1154_),
    .A2(_1156_),
    .B1(_1159_),
    .B2(_1160_),
    .ZN(_1161_));
 AND2_X1 _3774_ (.A1(_1153_),
    .A2(_1161_),
    .ZN(_1162_));
 NAND4_X4 _3775_ (.A1(_0977_),
    .A2(_0984_),
    .A3(_1027_),
    .A4(_1053_),
    .ZN(_1163_));
 AND2_X1 _3776_ (.A1(_0390_),
    .A2(_1058_),
    .ZN(_1164_));
 NAND2_X1 _3777_ (.A1(net11),
    .A2(_1074_),
    .ZN(_1165_));
 INV_X1 _3778_ (.A(_1165_),
    .ZN(_1166_));
 OAI21_X1 _3779_ (.A(_1132_),
    .B1(_1164_),
    .B2(_1166_),
    .ZN(_1167_));
 AND2_X1 _3780_ (.A1(net10),
    .A2(_1058_),
    .ZN(_1168_));
 AND2_X1 _3781_ (.A1(net9),
    .A2(_1074_),
    .ZN(_1169_));
 OAI21_X1 _3782_ (.A(_1092_),
    .B1(_1168_),
    .B2(_1169_),
    .ZN(_1170_));
 AND2_X1 _3783_ (.A1(_1167_),
    .A2(_1170_),
    .ZN(_1171_));
 NAND2_X1 _3784_ (.A1(net14),
    .A2(_0987_),
    .ZN(_1172_));
 NAND2_X1 _3785_ (.A1(net15),
    .A2(_1057_),
    .ZN(_1173_));
 AOI221_X2 _3786_ (.A(_0990_),
    .B1(_1172_),
    .B2(_1173_),
    .C1(_0995_),
    .C2(_0991_),
    .ZN(_1174_));
 NAND2_X1 _3787_ (.A1(_1074_),
    .A2(_0998_),
    .ZN(_1175_));
 INV_X1 _3788_ (.A(_1175_),
    .ZN(_1176_));
 AOI21_X4 _3789_ (.A(_1174_),
    .B1(_1176_),
    .B2(_1132_),
    .ZN(_1177_));
 OAI211_X4 _3790_ (.A(_1027_),
    .B(_1053_),
    .C1(_1063_),
    .C2(_1066_),
    .ZN(_1178_));
 OAI22_X4 _3791_ (.A1(_1163_),
    .A2(_1171_),
    .B1(_1177_),
    .B2(_1178_),
    .ZN(_1179_));
 NOR2_X1 _3792_ (.A1(_1153_),
    .A2(_1179_),
    .ZN(_1180_));
 OAI33_X1 _3793_ (.A1(_1151_),
    .A2(_1118_),
    .A3(_1152_),
    .B1(_1125_),
    .B2(_1162_),
    .B3(_1180_),
    .ZN(_0115_));
 NAND2_X1 _3794_ (.A1(_0392_),
    .A2(_1121_),
    .ZN(_1181_));
 CLKBUF_X3 _3795_ (.A(_1105_),
    .Z(_1182_));
 MUX2_X1 _3796_ (.A(_1072_),
    .B(_1077_),
    .S(_1060_),
    .Z(_1183_));
 AOI22_X2 _3797_ (.A1(_1182_),
    .A2(_1112_),
    .B1(_1183_),
    .B2(_1154_),
    .ZN(_1184_));
 AND2_X2 _3798_ (.A1(_1123_),
    .A2(_1039_),
    .ZN(_1185_));
 NAND2_X2 _3799_ (.A1(_1153_),
    .A2(_1185_),
    .ZN(_1186_));
 NOR2_X2 _3800_ (.A1(_1041_),
    .A2(_1087_),
    .ZN(_1187_));
 NAND2_X1 _3801_ (.A1(_1039_),
    .A2(_1187_),
    .ZN(_1188_));
 CLKBUF_X3 _3802_ (.A(_1097_),
    .Z(_1189_));
 NAND2_X1 _3803_ (.A1(_1189_),
    .A2(_1103_),
    .ZN(_1190_));
 OR2_X1 _3804_ (.A1(_1189_),
    .A2(_1114_),
    .ZN(_1191_));
 AOI21_X2 _3805_ (.A(_1055_),
    .B1(_1190_),
    .B2(_1191_),
    .ZN(_1192_));
 INV_X1 _3806_ (.A(_1192_),
    .ZN(_1193_));
 OAI221_X1 _3807_ (.A(_1181_),
    .B1(_1184_),
    .B2(_1186_),
    .C1(_1188_),
    .C2(_1193_),
    .ZN(_0116_));
 NAND2_X1 _3808_ (.A1(_0405_),
    .A2(_1121_),
    .ZN(_1194_));
 MUX2_X1 _3809_ (.A(_0396_),
    .B(_0393_),
    .S(_1139_),
    .Z(_1195_));
 MUX2_X1 _3810_ (.A(_1077_),
    .B(_1195_),
    .S(_1060_),
    .Z(_1196_));
 NAND3_X1 _3811_ (.A1(_0397_),
    .A2(_1075_),
    .A3(_1093_),
    .ZN(_1197_));
 NAND3_X1 _3812_ (.A1(_0389_),
    .A2(_1079_),
    .A3(_1093_),
    .ZN(_1198_));
 OAI21_X1 _3813_ (.A(_1132_),
    .B1(_1168_),
    .B2(_1169_),
    .ZN(_1199_));
 NAND3_X1 _3814_ (.A1(_1197_),
    .A2(_1198_),
    .A3(_1199_),
    .ZN(_1200_));
 AOI22_X2 _3815_ (.A1(_1154_),
    .A2(_1196_),
    .B1(_1200_),
    .B2(_1160_),
    .ZN(_1201_));
 AOI21_X1 _3816_ (.A(_1092_),
    .B1(_1172_),
    .B2(_1173_),
    .ZN(_1202_));
 NAND2_X1 _3817_ (.A1(_0390_),
    .A2(_1058_),
    .ZN(_1203_));
 AOI21_X1 _3818_ (.A(_1139_),
    .B1(_1203_),
    .B2(_1165_),
    .ZN(_1204_));
 OAI21_X1 _3819_ (.A(_1189_),
    .B1(_1202_),
    .B2(_1204_),
    .ZN(_1205_));
 NAND3_X1 _3820_ (.A1(_1182_),
    .A2(_1093_),
    .A3(_1176_),
    .ZN(_1206_));
 NAND2_X1 _3821_ (.A1(_1205_),
    .A2(_1206_),
    .ZN(_1207_));
 NAND2_X1 _3822_ (.A1(_1185_),
    .A2(_1207_),
    .ZN(_1208_));
 NAND2_X1 _3823_ (.A1(_1149_),
    .A2(_1137_),
    .ZN(_1209_));
 OAI221_X1 _3824_ (.A(_1194_),
    .B1(_1201_),
    .B2(_1186_),
    .C1(_1208_),
    .C2(_1209_),
    .ZN(_0117_));
 NAND2_X1 _3825_ (.A1(_0396_),
    .A2(_1121_),
    .ZN(_1210_));
 AND2_X1 _3826_ (.A1(_1154_),
    .A2(_1145_),
    .ZN(_1211_));
 NAND2_X1 _3827_ (.A1(_1182_),
    .A2(_1146_),
    .ZN(_1212_));
 NOR2_X1 _3828_ (.A1(_1138_),
    .A2(_1142_),
    .ZN(_1213_));
 OAI21_X1 _3829_ (.A(_1212_),
    .B1(_1213_),
    .B2(_1182_),
    .ZN(_1214_));
 CLKBUF_X3 _3830_ (.A(_1088_),
    .Z(_1215_));
 AOI22_X1 _3831_ (.A1(_1149_),
    .A2(_1211_),
    .B1(_1214_),
    .B2(_1215_),
    .ZN(_1216_));
 OAI21_X1 _3832_ (.A(_1210_),
    .B1(_1216_),
    .B2(_1125_),
    .ZN(_0118_));
 NAND2_X1 _3833_ (.A1(_0395_),
    .A2(_1121_),
    .ZN(_1217_));
 NOR2_X2 _3834_ (.A1(_1163_),
    .A2(_1177_),
    .ZN(_1218_));
 NAND2_X1 _3835_ (.A1(_1167_),
    .A2(_1170_),
    .ZN(_1219_));
 MUX2_X1 _3836_ (.A(_1159_),
    .B(_1219_),
    .S(_1182_),
    .Z(_1220_));
 AOI22_X1 _3837_ (.A1(_1149_),
    .A2(_1218_),
    .B1(_1220_),
    .B2(_1215_),
    .ZN(_1221_));
 OAI21_X1 _3838_ (.A(_1217_),
    .B1(_1221_),
    .B2(_1125_),
    .ZN(_0119_));
 NAND2_X1 _3839_ (.A1(_0995_),
    .A2(_1005_),
    .ZN(_1222_));
 CLKBUF_X3 _3840_ (.A(_1222_),
    .Z(_1223_));
 NAND2_X1 _3841_ (.A1(_0393_),
    .A2(_1223_),
    .ZN(_1224_));
 AOI21_X4 _3842_ (.A(_1055_),
    .B1(_1038_),
    .B2(_1035_),
    .ZN(_1225_));
 NAND3_X1 _3843_ (.A1(_1124_),
    .A2(_1152_),
    .A3(_1225_),
    .ZN(_1226_));
 OAI21_X1 _3844_ (.A(_1224_),
    .B1(_1226_),
    .B2(_1116_),
    .ZN(_1227_));
 AND2_X1 _3845_ (.A1(_1000_),
    .A2(_1227_),
    .ZN(_0120_));
 NAND2_X1 _3846_ (.A1(_0397_),
    .A2(_1121_),
    .ZN(_1228_));
 NOR4_X2 _3847_ (.A1(_1041_),
    .A2(_1132_),
    .A3(_1163_),
    .A4(_1175_),
    .ZN(_1229_));
 OR2_X1 _3848_ (.A1(_1202_),
    .A2(_1204_),
    .ZN(_1230_));
 MUX2_X1 _3849_ (.A(_1200_),
    .B(_1230_),
    .S(_1105_),
    .Z(_1231_));
 AOI21_X1 _3850_ (.A(_1229_),
    .B1(_1231_),
    .B2(_1215_),
    .ZN(_1232_));
 OAI21_X1 _3851_ (.A(_1228_),
    .B1(_1232_),
    .B2(_1125_),
    .ZN(_0121_));
 NAND2_X1 _3852_ (.A1(_0389_),
    .A2(_1223_),
    .ZN(_1233_));
 NOR2_X4 _3853_ (.A1(_0964_),
    .A2(_0973_),
    .ZN(_1234_));
 NAND2_X1 _3854_ (.A1(_1225_),
    .A2(_1234_),
    .ZN(_1235_));
 OR3_X1 _3855_ (.A1(_1222_),
    .A2(_1148_),
    .A3(_1235_),
    .ZN(_1236_));
 AOI21_X1 _3856_ (.A(_1118_),
    .B1(_1233_),
    .B2(_1236_),
    .ZN(_0122_));
 NAND2_X1 _3857_ (.A1(net9),
    .A2(_1223_),
    .ZN(_1237_));
 AND2_X1 _3858_ (.A1(_1225_),
    .A2(_1234_),
    .ZN(_1238_));
 NAND3_X1 _3859_ (.A1(_1152_),
    .A2(_1179_),
    .A3(_1238_),
    .ZN(_1239_));
 AOI21_X1 _3860_ (.A(_1118_),
    .B1(_1237_),
    .B2(_1239_),
    .ZN(_0123_));
 MUX2_X1 _3861_ (.A(_0402_),
    .B(_0392_),
    .S(_1139_),
    .Z(_1240_));
 MUX2_X1 _3862_ (.A(_1083_),
    .B(_1240_),
    .S(_1060_),
    .Z(_1241_));
 AOI22_X1 _3863_ (.A1(_1160_),
    .A2(_1196_),
    .B1(_1241_),
    .B2(_1154_),
    .ZN(_1242_));
 AND2_X1 _3864_ (.A1(_1187_),
    .A2(_1242_),
    .ZN(_1243_));
 OR2_X1 _3865_ (.A1(_1124_),
    .A2(_1229_),
    .ZN(_1244_));
 AOI21_X1 _3866_ (.A(_1244_),
    .B1(_1231_),
    .B2(_1215_),
    .ZN(_1245_));
 AND2_X1 _3867_ (.A1(_0994_),
    .A2(_1039_),
    .ZN(_1246_));
 NAND2_X2 _3868_ (.A1(_1041_),
    .A2(_1123_),
    .ZN(_1247_));
 NOR2_X1 _3869_ (.A1(_2047_),
    .A2(_1139_),
    .ZN(_1248_));
 AND2_X1 _3870_ (.A1(net23),
    .A2(_1139_),
    .ZN(_1249_));
 OAI21_X1 _3871_ (.A(_1079_),
    .B1(_1248_),
    .B2(_1249_),
    .ZN(_1250_));
 NOR2_X1 _3872_ (.A1(_1094_),
    .A2(_1059_),
    .ZN(_1251_));
 AOI21_X1 _3873_ (.A(_1105_),
    .B1(_1132_),
    .B2(_1251_),
    .ZN(_1252_));
 OAI211_X2 _3874_ (.A(_0400_),
    .B(_1068_),
    .C1(_0981_),
    .C2(_1069_),
    .ZN(_1253_));
 INV_X1 _3875_ (.A(net29),
    .ZN(_1254_));
 OAI211_X2 _3876_ (.A(_1079_),
    .B(_1253_),
    .C1(_1092_),
    .C2(_1254_),
    .ZN(_1255_));
 OAI21_X1 _3877_ (.A(_1255_),
    .B1(_1090_),
    .B2(_1079_),
    .ZN(_1256_));
 AOI221_X2 _3878_ (.A(_1055_),
    .B1(_1250_),
    .B2(_1252_),
    .C1(_1256_),
    .C2(_1105_),
    .ZN(_1257_));
 OAI21_X1 _3879_ (.A(_1246_),
    .B1(_1247_),
    .B2(_1257_),
    .ZN(_1258_));
 NOR3_X1 _3880_ (.A1(_1243_),
    .A2(_1245_),
    .A3(_1258_),
    .ZN(_0124_));
 NAND2_X1 _3881_ (.A1(net10),
    .A2(_1223_),
    .ZN(_1259_));
 NAND3_X1 _3882_ (.A1(_1152_),
    .A2(_1192_),
    .A3(_1238_),
    .ZN(_1260_));
 AOI21_X1 _3883_ (.A(_1118_),
    .B1(_1259_),
    .B2(_1260_),
    .ZN(_0125_));
 NAND2_X1 _3884_ (.A1(net11),
    .A2(_1223_),
    .ZN(_1261_));
 AOI21_X2 _3885_ (.A(_1055_),
    .B1(_1205_),
    .B2(_1206_),
    .ZN(_1262_));
 NAND3_X1 _3886_ (.A1(_1152_),
    .A2(_1238_),
    .A3(_1262_),
    .ZN(_1263_));
 AOI21_X1 _3887_ (.A(_1118_),
    .B1(_1261_),
    .B2(_1263_),
    .ZN(_0126_));
 NAND2_X1 _3888_ (.A1(_0390_),
    .A2(_1223_),
    .ZN(_1264_));
 NAND3_X1 _3889_ (.A1(_1152_),
    .A2(_1211_),
    .A3(_1238_),
    .ZN(_1265_));
 AOI21_X1 _3890_ (.A(_1118_),
    .B1(_1264_),
    .B2(_1265_),
    .ZN(_0127_));
 NAND2_X1 _3891_ (.A1(net14),
    .A2(_1223_),
    .ZN(_1266_));
 NAND3_X1 _3892_ (.A1(_1152_),
    .A2(_1218_),
    .A3(_1238_),
    .ZN(_1267_));
 AOI21_X1 _3893_ (.A(_1118_),
    .B1(_1266_),
    .B2(_1267_),
    .ZN(_0128_));
 NAND2_X1 _3894_ (.A1(net15),
    .A2(_1223_),
    .ZN(_1268_));
 NAND3_X1 _3895_ (.A1(_1152_),
    .A2(_1115_),
    .A3(_1238_),
    .ZN(_1269_));
 AOI21_X1 _3896_ (.A(_1118_),
    .B1(_1268_),
    .B2(_1269_),
    .ZN(_0129_));
 NAND3_X1 _3897_ (.A1(_1075_),
    .A2(_1093_),
    .A3(_1154_),
    .ZN(_1270_));
 OAI21_X1 _3898_ (.A(_1152_),
    .B1(_1235_),
    .B2(_1270_),
    .ZN(_1271_));
 AND3_X1 _3899_ (.A1(_1750_),
    .A2(_0998_),
    .A3(_1271_),
    .ZN(_0130_));
 NAND2_X1 _3900_ (.A1(net1),
    .A2(_1121_),
    .ZN(_1272_));
 NAND2_X1 _3901_ (.A1(_0964_),
    .A2(_1123_),
    .ZN(_1273_));
 AOI21_X1 _3902_ (.A(_1273_),
    .B1(_1143_),
    .B2(_1136_),
    .ZN(_1274_));
 NOR2_X4 _3903_ (.A1(_0964_),
    .A2(_1123_),
    .ZN(_1275_));
 AND3_X1 _3904_ (.A1(_1137_),
    .A2(_1147_),
    .A3(_1275_),
    .ZN(_1276_));
 OAI21_X1 _3905_ (.A(_1246_),
    .B1(_1274_),
    .B2(_1276_),
    .ZN(_1277_));
 NOR3_X1 _3906_ (.A1(_1060_),
    .A2(_1248_),
    .A3(_1249_),
    .ZN(_1278_));
 NOR2_X1 _3907_ (.A1(_1094_),
    .A2(_1132_),
    .ZN(_1279_));
 AND2_X1 _3908_ (.A1(net26),
    .A2(_1132_),
    .ZN(_1280_));
 NOR3_X1 _3909_ (.A1(_1075_),
    .A2(_1279_),
    .A3(_1280_),
    .ZN(_1281_));
 INV_X1 _3910_ (.A(_0400_),
    .ZN(_1282_));
 AOI211_X2 _3911_ (.A(_1282_),
    .B(_0990_),
    .C1(_0995_),
    .C2(_0991_),
    .ZN(_1283_));
 AOI211_X2 _3912_ (.A(_1058_),
    .B(_1283_),
    .C1(_1139_),
    .C2(net29),
    .ZN(_1284_));
 INV_X1 _3913_ (.A(net28),
    .ZN(_1285_));
 AOI211_X2 _3914_ (.A(_1285_),
    .B(_0990_),
    .C1(_0995_),
    .C2(_0991_),
    .ZN(_1286_));
 AOI211_X2 _3915_ (.A(_0988_),
    .B(_1286_),
    .C1(_1139_),
    .C2(_0404_),
    .ZN(_1287_));
 OAI33_X1 _3916_ (.A1(_1163_),
    .A2(_1278_),
    .A3(_1281_),
    .B1(_1284_),
    .B2(_1287_),
    .B3(_1178_),
    .ZN(_1288_));
 NAND3_X1 _3917_ (.A1(_1246_),
    .A2(_1234_),
    .A3(_1288_),
    .ZN(_1289_));
 NAND3_X1 _3918_ (.A1(_1272_),
    .A2(_1277_),
    .A3(_1289_),
    .ZN(_0131_));
 AND2_X1 _3919_ (.A1(_1039_),
    .A2(_1275_),
    .ZN(_1290_));
 AOI22_X1 _3920_ (.A1(net12),
    .A2(_1121_),
    .B1(_1179_),
    .B2(_1290_),
    .ZN(_1291_));
 NOR2_X1 _3921_ (.A1(_1075_),
    .A2(_1089_),
    .ZN(_1292_));
 NOR3_X1 _3922_ (.A1(_1060_),
    .A2(_1279_),
    .A3(_1280_),
    .ZN(_1293_));
 NOR3_X1 _3923_ (.A1(_1182_),
    .A2(_1292_),
    .A3(_1293_),
    .ZN(_1294_));
 MUX2_X1 _3924_ (.A(net28),
    .B(_0404_),
    .S(_1080_),
    .Z(_1295_));
 MUX2_X1 _3925_ (.A(_1081_),
    .B(_1295_),
    .S(_0988_),
    .Z(_1296_));
 AOI21_X1 _3926_ (.A(_1294_),
    .B1(_1296_),
    .B2(_1182_),
    .ZN(_1297_));
 OAI221_X1 _3927_ (.A(_1291_),
    .B1(_1297_),
    .B2(_1186_),
    .C1(_1188_),
    .C2(_1161_),
    .ZN(_0132_));
 AOI22_X1 _3928_ (.A1(net23),
    .A2(_1121_),
    .B1(_1192_),
    .B2(_1290_),
    .ZN(_1298_));
 OR2_X1 _3929_ (.A1(_1184_),
    .A2(_1188_),
    .ZN(_1299_));
 MUX2_X1 _3930_ (.A(_1081_),
    .B(_1083_),
    .S(_1060_),
    .Z(_1300_));
 MUX2_X1 _3931_ (.A(_1091_),
    .B(_1300_),
    .S(_1182_),
    .Z(_1301_));
 NAND3_X1 _3932_ (.A1(_1215_),
    .A2(_1185_),
    .A3(_1301_),
    .ZN(_1302_));
 NAND3_X1 _3933_ (.A1(_1298_),
    .A2(_1299_),
    .A3(_1302_),
    .ZN(_0133_));
 AOI22_X1 _3934_ (.A1(net26),
    .A2(_1121_),
    .B1(_1262_),
    .B2(_1290_),
    .ZN(_1303_));
 NOR2_X1 _3935_ (.A1(_1182_),
    .A2(_1256_),
    .ZN(_1304_));
 AOI21_X1 _3936_ (.A(_1304_),
    .B1(_1241_),
    .B2(_1182_),
    .ZN(_1305_));
 OAI221_X1 _3937_ (.A(_1303_),
    .B1(_1305_),
    .B2(_1186_),
    .C1(_1188_),
    .C2(_1201_),
    .ZN(_0134_));
 NAND3_X1 _3938_ (.A1(_1153_),
    .A2(_1154_),
    .A3(_1145_),
    .ZN(_1306_));
 NAND2_X1 _3939_ (.A1(_1087_),
    .A2(_1306_),
    .ZN(_1307_));
 AOI22_X1 _3940_ (.A1(_0400_),
    .A2(_1120_),
    .B1(_1307_),
    .B2(_1039_),
    .ZN(_1308_));
 AOI21_X1 _3941_ (.A(_1087_),
    .B1(_1223_),
    .B2(_0400_),
    .ZN(_1309_));
 OR2_X1 _3942_ (.A1(_1130_),
    .A2(_1135_),
    .ZN(_1310_));
 NOR2_X1 _3943_ (.A1(_1284_),
    .A2(_1287_),
    .ZN(_1311_));
 MUX2_X1 _3944_ (.A(_1310_),
    .B(_1311_),
    .S(_1189_),
    .Z(_1312_));
 AOI22_X1 _3945_ (.A1(_1056_),
    .A2(_1214_),
    .B1(_1312_),
    .B2(_1215_),
    .ZN(_1313_));
 AOI21_X1 _3946_ (.A(_1308_),
    .B1(_1309_),
    .B2(_1313_),
    .ZN(_0135_));
 NOR2_X2 _3947_ (.A1(_1055_),
    .A2(_1273_),
    .ZN(_1314_));
 NAND3_X1 _3948_ (.A1(_1246_),
    .A2(_1220_),
    .A3(_1314_),
    .ZN(_1315_));
 AOI221_X1 _3949_ (.A(_1087_),
    .B1(_1160_),
    .B2(_1156_),
    .C1(_1296_),
    .C2(_1127_),
    .ZN(_1316_));
 OAI21_X1 _3950_ (.A(_1041_),
    .B1(_1124_),
    .B2(_1218_),
    .ZN(_1317_));
 OR2_X1 _3951_ (.A1(_1316_),
    .A2(_1317_),
    .ZN(_1318_));
 NAND2_X1 _3952_ (.A1(_1000_),
    .A2(_1223_),
    .ZN(_1319_));
 OAI221_X2 _3953_ (.A(_1315_),
    .B1(_1318_),
    .B2(_1040_),
    .C1(_1285_),
    .C2(_1319_),
    .ZN(_0136_));
 NAND3_X1 _3954_ (.A1(_1153_),
    .A2(_1085_),
    .A3(_1185_),
    .ZN(_1320_));
 NAND3_X1 _3955_ (.A1(_1189_),
    .A2(_1137_),
    .A3(_1111_),
    .ZN(_1321_));
 INV_X1 _3956_ (.A(_1103_),
    .ZN(_1322_));
 OAI21_X1 _3957_ (.A(_1321_),
    .B1(_1178_),
    .B2(_1322_),
    .ZN(_1323_));
 AOI22_X2 _3958_ (.A1(_1323_),
    .A2(_1187_),
    .B1(_1275_),
    .B2(_1115_),
    .ZN(_1324_));
 OAI221_X2 _3959_ (.A(_1320_),
    .B1(_1324_),
    .B2(_1040_),
    .C1(_1254_),
    .C2(_1319_),
    .ZN(_0137_));
 AND4_X1 _3960_ (.A1(_1093_),
    .A2(_1154_),
    .A3(_1176_),
    .A4(_1275_),
    .ZN(_1325_));
 AOI22_X1 _3961_ (.A1(_0404_),
    .A2(_1120_),
    .B1(_1325_),
    .B2(_1246_),
    .ZN(_1326_));
 NAND2_X1 _3962_ (.A1(_1185_),
    .A2(_1231_),
    .ZN(_1327_));
 OAI221_X1 _3963_ (.A(_1326_),
    .B1(_1327_),
    .B2(_1209_),
    .C1(_1186_),
    .C2(_1242_),
    .ZN(_0138_));
 NOR3_X4 _3964_ (.A1(_0995_),
    .A2(_1118_),
    .A3(_1004_),
    .ZN(_1328_));
 NAND3_X4 _3965_ (.A1(_0994_),
    .A2(_1225_),
    .A3(_1328_),
    .ZN(_1329_));
 MUX2_X1 _3966_ (.A(net47),
    .B(net51),
    .S(_1070_),
    .Z(_1330_));
 MUX2_X1 _3967_ (.A(net50),
    .B(net52),
    .S(_1070_),
    .Z(_1331_));
 MUX2_X1 _3968_ (.A(_1330_),
    .B(_1331_),
    .S(_1057_),
    .Z(_1332_));
 INV_X1 _3969_ (.A(net33),
    .ZN(_1333_));
 MUX2_X1 _3970_ (.A(_2050_),
    .B(_1333_),
    .S(_0987_),
    .Z(_1334_));
 NOR2_X1 _3971_ (.A1(_0992_),
    .A2(_1334_),
    .ZN(_1335_));
 MUX2_X1 _3972_ (.A(_1332_),
    .B(_1335_),
    .S(_1067_),
    .Z(_1336_));
 AOI211_X4 _3973_ (.A(_2083_),
    .B(_0990_),
    .C1(_0961_),
    .C2(_0991_),
    .ZN(_1337_));
 AOI211_X2 _3974_ (.A(_0986_),
    .B(_1337_),
    .C1(_1071_),
    .C2(_1575_),
    .ZN(_1338_));
 MUX2_X1 _3975_ (.A(_2086_),
    .B(_2080_),
    .S(_1071_),
    .Z(_1339_));
 AOI21_X1 _3976_ (.A(_1338_),
    .B1(_1339_),
    .B2(_1074_),
    .ZN(_1340_));
 NAND3_X1 _3977_ (.A1(_1074_),
    .A2(_1571_),
    .A3(_0992_),
    .ZN(_1341_));
 NAND3_X1 _3978_ (.A1(_1058_),
    .A2(_1572_),
    .A3(_0992_),
    .ZN(_1342_));
 NAND3_X1 _3979_ (.A1(_1074_),
    .A2(_1573_),
    .A3(_1076_),
    .ZN(_1343_));
 NAND3_X1 _3980_ (.A1(_1057_),
    .A2(_1574_),
    .A3(_1076_),
    .ZN(_1344_));
 NAND4_X1 _3981_ (.A1(_1341_),
    .A2(_1342_),
    .A3(_1343_),
    .A4(_1344_),
    .ZN(_1345_));
 MUX2_X1 _3982_ (.A(_1340_),
    .B(_1345_),
    .S(_1067_),
    .Z(_1346_));
 AOI221_X2 _3983_ (.A(_1087_),
    .B1(_1088_),
    .B2(_1336_),
    .C1(_1346_),
    .C2(_1056_),
    .ZN(_1347_));
 MUX2_X1 _3984_ (.A(_1579_),
    .B(net39),
    .S(_1076_),
    .Z(_1348_));
 NOR3_X2 _3985_ (.A1(_1060_),
    .A2(_1067_),
    .A3(_1348_),
    .ZN(_1349_));
 MUX2_X1 _3986_ (.A(_1580_),
    .B(_1581_),
    .S(_1131_),
    .Z(_1350_));
 NOR3_X2 _3987_ (.A1(_1075_),
    .A2(_1067_),
    .A3(_1350_),
    .ZN(_1351_));
 MUX2_X1 _3988_ (.A(_1576_),
    .B(_1577_),
    .S(_1080_),
    .Z(_1352_));
 NOR3_X2 _3989_ (.A1(_1079_),
    .A2(_1105_),
    .A3(_1352_),
    .ZN(_1353_));
 MUX2_X1 _3990_ (.A(net37),
    .B(_1578_),
    .S(_1076_),
    .Z(_1354_));
 NOR3_X2 _3991_ (.A1(_1075_),
    .A2(_0985_),
    .A3(_1354_),
    .ZN(_1355_));
 NOR4_X4 _3992_ (.A1(_1349_),
    .A2(_1351_),
    .A3(_1353_),
    .A4(_1355_),
    .ZN(_1356_));
 MUX2_X1 _3993_ (.A(_1582_),
    .B(_1003_),
    .S(_1057_),
    .Z(_1357_));
 AND3_X2 _3994_ (.A1(_1093_),
    .A2(_1127_),
    .A3(_1357_),
    .ZN(_1358_));
 AOI22_X4 _3995_ (.A1(_1088_),
    .A2(_1356_),
    .B1(_1358_),
    .B2(_1149_),
    .ZN(_1359_));
 AOI211_X2 _3996_ (.A(_1329_),
    .B(_1347_),
    .C1(_1359_),
    .C2(_1087_),
    .ZN(_0139_));
 MUX2_X1 _3997_ (.A(net39),
    .B(_1580_),
    .S(_0986_),
    .Z(_1360_));
 MUX2_X1 _3998_ (.A(_1582_),
    .B(_1581_),
    .S(_2118_),
    .Z(_1361_));
 MUX2_X1 _3999_ (.A(_1360_),
    .B(_1361_),
    .S(_1080_),
    .Z(_1362_));
 AND4_X1 _4000_ (.A1(_1041_),
    .A2(_0985_),
    .A3(_1100_),
    .A4(_1362_),
    .ZN(_1363_));
 AOI211_X2 _4001_ (.A(_2071_),
    .B(_0990_),
    .C1(_0971_),
    .C2(_0991_),
    .ZN(_1364_));
 AOI211_X2 _4002_ (.A(_1057_),
    .B(_1364_),
    .C1(_1071_),
    .C2(_1578_),
    .ZN(_1365_));
 AOI211_X4 _4003_ (.A(_2104_),
    .B(_0990_),
    .C1(_0971_),
    .C2(_0991_),
    .ZN(_1366_));
 AOI211_X2 _4004_ (.A(_0986_),
    .B(_1366_),
    .C1(_1071_),
    .C2(_1579_),
    .ZN(_1367_));
 NOR4_X2 _4005_ (.A1(_0963_),
    .A2(_0985_),
    .A3(_1365_),
    .A4(_1367_),
    .ZN(_1368_));
 NAND2_X1 _4006_ (.A1(_0987_),
    .A2(_1003_),
    .ZN(_1369_));
 NOR3_X2 _4007_ (.A1(_1132_),
    .A2(_1163_),
    .A3(_1369_),
    .ZN(_1370_));
 AOI221_X2 _4008_ (.A(_1363_),
    .B1(_1368_),
    .B2(_1100_),
    .C1(_1370_),
    .C2(_0964_),
    .ZN(_1371_));
 AND2_X1 _4009_ (.A1(_1087_),
    .A2(_1371_),
    .ZN(_1372_));
 AOI211_X4 _4010_ (.A(_2080_),
    .B(_0990_),
    .C1(_0971_),
    .C2(_0991_),
    .ZN(_1373_));
 AOI211_X2 _4011_ (.A(_0987_),
    .B(_1373_),
    .C1(_1080_),
    .C2(_1576_),
    .ZN(_1374_));
 AOI211_X2 _4012_ (.A(_1057_),
    .B(_1337_),
    .C1(_1071_),
    .C2(_1575_),
    .ZN(_1375_));
 NOR3_X1 _4013_ (.A1(_1178_),
    .A2(_1374_),
    .A3(_1375_),
    .ZN(_1376_));
 MUX2_X1 _4014_ (.A(_1573_),
    .B(_1572_),
    .S(_0986_),
    .Z(_1377_));
 MUX2_X1 _4015_ (.A(net34),
    .B(_1574_),
    .S(_0987_),
    .Z(_1378_));
 MUX2_X1 _4016_ (.A(_1377_),
    .B(_1378_),
    .S(_1131_),
    .Z(_1379_));
 AND3_X1 _4017_ (.A1(_1097_),
    .A2(_1137_),
    .A3(_1379_),
    .ZN(_1380_));
 NOR3_X1 _4018_ (.A1(_1273_),
    .A2(_1376_),
    .A3(_1380_),
    .ZN(_1381_));
 AOI21_X1 _4019_ (.A(_1059_),
    .B1(net38),
    .B2(_1139_),
    .ZN(_1382_));
 MUX2_X1 _4020_ (.A(net33),
    .B(net47),
    .S(_1080_),
    .Z(_1383_));
 INV_X1 _4021_ (.A(_1383_),
    .ZN(_1384_));
 AOI21_X1 _4022_ (.A(_1382_),
    .B1(_1384_),
    .B2(_1079_),
    .ZN(_1385_));
 MUX2_X1 _4023_ (.A(net51),
    .B(_1571_),
    .S(_1080_),
    .Z(_1386_));
 MUX2_X1 _4024_ (.A(_1331_),
    .B(_1386_),
    .S(_1079_),
    .Z(_1387_));
 AOI221_X2 _4025_ (.A(_1247_),
    .B1(_1385_),
    .B2(_1127_),
    .C1(_1387_),
    .C2(_1160_),
    .ZN(_1388_));
 NOR4_X1 _4026_ (.A1(_1329_),
    .A2(_1372_),
    .A3(_1381_),
    .A4(_1388_),
    .ZN(_0150_));
 NAND2_X1 _4027_ (.A1(_1741_),
    .A2(inexact_stage2),
    .ZN(_1389_));
 AOI21_X1 _4028_ (.A(_1389_),
    .B1(_1680_),
    .B2(_1589_),
    .ZN(_0028_));
 CLKBUF_X3 _4029_ (.A(_1586_),
    .Z(_1390_));
 NOR4_X1 _4030_ (.A1(\aligned_a_mant[1] ),
    .A2(_0451_),
    .A3(\aligned_b_mant[1] ),
    .A4(_0452_),
    .ZN(_1391_));
 NOR2_X1 _4031_ (.A1(_1390_),
    .A2(_1391_),
    .ZN(_0029_));
 BUF_X2 _4032_ (.A(_1740_),
    .Z(_1392_));
 AND2_X1 _4033_ (.A1(_1392_),
    .A2(invalid_op_stage2),
    .ZN(_0030_));
 NAND2_X1 _4034_ (.A1(_2123_),
    .A2(_0387_),
    .ZN(_1393_));
 NAND2_X1 _4035_ (.A1(_0429_),
    .A2(_1393_),
    .ZN(_1394_));
 AOI221_X1 _4036_ (.A(invalid_op_stage2),
    .B1(_0387_),
    .B2(_0409_),
    .C1(_1394_),
    .C2(_0419_),
    .ZN(_1395_));
 NOR2_X1 _4037_ (.A1(_1390_),
    .A2(_1395_),
    .ZN(_0031_));
 NOR2_X1 _4038_ (.A1(_1390_),
    .A2(_0995_),
    .ZN(_0032_));
 NAND2_X2 _4039_ (.A1(_1117_),
    .A2(_1222_),
    .ZN(_1396_));
 BUF_X4 _4040_ (.A(_1396_),
    .Z(_1397_));
 MUX2_X1 _4041_ (.A(_2116_),
    .B(_2119_),
    .S(_1397_),
    .Z(_1398_));
 NOR2_X1 _4042_ (.A1(_1390_),
    .A2(_1398_),
    .ZN(_0033_));
 MUX2_X1 _4043_ (.A(_1994_),
    .B(_1998_),
    .S(_1397_),
    .Z(_1399_));
 NOR2_X1 _4044_ (.A1(_1390_),
    .A2(_1399_),
    .ZN(_0034_));
 MUX2_X1 _4045_ (.A(_2037_),
    .B(_2040_),
    .S(_1397_),
    .Z(_1400_));
 NOR2_X1 _4046_ (.A1(_1390_),
    .A2(_1400_),
    .ZN(_0035_));
 MUX2_X1 _4047_ (.A(_2031_),
    .B(_2034_),
    .S(_1397_),
    .Z(_1401_));
 NOR2_X1 _4048_ (.A1(_1390_),
    .A2(_1401_),
    .ZN(_0036_));
 MUX2_X1 _4049_ (.A(_2025_),
    .B(_2028_),
    .S(_1396_),
    .Z(_1402_));
 NOR2_X1 _4050_ (.A1(_1390_),
    .A2(_1402_),
    .ZN(_0037_));
 MUX2_X1 _4051_ (.A(_2019_),
    .B(_2022_),
    .S(_1396_),
    .Z(_1403_));
 NOR2_X1 _4052_ (.A1(_1390_),
    .A2(_1403_),
    .ZN(_0038_));
 MUX2_X1 _4053_ (.A(_2013_),
    .B(_2016_),
    .S(_1396_),
    .Z(_1404_));
 NOR2_X1 _4054_ (.A1(_1390_),
    .A2(_1404_),
    .ZN(_0039_));
 MUX2_X1 _4055_ (.A(_2007_),
    .B(_2010_),
    .S(_1396_),
    .Z(_1405_));
 NOR2_X1 _4056_ (.A1(_1714_),
    .A2(_1405_),
    .ZN(_0040_));
 NOR3_X1 _4057_ (.A1(_1837_),
    .A2(_1589_),
    .A3(_1744_),
    .ZN(_0041_));
 AND2_X1 _4058_ (.A1(_1392_),
    .A2(\final_mant[0] ),
    .ZN(_0042_));
 AND2_X1 _4059_ (.A1(_1392_),
    .A2(\final_mant[10] ),
    .ZN(_0043_));
 AND2_X1 _4060_ (.A1(_1392_),
    .A2(\final_mant[11] ),
    .ZN(_0044_));
 AND2_X1 _4061_ (.A1(_1392_),
    .A2(\final_mant[12] ),
    .ZN(_0045_));
 AND2_X1 _4062_ (.A1(_1392_),
    .A2(\final_mant[13] ),
    .ZN(_0046_));
 AND2_X1 _4063_ (.A1(_1392_),
    .A2(\final_mant[14] ),
    .ZN(_0047_));
 AND2_X1 _4064_ (.A1(_1392_),
    .A2(\final_mant[15] ),
    .ZN(_0048_));
 AND2_X1 _4065_ (.A1(_1392_),
    .A2(\final_mant[16] ),
    .ZN(_0049_));
 AND2_X1 _4066_ (.A1(_1392_),
    .A2(\final_mant[17] ),
    .ZN(_0050_));
 BUF_X2 _4067_ (.A(_1740_),
    .Z(_1406_));
 AND2_X1 _4068_ (.A1(_1406_),
    .A2(\final_mant[18] ),
    .ZN(_0051_));
 AND2_X1 _4069_ (.A1(_1406_),
    .A2(\final_mant[19] ),
    .ZN(_0052_));
 AND2_X1 _4070_ (.A1(_1406_),
    .A2(\final_mant[1] ),
    .ZN(_0053_));
 AND2_X1 _4071_ (.A1(_1406_),
    .A2(\final_mant[20] ),
    .ZN(_0054_));
 AND2_X1 _4072_ (.A1(_1406_),
    .A2(\final_mant[21] ),
    .ZN(_0055_));
 AND2_X1 _4073_ (.A1(_1406_),
    .A2(\final_mant[22] ),
    .ZN(_0056_));
 NOR2_X1 _4074_ (.A1(_1714_),
    .A2(_1749_),
    .ZN(_0057_));
 AND2_X1 _4075_ (.A1(_1406_),
    .A2(\final_exp[1] ),
    .ZN(_0058_));
 NOR2_X1 _4076_ (.A1(_1714_),
    .A2(_1761_),
    .ZN(_0059_));
 NOR2_X1 _4077_ (.A1(_1714_),
    .A2(_1771_),
    .ZN(_0060_));
 NOR2_X1 _4078_ (.A1(_1714_),
    .A2(_1781_),
    .ZN(_0061_));
 NOR2_X1 _4079_ (.A1(_1714_),
    .A2(_1788_),
    .ZN(_0062_));
 AND2_X1 _4080_ (.A1(_1406_),
    .A2(\final_exp[6] ),
    .ZN(_0063_));
 AND2_X1 _4081_ (.A1(_1406_),
    .A2(\final_mant[2] ),
    .ZN(_0064_));
 AND2_X1 _4082_ (.A1(_1406_),
    .A2(\final_exp[7] ),
    .ZN(_0065_));
 BUF_X2 _4083_ (.A(_1740_),
    .Z(_1407_));
 AND2_X1 _4084_ (.A1(_1407_),
    .A2(result_sign_stage2),
    .ZN(_0066_));
 AND2_X1 _4085_ (.A1(_1407_),
    .A2(\final_mant[3] ),
    .ZN(_0067_));
 AND2_X1 _4086_ (.A1(_1407_),
    .A2(\final_mant[4] ),
    .ZN(_0068_));
 AND2_X1 _4087_ (.A1(_1407_),
    .A2(\final_mant[5] ),
    .ZN(_0069_));
 AND2_X1 _4088_ (.A1(_1407_),
    .A2(\final_mant[6] ),
    .ZN(_0070_));
 AND2_X1 _4089_ (.A1(_1407_),
    .A2(\final_mant[7] ),
    .ZN(_0071_));
 AND2_X1 _4090_ (.A1(_1407_),
    .A2(\final_mant[8] ),
    .ZN(_0072_));
 AND2_X1 _4091_ (.A1(_1407_),
    .A2(\final_mant[9] ),
    .ZN(_0073_));
 AND2_X1 _4092_ (.A1(_1407_),
    .A2(\larger_exp_stage1[0] ),
    .ZN(_0074_));
 AND2_X1 _4093_ (.A1(_1407_),
    .A2(\larger_exp_stage1[1] ),
    .ZN(_0075_));
 CLKBUF_X2 _4094_ (.A(_1740_),
    .Z(_1408_));
 AND2_X1 _4095_ (.A1(_1408_),
    .A2(\larger_exp_stage1[2] ),
    .ZN(_0076_));
 AND2_X1 _4096_ (.A1(_1408_),
    .A2(\larger_exp_stage1[3] ),
    .ZN(_0077_));
 AND2_X1 _4097_ (.A1(_1408_),
    .A2(\larger_exp_stage1[4] ),
    .ZN(_0078_));
 AND2_X1 _4098_ (.A1(_1408_),
    .A2(\larger_exp_stage1[5] ),
    .ZN(_0079_));
 AND2_X1 _4099_ (.A1(_1408_),
    .A2(\larger_exp_stage1[6] ),
    .ZN(_0080_));
 AND2_X1 _4100_ (.A1(_1408_),
    .A2(\larger_exp_stage1[7] ),
    .ZN(_0081_));
 AND2_X1 _4101_ (.A1(_1408_),
    .A2(valid_stage2),
    .ZN(_0084_));
 AND2_X1 _4102_ (.A1(_1408_),
    .A2(net53),
    .ZN(_0085_));
 AND2_X1 _4103_ (.A1(_1408_),
    .A2(valid_stage1),
    .ZN(_0086_));
 AND2_X1 _4104_ (.A1(_1408_),
    .A2(net25),
    .ZN(_0087_));
 NOR3_X1 _4105_ (.A1(_0831_),
    .A2(_0419_),
    .A3(_0387_),
    .ZN(_1409_));
 NAND2_X1 _4106_ (.A1(_0835_),
    .A2(_0826_),
    .ZN(_1410_));
 NAND3_X1 _4107_ (.A1(_2306_),
    .A2(_0815_),
    .A3(_0806_),
    .ZN(_1411_));
 AOI21_X1 _4108_ (.A(_0746_),
    .B1(_0748_),
    .B2(_0631_),
    .ZN(_1412_));
 AOI21_X1 _4109_ (.A(_0790_),
    .B1(_1411_),
    .B2(_1412_),
    .ZN(_1413_));
 OAI21_X1 _4110_ (.A(_0806_),
    .B1(_2330_),
    .B2(_0815_),
    .ZN(_1414_));
 AOI21_X1 _4111_ (.A(_0500_),
    .B1(_1414_),
    .B2(_0835_),
    .ZN(_1415_));
 AOI21_X1 _4112_ (.A(_2320_),
    .B1(_2312_),
    .B2(_0764_),
    .ZN(_1416_));
 OAI21_X1 _4113_ (.A(_0818_),
    .B1(_1416_),
    .B2(_0815_),
    .ZN(_1417_));
 AOI21_X1 _4114_ (.A(_2336_),
    .B1(_1417_),
    .B2(_0805_),
    .ZN(_1418_));
 NAND2_X1 _4115_ (.A1(_0411_),
    .A2(_1418_),
    .ZN(_1419_));
 AOI21_X1 _4116_ (.A(_2317_),
    .B1(_2309_),
    .B2(_0764_),
    .ZN(_1420_));
 OAI21_X1 _4117_ (.A(_0816_),
    .B1(_1420_),
    .B2(_0815_),
    .ZN(_1421_));
 AOI21_X1 _4118_ (.A(_2333_),
    .B1(_1421_),
    .B2(_0805_),
    .ZN(_1422_));
 NAND2_X1 _4119_ (.A1(_0738_),
    .A2(_1422_),
    .ZN(_1423_));
 NOR4_X1 _4120_ (.A1(_0780_),
    .A2(_0766_),
    .A3(_0815_),
    .A4(_0806_),
    .ZN(_1424_));
 AOI221_X2 _4121_ (.A(_0465_),
    .B1(_1419_),
    .B2(_1423_),
    .C1(_1424_),
    .C2(_0761_),
    .ZN(_1425_));
 OAI221_X1 _4122_ (.A(_1409_),
    .B1(_1410_),
    .B2(_1413_),
    .C1(_1415_),
    .C2(_1425_),
    .ZN(_1426_));
 NAND2_X1 _4123_ (.A1(_0831_),
    .A2(_0431_),
    .ZN(_1427_));
 OR2_X1 _4124_ (.A1(_1415_),
    .A2(_1425_),
    .ZN(_1428_));
 OAI21_X1 _4125_ (.A(_1426_),
    .B1(_1427_),
    .B2(_1428_),
    .ZN(_1429_));
 NOR3_X1 _4126_ (.A1(_1413_),
    .A2(_1410_),
    .A3(_1427_),
    .ZN(_1430_));
 NOR3_X1 _4127_ (.A1(_1837_),
    .A2(_1429_),
    .A3(_1430_),
    .ZN(_0103_));
 AND3_X1 _4128_ (.A1(_0994_),
    .A2(_1225_),
    .A3(_1328_),
    .ZN(_1431_));
 NAND2_X4 _4129_ (.A1(_1124_),
    .A2(_1431_),
    .ZN(_1432_));
 MUX2_X1 _4130_ (.A(net36),
    .B(_1576_),
    .S(_1131_),
    .Z(_1433_));
 MUX2_X1 _4131_ (.A(_1575_),
    .B(net37),
    .S(_1080_),
    .Z(_1434_));
 MUX2_X1 _4132_ (.A(_1433_),
    .B(_1434_),
    .S(_1059_),
    .Z(_1435_));
 MUX2_X1 _4133_ (.A(_1573_),
    .B(net34),
    .S(_1131_),
    .Z(_1436_));
 MUX2_X1 _4134_ (.A(_1574_),
    .B(net35),
    .S(_1131_),
    .Z(_1437_));
 MUX2_X1 _4135_ (.A(_1436_),
    .B(_1437_),
    .S(_1079_),
    .Z(_1438_));
 MUX2_X1 _4136_ (.A(_1435_),
    .B(_1438_),
    .S(_1097_),
    .Z(_1439_));
 NAND2_X1 _4137_ (.A1(_0987_),
    .A2(_1579_),
    .ZN(_1440_));
 NAND2_X1 _4138_ (.A1(_1057_),
    .A2(_1580_),
    .ZN(_1441_));
 AOI21_X1 _4139_ (.A(_1092_),
    .B1(_1440_),
    .B2(_1441_),
    .ZN(_1442_));
 NAND2_X1 _4140_ (.A1(_1074_),
    .A2(_1577_),
    .ZN(_1443_));
 NAND2_X1 _4141_ (.A1(_1058_),
    .A2(_1578_),
    .ZN(_1444_));
 AOI21_X1 _4142_ (.A(_1139_),
    .B1(_1443_),
    .B2(_1444_),
    .ZN(_1445_));
 NOR2_X1 _4143_ (.A1(_1442_),
    .A2(_1445_),
    .ZN(_1446_));
 MUX2_X1 _4144_ (.A(_1581_),
    .B(net39),
    .S(_0986_),
    .Z(_1447_));
 MUX2_X1 _4145_ (.A(_1357_),
    .B(_1447_),
    .S(_1092_),
    .Z(_1448_));
 NAND2_X2 _4146_ (.A1(_1137_),
    .A2(_1448_),
    .ZN(_1449_));
 OAI22_X4 _4147_ (.A1(_1163_),
    .A2(_1446_),
    .B1(_1449_),
    .B2(_1097_),
    .ZN(_1450_));
 AOI22_X2 _4148_ (.A1(_1215_),
    .A2(_1439_),
    .B1(_1450_),
    .B2(_1149_),
    .ZN(_1451_));
 NAND2_X4 _4149_ (.A1(_1740_),
    .A2(_1397_),
    .ZN(_1452_));
 OAI22_X2 _4150_ (.A1(_1432_),
    .A2(_1451_),
    .B1(_1452_),
    .B2(_2092_),
    .ZN(_0140_));
 NOR2_X4 _4151_ (.A1(_0999_),
    .A2(_1152_),
    .ZN(_1453_));
 INV_X1 _4152_ (.A(_1369_),
    .ZN(_1454_));
 MUX2_X1 _4153_ (.A(_1454_),
    .B(_1361_),
    .S(_0992_),
    .Z(_1455_));
 MUX2_X1 _4154_ (.A(_1578_),
    .B(_1580_),
    .S(_1076_),
    .Z(_1456_));
 MUX2_X1 _4155_ (.A(_1348_),
    .B(_1456_),
    .S(_0988_),
    .Z(_1457_));
 MUX2_X1 _4156_ (.A(_1455_),
    .B(_1457_),
    .S(_1097_),
    .Z(_1458_));
 NOR2_X1 _4157_ (.A1(_1153_),
    .A2(_1458_),
    .ZN(_1459_));
 MUX2_X1 _4158_ (.A(_1352_),
    .B(_1434_),
    .S(_0988_),
    .Z(_1460_));
 MUX2_X1 _4159_ (.A(net34),
    .B(net36),
    .S(_1131_),
    .Z(_1461_));
 MUX2_X1 _4160_ (.A(_1461_),
    .B(_1437_),
    .S(_0988_),
    .Z(_1462_));
 MUX2_X1 _4161_ (.A(_1460_),
    .B(_1462_),
    .S(_1097_),
    .Z(_1463_));
 NOR2_X1 _4162_ (.A1(_1149_),
    .A2(_1463_),
    .ZN(_1464_));
 OAI33_X1 _4163_ (.A1(_1813_),
    .A2(_2089_),
    .A3(_1453_),
    .B1(_1459_),
    .B2(_1464_),
    .B3(_1432_),
    .ZN(_0141_));
 NAND2_X1 _4164_ (.A1(_1440_),
    .A2(_1441_),
    .ZN(_1465_));
 MUX2_X1 _4165_ (.A(_1447_),
    .B(_1465_),
    .S(_1069_),
    .Z(_1466_));
 MUX2_X1 _4166_ (.A(_1447_),
    .B(_1465_),
    .S(_0989_),
    .Z(_1467_));
 MUX2_X1 _4167_ (.A(_1466_),
    .B(_1467_),
    .S(_0981_),
    .Z(_1468_));
 INV_X1 _4168_ (.A(_1468_),
    .ZN(_1469_));
 NAND2_X1 _4169_ (.A1(_1093_),
    .A2(_1357_),
    .ZN(_1470_));
 OAI22_X4 _4170_ (.A1(_1163_),
    .A2(_1469_),
    .B1(_1470_),
    .B2(_1178_),
    .ZN(_1471_));
 MUX2_X1 _4171_ (.A(_1352_),
    .B(_1354_),
    .S(_1059_),
    .Z(_1472_));
 MUX2_X1 _4172_ (.A(_1340_),
    .B(_1472_),
    .S(_1105_),
    .Z(_1473_));
 AOI22_X1 _4173_ (.A1(_1149_),
    .A2(_1471_),
    .B1(_1473_),
    .B2(_1215_),
    .ZN(_1474_));
 OAI22_X1 _4174_ (.A1(_2086_),
    .A2(_1452_),
    .B1(_1474_),
    .B2(_1432_),
    .ZN(_0142_));
 AOI21_X1 _4175_ (.A(_1092_),
    .B1(_1361_),
    .B2(_1067_),
    .ZN(_1475_));
 OAI21_X1 _4176_ (.A(_1369_),
    .B1(_1066_),
    .B2(_1063_),
    .ZN(_1476_));
 OAI21_X1 _4177_ (.A(_1476_),
    .B1(_1360_),
    .B2(_0985_),
    .ZN(_1477_));
 AOI21_X2 _4178_ (.A(_1475_),
    .B1(_1477_),
    .B2(_1093_),
    .ZN(_1478_));
 AOI21_X1 _4179_ (.A(_1153_),
    .B1(_1137_),
    .B2(_1478_),
    .ZN(_1479_));
 OAI33_X1 _4180_ (.A1(_1178_),
    .A2(_1365_),
    .A3(_1367_),
    .B1(_1374_),
    .B2(_1375_),
    .B3(_1163_),
    .ZN(_1480_));
 NOR2_X1 _4181_ (.A1(_1149_),
    .A2(_1480_),
    .ZN(_1481_));
 OAI33_X1 _4182_ (.A1(_1813_),
    .A2(_2083_),
    .A3(_1453_),
    .B1(_1479_),
    .B2(_1481_),
    .B3(_1432_),
    .ZN(_0143_));
 OR2_X1 _4183_ (.A1(_1442_),
    .A2(_1445_),
    .ZN(_1482_));
 AOI22_X1 _4184_ (.A1(_1154_),
    .A2(_1435_),
    .B1(_1482_),
    .B2(_1160_),
    .ZN(_1483_));
 NAND3_X1 _4185_ (.A1(_1189_),
    .A2(_1137_),
    .A3(_1448_),
    .ZN(_1484_));
 MUX2_X1 _4186_ (.A(_1483_),
    .B(_1484_),
    .S(_1149_),
    .Z(_1485_));
 OAI22_X1 _4187_ (.A1(_2080_),
    .A2(_1452_),
    .B1(_1485_),
    .B2(_1432_),
    .ZN(_0144_));
 AND3_X1 _4188_ (.A1(_0964_),
    .A2(_1189_),
    .A3(_1455_),
    .ZN(_1486_));
 MUX2_X1 _4189_ (.A(_1457_),
    .B(_1460_),
    .S(_1189_),
    .Z(_1487_));
 AOI21_X1 _4190_ (.A(_1486_),
    .B1(_1487_),
    .B2(_1153_),
    .ZN(_1488_));
 OAI22_X1 _4191_ (.A1(_2077_),
    .A2(_1452_),
    .B1(_1488_),
    .B2(_1432_),
    .ZN(_0145_));
 OAI22_X2 _4192_ (.A1(_1359_),
    .A2(_1432_),
    .B1(_1452_),
    .B2(_2074_),
    .ZN(_0146_));
 NOR3_X2 _4193_ (.A1(_0995_),
    .A2(_0999_),
    .A3(_1004_),
    .ZN(_1489_));
 NAND3_X1 _4194_ (.A1(_1124_),
    .A2(_1225_),
    .A3(_1489_),
    .ZN(_1490_));
 OAI22_X1 _4195_ (.A1(_1490_),
    .A2(_1371_),
    .B1(_1453_),
    .B2(_2071_),
    .ZN(_1491_));
 AND2_X1 _4196_ (.A1(_1750_),
    .A2(_1491_),
    .ZN(_0147_));
 AND3_X2 _4197_ (.A1(_1225_),
    .A2(_1234_),
    .A3(_1489_),
    .ZN(_1492_));
 AOI22_X2 _4198_ (.A1(_1577_),
    .A2(_1397_),
    .B1(_1450_),
    .B2(_1492_),
    .ZN(_1493_));
 NOR2_X1 _4199_ (.A1(_1714_),
    .A2(_1493_),
    .ZN(_0148_));
 NAND2_X1 _4200_ (.A1(_1458_),
    .A2(_1492_),
    .ZN(_1494_));
 NAND2_X1 _4201_ (.A1(_1578_),
    .A2(_1397_),
    .ZN(_1495_));
 AOI21_X1 _4202_ (.A(_1813_),
    .B1(_1494_),
    .B2(_1495_),
    .ZN(_0149_));
 NAND2_X1 _4203_ (.A1(_1153_),
    .A2(_1471_),
    .ZN(_1496_));
 OAI22_X2 _4204_ (.A1(_2098_),
    .A2(_1452_),
    .B1(_1496_),
    .B2(_1432_),
    .ZN(_0151_));
 AOI22_X1 _4205_ (.A1(_1580_),
    .A2(_1397_),
    .B1(_1478_),
    .B2(_1492_),
    .ZN(_1497_));
 NOR2_X1 _4206_ (.A1(_1714_),
    .A2(_1497_),
    .ZN(_0152_));
 NAND3_X1 _4207_ (.A1(_1225_),
    .A2(_1234_),
    .A3(_1489_),
    .ZN(_1498_));
 OAI22_X1 _4208_ (.A1(_2110_),
    .A2(_1453_),
    .B1(_1484_),
    .B2(_1498_),
    .ZN(_1499_));
 AND2_X1 _4209_ (.A1(_1750_),
    .A2(_1499_),
    .ZN(_0153_));
 NAND2_X1 _4210_ (.A1(_1581_),
    .A2(_1397_),
    .ZN(_1500_));
 NAND3_X1 _4211_ (.A1(_1154_),
    .A2(_1455_),
    .A3(_1492_),
    .ZN(_1501_));
 AOI21_X1 _4212_ (.A(_1813_),
    .B1(_1500_),
    .B2(_1501_),
    .ZN(_0154_));
 AOI22_X2 _4213_ (.A1(_1582_),
    .A2(_1397_),
    .B1(_1492_),
    .B2(_1358_),
    .ZN(_1502_));
 NOR2_X1 _4214_ (.A1(_1714_),
    .A2(_1502_),
    .ZN(_0155_));
 OAI21_X1 _4215_ (.A(_1453_),
    .B1(_1498_),
    .B2(_1270_),
    .ZN(_1503_));
 AND3_X1 _4216_ (.A1(_1750_),
    .A2(_1003_),
    .A3(_1503_),
    .ZN(_0156_));
 NOR2_X1 _4217_ (.A1(_1055_),
    .A2(_1247_),
    .ZN(_1504_));
 MUX2_X1 _4218_ (.A(net52),
    .B(_1572_),
    .S(_1076_),
    .Z(_1505_));
 MUX2_X1 _4219_ (.A(_1386_),
    .B(_1505_),
    .S(_1059_),
    .Z(_1506_));
 MUX2_X1 _4220_ (.A(net38),
    .B(net50),
    .S(_1076_),
    .Z(_1507_));
 MUX2_X1 _4221_ (.A(_1383_),
    .B(_1507_),
    .S(_1059_),
    .Z(_1508_));
 MUX2_X1 _4222_ (.A(_1506_),
    .B(_1508_),
    .S(_1097_),
    .Z(_1509_));
 AOI222_X2 _4223_ (.A1(_1314_),
    .A2(_1439_),
    .B1(_1450_),
    .B2(_1275_),
    .C1(_1504_),
    .C2(_1509_),
    .ZN(_1510_));
 OAI22_X1 _4224_ (.A1(_1333_),
    .A2(_1452_),
    .B1(_1510_),
    .B2(_1329_),
    .ZN(_0157_));
 AOI21_X1 _4225_ (.A(_1124_),
    .B1(_1215_),
    .B2(_1458_),
    .ZN(_1511_));
 AOI221_X2 _4226_ (.A(_1041_),
    .B1(_1160_),
    .B2(_1460_),
    .C1(_1462_),
    .C2(_1127_),
    .ZN(_1512_));
 NOR2_X1 _4227_ (.A1(_1060_),
    .A2(_1507_),
    .ZN(_1513_));
 OAI21_X1 _4228_ (.A(_1127_),
    .B1(_1330_),
    .B2(_1075_),
    .ZN(_1514_));
 NOR2_X1 _4229_ (.A1(_1513_),
    .A2(_1514_),
    .ZN(_1515_));
 MUX2_X1 _4230_ (.A(_1571_),
    .B(net52),
    .S(_0987_),
    .Z(_1516_));
 MUX2_X1 _4231_ (.A(_1377_),
    .B(_1516_),
    .S(_0992_),
    .Z(_1517_));
 NAND2_X1 _4232_ (.A1(_1100_),
    .A2(_1517_),
    .ZN(_1518_));
 OAI21_X1 _4233_ (.A(_1234_),
    .B1(_1518_),
    .B2(_1189_),
    .ZN(_1519_));
 OAI21_X1 _4234_ (.A(_1431_),
    .B1(_1515_),
    .B2(_1519_),
    .ZN(_1520_));
 OAI33_X1 _4235_ (.A1(_1813_),
    .A2(_2050_),
    .A3(_1453_),
    .B1(_1511_),
    .B2(_1512_),
    .B3(_1520_),
    .ZN(_0158_));
 AOI221_X1 _4236_ (.A(_1247_),
    .B1(_1332_),
    .B2(_1127_),
    .C1(_1345_),
    .C2(_1160_),
    .ZN(_1521_));
 OAI21_X1 _4237_ (.A(_1431_),
    .B1(_1471_),
    .B2(_1124_),
    .ZN(_1522_));
 NOR2_X1 _4238_ (.A1(_1087_),
    .A2(_1055_),
    .ZN(_1523_));
 AOI21_X1 _4239_ (.A(_1153_),
    .B1(_1473_),
    .B2(_1523_),
    .ZN(_1524_));
 OAI33_X1 _4240_ (.A1(_1813_),
    .A2(_2056_),
    .A3(_1453_),
    .B1(_1521_),
    .B2(_1522_),
    .B3(_1524_),
    .ZN(_0159_));
 AND2_X1 _4241_ (.A1(_1100_),
    .A2(_1379_),
    .ZN(_1525_));
 AOI221_X2 _4242_ (.A(_1247_),
    .B1(_1525_),
    .B2(_1105_),
    .C1(_1387_),
    .C2(_1127_),
    .ZN(_1526_));
 AOI221_X2 _4243_ (.A(_1234_),
    .B1(_1480_),
    .B2(_1123_),
    .C1(_1478_),
    .C2(_1088_),
    .ZN(_1527_));
 OAI33_X1 _4244_ (.A1(_1813_),
    .A2(_2053_),
    .A3(_1453_),
    .B1(_1526_),
    .B2(_1527_),
    .B3(_1329_),
    .ZN(_0160_));
 NOR2_X1 _4245_ (.A1(_1060_),
    .A2(_1386_),
    .ZN(_1528_));
 NOR2_X1 _4246_ (.A1(_1075_),
    .A2(_1505_),
    .ZN(_1529_));
 NAND2_X1 _4247_ (.A1(_1123_),
    .A2(_1137_),
    .ZN(_1530_));
 OAI33_X1 _4248_ (.A1(_0964_),
    .A2(_1124_),
    .A3(_1449_),
    .B1(_1528_),
    .B2(_1529_),
    .B3(_1530_),
    .ZN(_1531_));
 MUX2_X1 _4249_ (.A(_2092_),
    .B(_2086_),
    .S(_1131_),
    .Z(_1532_));
 MUX2_X1 _4250_ (.A(_2089_),
    .B(_2083_),
    .S(_1076_),
    .Z(_1533_));
 MUX2_X1 _4251_ (.A(_1532_),
    .B(_1533_),
    .S(_1079_),
    .Z(_1534_));
 OAI21_X1 _4252_ (.A(_1041_),
    .B1(_1178_),
    .B2(_1534_),
    .ZN(_1535_));
 AOI22_X1 _4253_ (.A1(_1189_),
    .A2(_1531_),
    .B1(_1535_),
    .B2(_1124_),
    .ZN(_1536_));
 AND2_X1 _4254_ (.A1(_1187_),
    .A2(_1483_),
    .ZN(_1537_));
 OAI33_X1 _4255_ (.A1(_1813_),
    .A2(_2068_),
    .A3(_1453_),
    .B1(_1536_),
    .B2(_1537_),
    .B3(_1329_),
    .ZN(_0161_));
 AOI21_X1 _4256_ (.A(_1123_),
    .B1(_1067_),
    .B2(_1455_),
    .ZN(_1538_));
 NOR2_X1 _4257_ (.A1(_0973_),
    .A2(_1105_),
    .ZN(_1539_));
 MUX2_X1 _4258_ (.A(_1339_),
    .B(_1533_),
    .S(_0988_),
    .Z(_1540_));
 NOR2_X1 _4259_ (.A1(_0973_),
    .A2(_1097_),
    .ZN(_1541_));
 AOI221_X1 _4260_ (.A(_1538_),
    .B1(_1539_),
    .B2(_1518_),
    .C1(_1540_),
    .C2(_1541_),
    .ZN(_1542_));
 AOI22_X1 _4261_ (.A1(_1314_),
    .A2(_1487_),
    .B1(_1542_),
    .B2(_1215_),
    .ZN(_1543_));
 OAI22_X1 _4262_ (.A1(_2065_),
    .A2(_1452_),
    .B1(_1543_),
    .B2(_1329_),
    .ZN(_0162_));
 AOI222_X2 _4263_ (.A1(_1504_),
    .A2(_1346_),
    .B1(_1356_),
    .B2(_1314_),
    .C1(_1358_),
    .C2(_1275_),
    .ZN(_1544_));
 OAI22_X1 _4264_ (.A1(_2062_),
    .A2(_1452_),
    .B1(_1544_),
    .B2(_1329_),
    .ZN(_0163_));
 OAI21_X1 _4265_ (.A(_1234_),
    .B1(_1376_),
    .B2(_1380_),
    .ZN(_1545_));
 NOR2_X1 _4266_ (.A1(_1132_),
    .A2(_1360_),
    .ZN(_1546_));
 NOR2_X1 _4267_ (.A1(_1093_),
    .A2(_1361_),
    .ZN(_1547_));
 OAI33_X1 _4268_ (.A1(_1178_),
    .A2(_1546_),
    .A3(_1547_),
    .B1(_1365_),
    .B2(_1367_),
    .B3(_1163_),
    .ZN(_1548_));
 AOI22_X1 _4269_ (.A1(_1275_),
    .A2(_1370_),
    .B1(_1548_),
    .B2(_1187_),
    .ZN(_1549_));
 AND2_X1 _4270_ (.A1(_1545_),
    .A2(_1549_),
    .ZN(_1550_));
 OAI22_X1 _4271_ (.A1(_2059_),
    .A2(_1452_),
    .B1(_1550_),
    .B2(_1329_),
    .ZN(_0164_));
 AND2_X1 _4272_ (.A1(_1750_),
    .A2(net49),
    .ZN(_0165_));
 FA_X1 _4273_ (.A(_1994_),
    .B(net41),
    .CI(_1995_),
    .CO(_1996_),
    .S(_1997_));
 FA_X1 _4274_ (.A(net17),
    .B(_1998_),
    .CI(_1999_),
    .CO(_2000_),
    .S(_2001_));
 FA_X1 _4275_ (.A(_2002_),
    .B(_2003_),
    .CI(_2004_),
    .CO(_2005_),
    .S(_2006_));
 HA_X1 _4276_ (.A(_2007_),
    .B(net48),
    .CO(_2008_),
    .S(_2009_));
 HA_X1 _4277_ (.A(net24),
    .B(_2010_),
    .CO(_2011_),
    .S(_2012_));
 HA_X1 _4278_ (.A(_2013_),
    .B(net46),
    .CO(_2014_),
    .S(_2015_));
 HA_X1 _4279_ (.A(net22),
    .B(_2016_),
    .CO(_2017_),
    .S(_2018_));
 HA_X1 _4280_ (.A(_2019_),
    .B(net45),
    .CO(_2020_),
    .S(_2021_));
 HA_X1 _4281_ (.A(net21),
    .B(_2022_),
    .CO(_2023_),
    .S(_2024_));
 HA_X1 _4282_ (.A(_2025_),
    .B(net44),
    .CO(_2026_),
    .S(_2027_));
 HA_X1 _4283_ (.A(net20),
    .B(_2028_),
    .CO(_2029_),
    .S(_2030_));
 HA_X1 _4284_ (.A(_2031_),
    .B(net43),
    .CO(_2032_),
    .S(_2033_));
 HA_X1 _4285_ (.A(net19),
    .B(_2034_),
    .CO(_2035_),
    .S(_2036_));
 HA_X1 _4286_ (.A(_2037_),
    .B(net42),
    .CO(_2038_),
    .S(_2039_));
 HA_X1 _4287_ (.A(net18),
    .B(_2040_),
    .CO(_2041_),
    .S(_2042_));
 HA_X1 _4288_ (.A(_1994_),
    .B(net41),
    .CO(_2043_),
    .S(_2044_));
 HA_X1 _4289_ (.A(net17),
    .B(_1998_),
    .CO(_2045_),
    .S(_2046_));
 HA_X1 _4290_ (.A(_2047_),
    .B(net33),
    .CO(_2048_),
    .S(_2049_));
 HA_X1 _4291_ (.A(net12),
    .B(_2050_),
    .CO(_2051_),
    .S(_2052_));
 HA_X1 _4292_ (.A(net26),
    .B(_2053_),
    .CO(_2054_),
    .S(_2055_));
 HA_X1 _4293_ (.A(net23),
    .B(_2056_),
    .CO(_2057_),
    .S(_2058_));
 HA_X1 _4294_ (.A(net30),
    .B(_2059_),
    .CO(_2060_),
    .S(_2061_));
 HA_X1 _4295_ (.A(net29),
    .B(_2062_),
    .CO(_2063_),
    .S(_2064_));
 HA_X1 _4296_ (.A(net28),
    .B(_2065_),
    .CO(_2066_),
    .S(_2067_));
 HA_X1 _4297_ (.A(net27),
    .B(_2068_),
    .CO(_2069_),
    .S(_2070_));
 HA_X1 _4298_ (.A(net7),
    .B(_2071_),
    .CO(_2072_),
    .S(_2073_));
 HA_X1 _4299_ (.A(net6),
    .B(_2074_),
    .CO(_2075_),
    .S(_2076_));
 HA_X1 _4300_ (.A(net5),
    .B(_2077_),
    .CO(_2078_),
    .S(_2079_));
 HA_X1 _4301_ (.A(net4),
    .B(_2080_),
    .CO(_2081_),
    .S(_2082_));
 HA_X1 _4302_ (.A(net3),
    .B(_2083_),
    .CO(_2084_),
    .S(_2085_));
 HA_X1 _4303_ (.A(net2),
    .B(_2086_),
    .CO(_2087_),
    .S(_2088_));
 HA_X1 _4304_ (.A(net32),
    .B(_2089_),
    .CO(_2090_),
    .S(_2091_));
 HA_X1 _4305_ (.A(net31),
    .B(_2092_),
    .CO(_2093_),
    .S(_2094_));
 HA_X1 _4306_ (.A(net11),
    .B(_2095_),
    .CO(_2096_),
    .S(_2097_));
 HA_X1 _4307_ (.A(net10),
    .B(_2098_),
    .CO(_2099_),
    .S(_2100_));
 HA_X1 _4308_ (.A(net9),
    .B(_2101_),
    .CO(_2102_),
    .S(_2103_));
 HA_X1 _4309_ (.A(net8),
    .B(_2104_),
    .CO(_2105_),
    .S(_2106_));
 HA_X1 _4310_ (.A(net14),
    .B(_2107_),
    .CO(_2108_),
    .S(_2109_));
 HA_X1 _4311_ (.A(net13),
    .B(_2110_),
    .CO(_2111_),
    .S(_2112_));
 HA_X1 _4312_ (.A(net15),
    .B(_2113_),
    .CO(_2114_),
    .S(_2115_));
 HA_X1 _4313_ (.A(_2116_),
    .B(net40),
    .CO(_2117_),
    .S(_2118_));
 HA_X1 _4314_ (.A(net16),
    .B(_2119_),
    .CO(_2120_),
    .S(_2121_));
 HA_X1 _4315_ (.A(net25),
    .B(net49),
    .CO(_2122_),
    .S(_2123_));
 HA_X1 _4316_ (.A(_2124_),
    .B(_2125_),
    .CO(_2003_),
    .S(_2126_));
 HA_X1 _4317_ (.A(\result_exp_stage2[0] ),
    .B(_2127_),
    .CO(_2128_),
    .S(_2129_));
 HA_X1 _4318_ (.A(_2002_),
    .B(_2004_),
    .CO(_2130_),
    .S(_2131_));
 HA_X1 _4319_ (.A(\result_exp_stage2[1] ),
    .B(_2132_),
    .CO(_2133_),
    .S(_2134_));
 HA_X1 _4320_ (.A(_2135_),
    .B(_2136_),
    .CO(_2137_),
    .S(_2138_));
 HA_X1 _4321_ (.A(\result_exp_stage2[2] ),
    .B(_2139_),
    .CO(_2140_),
    .S(_2141_));
 HA_X1 _4322_ (.A(_2124_),
    .B(_2002_),
    .CO(_2142_),
    .S(_2143_));
 HA_X1 _4323_ (.A(_2124_),
    .B(\result_exp_stage2[1] ),
    .CO(_2144_),
    .S(_2145_));
 HA_X1 _4324_ (.A(\result_exp_stage2[0] ),
    .B(\result_exp_stage2[1] ),
    .CO(_2146_),
    .S(_2147_));
 HA_X1 _4325_ (.A(_2148_),
    .B(\aligned_b_mant[2] ),
    .CO(_2149_),
    .S(_2150_));
 HA_X1 _4326_ (.A(\aligned_a_mant[2] ),
    .B(_2151_),
    .CO(_2152_),
    .S(_2153_));
 HA_X1 _4327_ (.A(\aligned_a_mant[2] ),
    .B(\aligned_b_mant[2] ),
    .CO(_2154_),
    .S(_2155_));
 HA_X1 _4328_ (.A(_2156_),
    .B(\aligned_b_mant[1] ),
    .CO(_2157_),
    .S(_2158_));
 HA_X1 _4329_ (.A(\aligned_a_mant[1] ),
    .B(_2159_),
    .CO(_2160_),
    .S(_2161_));
 HA_X1 _4330_ (.A(\aligned_a_mant[1] ),
    .B(\aligned_b_mant[1] ),
    .CO(_2162_),
    .S(_2163_));
 HA_X1 _4331_ (.A(_2164_),
    .B(\aligned_b_mant[3] ),
    .CO(_2165_),
    .S(_2166_));
 HA_X1 _4332_ (.A(\aligned_a_mant[3] ),
    .B(_2167_),
    .CO(_2168_),
    .S(_2169_));
 HA_X1 _4333_ (.A(\aligned_a_mant[3] ),
    .B(\aligned_b_mant[3] ),
    .CO(_2170_),
    .S(_2171_));
 HA_X1 _4334_ (.A(_2172_),
    .B(\aligned_b_mant[4] ),
    .CO(_2173_),
    .S(_2174_));
 HA_X1 _4335_ (.A(\aligned_a_mant[4] ),
    .B(_2175_),
    .CO(_2176_),
    .S(_2177_));
 HA_X1 _4336_ (.A(\aligned_a_mant[4] ),
    .B(\aligned_b_mant[4] ),
    .CO(_2178_),
    .S(_2179_));
 HA_X1 _4337_ (.A(_2180_),
    .B(\aligned_b_mant[5] ),
    .CO(_2181_),
    .S(_2182_));
 HA_X1 _4338_ (.A(\aligned_a_mant[5] ),
    .B(_2183_),
    .CO(_2184_),
    .S(_2185_));
 HA_X1 _4339_ (.A(\aligned_a_mant[5] ),
    .B(\aligned_b_mant[5] ),
    .CO(_2186_),
    .S(_2187_));
 HA_X1 _4340_ (.A(_2188_),
    .B(\aligned_b_mant[6] ),
    .CO(_2189_),
    .S(_2190_));
 HA_X1 _4341_ (.A(\aligned_a_mant[6] ),
    .B(_2191_),
    .CO(_2192_),
    .S(_2193_));
 HA_X1 _4342_ (.A(\aligned_a_mant[6] ),
    .B(\aligned_b_mant[6] ),
    .CO(_2194_),
    .S(_2195_));
 HA_X1 _4343_ (.A(_2196_),
    .B(\aligned_b_mant[7] ),
    .CO(_2197_),
    .S(_2198_));
 HA_X1 _4344_ (.A(\aligned_a_mant[7] ),
    .B(_2199_),
    .CO(_2200_),
    .S(_2201_));
 HA_X1 _4345_ (.A(\aligned_a_mant[7] ),
    .B(\aligned_b_mant[7] ),
    .CO(_2202_),
    .S(_2203_));
 HA_X1 _4346_ (.A(_2204_),
    .B(\aligned_b_mant[8] ),
    .CO(_2205_),
    .S(_2206_));
 HA_X1 _4347_ (.A(\aligned_a_mant[8] ),
    .B(_2207_),
    .CO(_2208_),
    .S(_2209_));
 HA_X1 _4348_ (.A(\aligned_a_mant[8] ),
    .B(\aligned_b_mant[8] ),
    .CO(_2210_),
    .S(_2211_));
 HA_X1 _4349_ (.A(_2212_),
    .B(\aligned_b_mant[9] ),
    .CO(_2213_),
    .S(_2214_));
 HA_X1 _4350_ (.A(\aligned_a_mant[9] ),
    .B(_2215_),
    .CO(_2216_),
    .S(_2217_));
 HA_X1 _4351_ (.A(\aligned_a_mant[9] ),
    .B(\aligned_b_mant[9] ),
    .CO(_2218_),
    .S(_2219_));
 HA_X1 _4352_ (.A(_2220_),
    .B(\aligned_b_mant[10] ),
    .CO(_2221_),
    .S(_2222_));
 HA_X1 _4353_ (.A(\aligned_a_mant[10] ),
    .B(_2223_),
    .CO(_2224_),
    .S(_2225_));
 HA_X1 _4354_ (.A(\aligned_a_mant[10] ),
    .B(\aligned_b_mant[10] ),
    .CO(_2226_),
    .S(_2227_));
 HA_X1 _4355_ (.A(_2228_),
    .B(\aligned_b_mant[11] ),
    .CO(_2229_),
    .S(_2230_));
 HA_X1 _4356_ (.A(\aligned_a_mant[11] ),
    .B(_2231_),
    .CO(_2232_),
    .S(_2233_));
 HA_X1 _4357_ (.A(\aligned_a_mant[11] ),
    .B(\aligned_b_mant[11] ),
    .CO(_2234_),
    .S(_2235_));
 HA_X1 _4358_ (.A(_2236_),
    .B(\aligned_b_mant[12] ),
    .CO(_2237_),
    .S(_2238_));
 HA_X1 _4359_ (.A(\aligned_a_mant[12] ),
    .B(_2239_),
    .CO(_2240_),
    .S(_2241_));
 HA_X1 _4360_ (.A(\aligned_a_mant[12] ),
    .B(\aligned_b_mant[12] ),
    .CO(_2242_),
    .S(_2243_));
 HA_X1 _4361_ (.A(_2244_),
    .B(\aligned_b_mant[13] ),
    .CO(_2245_),
    .S(_2246_));
 HA_X1 _4362_ (.A(\aligned_a_mant[13] ),
    .B(_2247_),
    .CO(_2248_),
    .S(_2249_));
 HA_X1 _4363_ (.A(\aligned_a_mant[13] ),
    .B(\aligned_b_mant[13] ),
    .CO(_2250_),
    .S(_2251_));
 HA_X1 _4364_ (.A(_2252_),
    .B(\aligned_b_mant[14] ),
    .CO(_2253_),
    .S(_2254_));
 HA_X1 _4365_ (.A(\aligned_a_mant[14] ),
    .B(_2255_),
    .CO(_2256_),
    .S(_2257_));
 HA_X1 _4366_ (.A(\aligned_a_mant[14] ),
    .B(\aligned_b_mant[14] ),
    .CO(_2258_),
    .S(_2259_));
 HA_X1 _4367_ (.A(_2260_),
    .B(\aligned_b_mant[15] ),
    .CO(_2261_),
    .S(_2262_));
 HA_X1 _4368_ (.A(\aligned_a_mant[15] ),
    .B(_2263_),
    .CO(_2264_),
    .S(_2265_));
 HA_X1 _4369_ (.A(\aligned_a_mant[15] ),
    .B(\aligned_b_mant[15] ),
    .CO(_2266_),
    .S(_2267_));
 HA_X1 _4370_ (.A(_2268_),
    .B(\aligned_b_mant[16] ),
    .CO(_2269_),
    .S(_2270_));
 HA_X1 _4371_ (.A(\aligned_a_mant[16] ),
    .B(_2271_),
    .CO(_2272_),
    .S(_2273_));
 HA_X1 _4372_ (.A(\aligned_a_mant[16] ),
    .B(\aligned_b_mant[16] ),
    .CO(_2274_),
    .S(_2275_));
 HA_X1 _4373_ (.A(_2276_),
    .B(\aligned_b_mant[17] ),
    .CO(_2277_),
    .S(_2278_));
 HA_X1 _4374_ (.A(\aligned_a_mant[17] ),
    .B(_2279_),
    .CO(_2280_),
    .S(_2281_));
 HA_X1 _4375_ (.A(\aligned_a_mant[17] ),
    .B(\aligned_b_mant[17] ),
    .CO(_2282_),
    .S(_2283_));
 HA_X1 _4376_ (.A(_2284_),
    .B(\aligned_b_mant[18] ),
    .CO(_2285_),
    .S(_2286_));
 HA_X1 _4377_ (.A(\aligned_a_mant[18] ),
    .B(_2287_),
    .CO(_2288_),
    .S(_2289_));
 HA_X1 _4378_ (.A(\aligned_a_mant[18] ),
    .B(\aligned_b_mant[18] ),
    .CO(_2290_),
    .S(_2291_));
 HA_X1 _4379_ (.A(_2292_),
    .B(\aligned_b_mant[19] ),
    .CO(_2293_),
    .S(_2294_));
 HA_X1 _4380_ (.A(\aligned_a_mant[19] ),
    .B(_2295_),
    .CO(_2296_),
    .S(_2297_));
 HA_X1 _4381_ (.A(\aligned_a_mant[19] ),
    .B(\aligned_b_mant[19] ),
    .CO(_2298_),
    .S(_2299_));
 HA_X1 _4382_ (.A(_2300_),
    .B(\aligned_b_mant[20] ),
    .CO(_2301_),
    .S(_2302_));
 HA_X1 _4383_ (.A(\aligned_a_mant[20] ),
    .B(_2303_),
    .CO(_2304_),
    .S(_2305_));
 HA_X1 _4384_ (.A(\aligned_a_mant[20] ),
    .B(\aligned_b_mant[20] ),
    .CO(_2306_),
    .S(_2307_));
 HA_X1 _4385_ (.A(_2308_),
    .B(\aligned_b_mant[21] ),
    .CO(_2309_),
    .S(_2310_));
 HA_X1 _4386_ (.A(\aligned_a_mant[21] ),
    .B(_2311_),
    .CO(_2312_),
    .S(_2313_));
 HA_X1 _4387_ (.A(\aligned_a_mant[21] ),
    .B(\aligned_b_mant[21] ),
    .CO(_2314_),
    .S(_2315_));
 HA_X1 _4388_ (.A(_2316_),
    .B(\aligned_b_mant[22] ),
    .CO(_2317_),
    .S(_2318_));
 HA_X1 _4389_ (.A(\aligned_a_mant[22] ),
    .B(_2319_),
    .CO(_2320_),
    .S(_2321_));
 HA_X1 _4390_ (.A(\aligned_a_mant[22] ),
    .B(\aligned_b_mant[22] ),
    .CO(_2322_),
    .S(_2323_));
 HA_X1 _4391_ (.A(_2324_),
    .B(\aligned_b_mant[23] ),
    .CO(_2325_),
    .S(_2326_));
 HA_X1 _4392_ (.A(\aligned_a_mant[23] ),
    .B(_2327_),
    .CO(_2328_),
    .S(_2329_));
 HA_X1 _4393_ (.A(\aligned_a_mant[23] ),
    .B(\aligned_b_mant[23] ),
    .CO(_2330_),
    .S(_2331_));
 HA_X1 _4394_ (.A(_2332_),
    .B(\aligned_b_mant[24] ),
    .CO(_2333_),
    .S(_2334_));
 HA_X1 _4395_ (.A(\aligned_a_mant[24] ),
    .B(_2335_),
    .CO(_2336_),
    .S(_2337_));
 HA_X1 _4396_ (.A(\aligned_a_mant[24] ),
    .B(\aligned_b_mant[24] ),
    .CO(_2338_),
    .S(_2339_));
 HA_X1 _4397_ (.A(_2340_),
    .B(\aligned_b_mant[25] ),
    .CO(_2341_),
    .S(_2342_));
 HA_X1 _4398_ (.A(\aligned_a_mant[25] ),
    .B(_2343_),
    .CO(_2344_),
    .S(_2345_));
 HA_X1 _4399_ (.A(\aligned_a_mant[25] ),
    .B(\aligned_b_mant[25] ),
    .CO(_2346_),
    .S(_2347_));
 DFF_X2 \a_sign_stage1$_SDFF_PN0_  (.D(_0087_),
    .CK(clknet_4_4_0_clk),
    .Q(a_sign_stage1),
    .QN(_1993_));
 DFF_X1 \add_result[10]$_SDFF_PP0_  (.D(_0088_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[10] ),
    .QN(_0008_));
 DFF_X1 \add_result[11]$_SDFF_PP0_  (.D(_0089_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[11] ),
    .QN(_0009_));
 DFF_X2 \add_result[12]$_SDFF_PP0_  (.D(_0090_),
    .CK(clknet_4_9_0_clk),
    .Q(\add_result[12] ),
    .QN(_0010_));
 DFF_X2 \add_result[13]$_SDFF_PP0_  (.D(_0091_),
    .CK(clknet_4_14_0_clk),
    .Q(\add_result[13] ),
    .QN(_0011_));
 DFF_X2 \add_result[14]$_SDFF_PP0_  (.D(_0092_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[14] ),
    .QN(_0012_));
 DFF_X1 \add_result[15]$_SDFF_PP0_  (.D(_0093_),
    .CK(clknet_4_15_0_clk),
    .Q(\add_result[15] ),
    .QN(_0013_));
 DFF_X1 \add_result[16]$_SDFF_PP0_  (.D(_0094_),
    .CK(clknet_4_13_0_clk),
    .Q(\add_result[16] ),
    .QN(_0014_));
 DFF_X2 \add_result[17]$_SDFF_PP0_  (.D(_0095_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[17] ),
    .QN(_0015_));
 DFF_X1 \add_result[18]$_SDFF_PP0_  (.D(_0096_),
    .CK(clknet_4_13_0_clk),
    .Q(\add_result[18] ),
    .QN(_0016_));
 DFF_X1 \add_result[19]$_SDFF_PP0_  (.D(_0097_),
    .CK(clknet_4_13_0_clk),
    .Q(\add_result[19] ),
    .QN(_0017_));
 DFF_X1 \add_result[20]$_SDFF_PP0_  (.D(_0098_),
    .CK(clknet_4_13_0_clk),
    .Q(\add_result[20] ),
    .QN(_0018_));
 DFF_X1 \add_result[21]$_SDFF_PP0_  (.D(_0099_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[21] ),
    .QN(_0019_));
 DFF_X2 \add_result[22]$_SDFF_PP0_  (.D(_0100_),
    .CK(clknet_4_7_0_clk),
    .Q(\add_result[22] ),
    .QN(_0023_));
 DFF_X2 \add_result[23]$_SDFF_PP0_  (.D(_0101_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[23] ),
    .QN(_0022_));
 DFF_X2 \add_result[24]$_SDFF_PP0_  (.D(_0102_),
    .CK(clknet_4_7_0_clk),
    .Q(\add_result[24] ),
    .QN(_0021_));
 DFF_X1 \add_result[25]$_SDFF_PN0_  (.D(_0103_),
    .CK(clknet_4_7_0_clk),
    .Q(\add_result[25] ),
    .QN(_1992_));
 DFF_X1 \add_result[26]$_SDFF_PP0_  (.D(_0104_),
    .CK(clknet_4_7_0_clk),
    .Q(\add_result[26] ),
    .QN(_0020_));
 DFF_X1 \add_result[2]$_SDFF_PP0_  (.D(_0105_),
    .CK(clknet_4_11_0_clk),
    .Q(\add_result[2] ),
    .QN(_0000_));
 DFF_X1 \add_result[3]$_SDFF_PP0_  (.D(_0106_),
    .CK(clknet_4_9_0_clk),
    .Q(\add_result[3] ),
    .QN(_0001_));
 DFF_X1 \add_result[4]$_SDFF_PP0_  (.D(_0107_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[4] ),
    .QN(_0002_));
 DFF_X1 \add_result[5]$_SDFF_PP0_  (.D(_0108_),
    .CK(clknet_4_11_0_clk),
    .Q(\add_result[5] ),
    .QN(_0003_));
 DFF_X1 \add_result[6]$_SDFF_PP0_  (.D(_0109_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[6] ),
    .QN(_0004_));
 DFF_X2 \add_result[7]$_SDFF_PP0_  (.D(_0110_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[7] ),
    .QN(_0005_));
 DFF_X2 \add_result[8]$_SDFF_PP0_  (.D(_0111_),
    .CK(clknet_4_12_0_clk),
    .Q(\add_result[8] ),
    .QN(_0006_));
 DFF_X2 \add_result[9]$_SDFF_PP0_  (.D(_0112_),
    .CK(clknet_4_9_0_clk),
    .Q(\add_result[9] ),
    .QN(_0007_));
 DFF_X1 \aligned_a_mant[0]$_SDFF_PP0_  (.D(_0113_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[0] ),
    .QN(_1991_));
 DFF_X1 \aligned_a_mant[10]$_SDFF_PP0_  (.D(_0114_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[10] ),
    .QN(_2220_));
 DFF_X1 \aligned_a_mant[11]$_SDFF_PP0_  (.D(_0115_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[11] ),
    .QN(_2228_));
 DFF_X1 \aligned_a_mant[12]$_SDFF_PP0_  (.D(_0116_),
    .CK(clknet_4_10_0_clk),
    .Q(\aligned_a_mant[12] ),
    .QN(_2236_));
 DFF_X1 \aligned_a_mant[13]$_SDFF_PP0_  (.D(_0117_),
    .CK(clknet_4_9_0_clk),
    .Q(\aligned_a_mant[13] ),
    .QN(_2244_));
 DFF_X1 \aligned_a_mant[14]$_SDFF_PP0_  (.D(_0118_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[14] ),
    .QN(_2252_));
 DFF_X1 \aligned_a_mant[15]$_SDFF_PP0_  (.D(_0119_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[15] ),
    .QN(_2260_));
 DFF_X1 \aligned_a_mant[16]$_SDFF_PP0_  (.D(_0120_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[16] ),
    .QN(_2268_));
 DFF_X1 \aligned_a_mant[17]$_SDFF_PP0_  (.D(_0121_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_a_mant[17] ),
    .QN(_2276_));
 DFF_X1 \aligned_a_mant[18]$_SDFF_PP0_  (.D(_0122_),
    .CK(clknet_4_3_0_clk),
    .Q(\aligned_a_mant[18] ),
    .QN(_2284_));
 DFF_X1 \aligned_a_mant[19]$_SDFF_PP0_  (.D(_0123_),
    .CK(clknet_4_3_0_clk),
    .Q(\aligned_a_mant[19] ),
    .QN(_2292_));
 DFF_X1 \aligned_a_mant[1]$_SDFF_PP0_  (.D(_0124_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[1] ),
    .QN(_2156_));
 DFF_X1 \aligned_a_mant[20]$_SDFF_PP0_  (.D(_0125_),
    .CK(clknet_4_3_0_clk),
    .Q(\aligned_a_mant[20] ),
    .QN(_2300_));
 DFF_X1 \aligned_a_mant[21]$_SDFF_PP0_  (.D(_0126_),
    .CK(clknet_4_2_0_clk),
    .Q(\aligned_a_mant[21] ),
    .QN(_2308_));
 DFF_X1 \aligned_a_mant[22]$_SDFF_PP0_  (.D(_0127_),
    .CK(clknet_4_3_0_clk),
    .Q(\aligned_a_mant[22] ),
    .QN(_2316_));
 DFF_X1 \aligned_a_mant[23]$_SDFF_PP0_  (.D(_0128_),
    .CK(clknet_4_2_0_clk),
    .Q(\aligned_a_mant[23] ),
    .QN(_2324_));
 DFF_X1 \aligned_a_mant[24]$_SDFF_PP0_  (.D(_0129_),
    .CK(clknet_4_2_0_clk),
    .Q(\aligned_a_mant[24] ),
    .QN(_2332_));
 DFF_X1 \aligned_a_mant[25]$_SDFF_PP0_  (.D(_0130_),
    .CK(clknet_4_6_0_clk),
    .Q(\aligned_a_mant[25] ),
    .QN(_2340_));
 DFF_X1 \aligned_a_mant[2]$_SDFF_PP0_  (.D(_0131_),
    .CK(clknet_4_10_0_clk),
    .Q(\aligned_a_mant[2] ),
    .QN(_2148_));
 DFF_X1 \aligned_a_mant[3]$_SDFF_PP0_  (.D(_0132_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[3] ),
    .QN(_2164_));
 DFF_X1 \aligned_a_mant[4]$_SDFF_PP0_  (.D(_0133_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[4] ),
    .QN(_2172_));
 DFF_X1 \aligned_a_mant[5]$_SDFF_PP0_  (.D(_0134_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[5] ),
    .QN(_2180_));
 DFF_X1 \aligned_a_mant[6]$_SDFF_PP0_  (.D(_0135_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[6] ),
    .QN(_2188_));
 DFF_X1 \aligned_a_mant[7]$_SDFF_PP0_  (.D(_0136_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_a_mant[7] ),
    .QN(_2196_));
 DFF_X1 \aligned_a_mant[8]$_SDFF_PP0_  (.D(_0137_),
    .CK(clknet_4_10_0_clk),
    .Q(\aligned_a_mant[8] ),
    .QN(_2204_));
 DFF_X1 \aligned_a_mant[9]$_SDFF_PP0_  (.D(_0138_),
    .CK(clknet_4_10_0_clk),
    .Q(\aligned_a_mant[9] ),
    .QN(_2212_));
 DFF_X1 \aligned_b_mant[0]$_SDFF_PP0_  (.D(_0139_),
    .CK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[0] ),
    .QN(_1990_));
 DFF_X1 \aligned_b_mant[10]$_SDFF_PN0_  (.D(_0140_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[10] ),
    .QN(_2223_));
 DFF_X1 \aligned_b_mant[11]$_SDFF_PN0_  (.D(_0141_),
    .CK(clknet_4_9_0_clk),
    .Q(\aligned_b_mant[11] ),
    .QN(_2231_));
 DFF_X1 \aligned_b_mant[12]$_SDFF_PN0_  (.D(_0142_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[12] ),
    .QN(_2239_));
 DFF_X1 \aligned_b_mant[13]$_SDFF_PN0_  (.D(_0143_),
    .CK(clknet_4_9_0_clk),
    .Q(\aligned_b_mant[13] ),
    .QN(_2247_));
 DFF_X1 \aligned_b_mant[14]$_SDFF_PN0_  (.D(_0144_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[14] ),
    .QN(_2255_));
 DFF_X1 \aligned_b_mant[15]$_SDFF_PN0_  (.D(_0145_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[15] ),
    .QN(_2263_));
 DFF_X1 \aligned_b_mant[16]$_SDFF_PN0_  (.D(_0146_),
    .CK(clknet_4_8_0_clk),
    .Q(\aligned_b_mant[16] ),
    .QN(_2271_));
 DFF_X1 \aligned_b_mant[17]$_SDFF_PN0_  (.D(_0147_),
    .CK(clknet_4_3_0_clk),
    .Q(\aligned_b_mant[17] ),
    .QN(_2279_));
 DFF_X1 \aligned_b_mant[18]$_SDFF_PN0_  (.D(_0148_),
    .CK(clknet_4_3_0_clk),
    .Q(\aligned_b_mant[18] ),
    .QN(_2287_));
 DFF_X1 \aligned_b_mant[19]$_SDFF_PN0_  (.D(_0149_),
    .CK(clknet_4_3_0_clk),
    .Q(\aligned_b_mant[19] ),
    .QN(_2295_));
 DFF_X2 \aligned_b_mant[1]$_SDFF_PP0_  (.D(_0150_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_b_mant[1] ),
    .QN(_2159_));
 DFF_X1 \aligned_b_mant[20]$_SDFF_PN0_  (.D(_0151_),
    .CK(clknet_4_3_0_clk),
    .Q(\aligned_b_mant[20] ),
    .QN(_2303_));
 DFF_X1 \aligned_b_mant[21]$_SDFF_PN0_  (.D(_0152_),
    .CK(clknet_4_3_0_clk),
    .Q(\aligned_b_mant[21] ),
    .QN(_2311_));
 DFF_X1 \aligned_b_mant[22]$_SDFF_PN0_  (.D(_0153_),
    .CK(clknet_4_2_0_clk),
    .Q(\aligned_b_mant[22] ),
    .QN(_2319_));
 DFF_X1 \aligned_b_mant[23]$_SDFF_PN0_  (.D(_0154_),
    .CK(clknet_4_2_0_clk),
    .Q(\aligned_b_mant[23] ),
    .QN(_2327_));
 DFF_X1 \aligned_b_mant[24]$_SDFF_PN0_  (.D(_0155_),
    .CK(clknet_4_2_0_clk),
    .Q(\aligned_b_mant[24] ),
    .QN(_2335_));
 DFF_X1 \aligned_b_mant[25]$_SDFF_PN0_  (.D(_0156_),
    .CK(clknet_4_6_0_clk),
    .Q(\aligned_b_mant[25] ),
    .QN(_2343_));
 DFF_X1 \aligned_b_mant[2]$_SDFF_PN0_  (.D(_0157_),
    .CK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[2] ),
    .QN(_2151_));
 DFF_X1 \aligned_b_mant[3]$_SDFF_PN0_  (.D(_0158_),
    .CK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[3] ),
    .QN(_2167_));
 DFF_X1 \aligned_b_mant[4]$_SDFF_PN0_  (.D(_0159_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_b_mant[4] ),
    .QN(_2175_));
 DFF_X1 \aligned_b_mant[5]$_SDFF_PN0_  (.D(_0160_),
    .CK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[5] ),
    .QN(_2183_));
 DFF_X1 \aligned_b_mant[6]$_SDFF_PN0_  (.D(_0161_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_b_mant[6] ),
    .QN(_2191_));
 DFF_X1 \aligned_b_mant[7]$_SDFF_PN0_  (.D(_0162_),
    .CK(clknet_4_10_0_clk),
    .Q(\aligned_b_mant[7] ),
    .QN(_2199_));
 DFF_X1 \aligned_b_mant[8]$_SDFF_PN0_  (.D(_0163_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_b_mant[8] ),
    .QN(_2207_));
 DFF_X1 \aligned_b_mant[9]$_SDFF_PN0_  (.D(_0164_),
    .CK(clknet_4_11_0_clk),
    .Q(\aligned_b_mant[9] ),
    .QN(_2215_));
 DFF_X2 \b_sign_stage1$_SDFF_PN0_  (.D(_0165_),
    .CK(clknet_4_4_0_clk),
    .Q(b_sign_stage1),
    .QN(_1989_));
 DFF_X1 \final_exp[0]$_DFFE_PP_  (.D(_0166_),
    .CK(clknet_4_4_0_clk),
    .Q(\final_exp[0] ),
    .QN(_1988_));
 DFF_X1 \final_exp[1]$_DFFE_PP_  (.D(_0167_),
    .CK(clknet_4_5_0_clk),
    .Q(\final_exp[1] ),
    .QN(_1987_));
 DFF_X1 \final_exp[2]$_DFFE_PP_  (.D(_0168_),
    .CK(clknet_4_4_0_clk),
    .Q(\final_exp[2] ),
    .QN(_1986_));
 DFF_X1 \final_exp[3]$_DFFE_PP_  (.D(_0169_),
    .CK(clknet_4_1_0_clk),
    .Q(\final_exp[3] ),
    .QN(_1985_));
 DFF_X1 \final_exp[4]$_DFFE_PP_  (.D(_0170_),
    .CK(clknet_4_4_0_clk),
    .Q(\final_exp[4] ),
    .QN(_1984_));
 DFF_X1 \final_exp[5]$_DFFE_PP_  (.D(_0171_),
    .CK(clknet_4_4_0_clk),
    .Q(\final_exp[5] ),
    .QN(_1983_));
 DFF_X1 \final_exp[6]$_DFFE_PP_  (.D(_0172_),
    .CK(clknet_4_5_0_clk),
    .Q(\final_exp[6] ),
    .QN(_1982_));
 DFF_X1 \final_exp[7]$_DFFE_PP_  (.D(_0173_),
    .CK(clknet_4_5_0_clk),
    .Q(\final_exp[7] ),
    .QN(_1981_));
 DFF_X1 \final_mant[0]$_DFFE_PP_  (.D(_0174_),
    .CK(clknet_4_15_0_clk),
    .Q(\final_mant[0] ),
    .QN(_1980_));
 DFF_X1 \final_mant[10]$_DFFE_PP_  (.D(_0175_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[10] ),
    .QN(_1979_));
 DFF_X1 \final_mant[11]$_DFFE_PP_  (.D(_0176_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[11] ),
    .QN(_1978_));
 DFF_X1 \final_mant[12]$_DFFE_PP_  (.D(_0177_),
    .CK(clknet_4_15_0_clk),
    .Q(\final_mant[12] ),
    .QN(_1977_));
 DFF_X1 \final_mant[13]$_DFFE_PP_  (.D(_0178_),
    .CK(clknet_4_15_0_clk),
    .Q(\final_mant[13] ),
    .QN(_1976_));
 DFF_X1 \final_mant[14]$_DFFE_PP_  (.D(_0179_),
    .CK(clknet_4_15_0_clk),
    .Q(\final_mant[14] ),
    .QN(_1975_));
 DFF_X1 \final_mant[15]$_DFFE_PP_  (.D(_0180_),
    .CK(clknet_4_15_0_clk),
    .Q(\final_mant[15] ),
    .QN(_1974_));
 DFF_X1 \final_mant[16]$_DFFE_PP_  (.D(_0181_),
    .CK(clknet_4_13_0_clk),
    .Q(\final_mant[16] ),
    .QN(_1973_));
 DFF_X1 \final_mant[17]$_DFFE_PP_  (.D(_0182_),
    .CK(clknet_4_13_0_clk),
    .Q(\final_mant[17] ),
    .QN(_1972_));
 DFF_X1 \final_mant[18]$_DFFE_PP_  (.D(_0183_),
    .CK(clknet_4_13_0_clk),
    .Q(\final_mant[18] ),
    .QN(_1971_));
 DFF_X1 \final_mant[19]$_DFFE_PP_  (.D(_0184_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[19] ),
    .QN(_1970_));
 DFF_X1 \final_mant[1]$_DFFE_PP_  (.D(_0185_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[1] ),
    .QN(_1969_));
 DFF_X1 \final_mant[20]$_DFFE_PP_  (.D(_0186_),
    .CK(clknet_4_13_0_clk),
    .Q(\final_mant[20] ),
    .QN(_1968_));
 DFF_X1 \final_mant[21]$_DFFE_PP_  (.D(_0187_),
    .CK(clknet_4_7_0_clk),
    .Q(\final_mant[21] ),
    .QN(_1967_));
 DFF_X1 \final_mant[22]$_DFFE_PP_  (.D(_0188_),
    .CK(clknet_4_13_0_clk),
    .Q(\final_mant[22] ),
    .QN(_1966_));
 DFF_X1 \final_mant[2]$_DFFE_PP_  (.D(_0189_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[2] ),
    .QN(_1965_));
 DFF_X1 \final_mant[3]$_DFFE_PP_  (.D(_0190_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[3] ),
    .QN(_1964_));
 DFF_X1 \final_mant[4]$_DFFE_PP_  (.D(_0191_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[4] ),
    .QN(_1963_));
 DFF_X1 \final_mant[5]$_DFFE_PP_  (.D(_0192_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[5] ),
    .QN(_1962_));
 DFF_X1 \final_mant[6]$_DFFE_PP_  (.D(_0193_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[6] ),
    .QN(_1961_));
 DFF_X1 \final_mant[7]$_DFFE_PP_  (.D(_0025_),
    .CK(clknet_4_12_0_clk),
    .Q(\final_mant[7] ),
    .QN(_1960_));
 DFF_X1 \final_mant[8]$_DFFE_PP_  (.D(_0026_),
    .CK(clknet_4_0_0_clk),
    .Q(\final_mant[8] ),
    .QN(_1959_));
 DFF_X1 \final_mant[9]$_DFFE_PP_  (.D(_0027_),
    .CK(clknet_4_14_0_clk),
    .Q(\final_mant[9] ),
    .QN(_1958_));
 DFF_X1 \inexact$_SDFF_PN0_  (.D(_0028_),
    .CK(clknet_4_13_0_clk),
    .Q(net54),
    .QN(_1957_));
 DFF_X1 \inexact_stage2$_SDFF_PN0_  (.D(_0029_),
    .CK(clknet_4_14_0_clk),
    .Q(inexact_stage2),
    .QN(_1956_));
 DFF_X1 \invalid_op$_SDFF_PN0_  (.D(_0030_),
    .CK(clknet_4_1_0_clk),
    .Q(net55),
    .QN(_1955_));
 DFF_X1 \invalid_op_stage2$_SDFFE_PN0P_  (.D(_0031_),
    .CK(clknet_4_2_0_clk),
    .Q(invalid_op_stage2),
    .QN(_1954_));
 DFF_X1 \is_a_larger_stage1$_SDFF_PN0_  (.D(_0032_),
    .CK(clknet_4_10_0_clk),
    .Q(is_a_larger_stage1),
    .QN(_1953_));
 DFF_X1 \larger_exp_stage1[0]$_SDFF_PN0_  (.D(_0033_),
    .CK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[0] ),
    .QN(_1952_));
 DFF_X1 \larger_exp_stage1[1]$_SDFF_PN0_  (.D(_0034_),
    .CK(clknet_4_6_0_clk),
    .Q(\larger_exp_stage1[1] ),
    .QN(_1951_));
 DFF_X1 \larger_exp_stage1[2]$_SDFF_PN0_  (.D(_0035_),
    .CK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[2] ),
    .QN(_1950_));
 DFF_X1 \larger_exp_stage1[3]$_SDFF_PN0_  (.D(_0036_),
    .CK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[3] ),
    .QN(_1949_));
 DFF_X1 \larger_exp_stage1[4]$_SDFF_PN0_  (.D(_0037_),
    .CK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[4] ),
    .QN(_1948_));
 DFF_X1 \larger_exp_stage1[5]$_SDFF_PN0_  (.D(_0038_),
    .CK(clknet_4_1_0_clk),
    .Q(\larger_exp_stage1[5] ),
    .QN(_1947_));
 DFF_X1 \larger_exp_stage1[6]$_SDFF_PN0_  (.D(_0039_),
    .CK(clknet_4_1_0_clk),
    .Q(\larger_exp_stage1[6] ),
    .QN(_1946_));
 DFF_X1 \larger_exp_stage1[7]$_SDFF_PN0_  (.D(_0040_),
    .CK(clknet_4_0_0_clk),
    .Q(\larger_exp_stage1[7] ),
    .QN(_1945_));
 DFF_X1 \overflow$_SDFF_PN0_  (.D(_0041_),
    .CK(clknet_4_5_0_clk),
    .Q(net56),
    .QN(_1944_));
 DFF_X1 \result[0]$_SDFF_PN0_  (.D(_0042_),
    .CK(clknet_4_15_0_clk),
    .Q(net57),
    .QN(_1943_));
 DFF_X1 \result[10]$_SDFF_PN0_  (.D(_0043_),
    .CK(clknet_4_15_0_clk),
    .Q(net58),
    .QN(_1942_));
 DFF_X1 \result[11]$_SDFF_PN0_  (.D(_0044_),
    .CK(clknet_4_15_0_clk),
    .Q(net59),
    .QN(_1941_));
 DFF_X1 \result[12]$_SDFF_PN0_  (.D(_0045_),
    .CK(clknet_4_15_0_clk),
    .Q(net60),
    .QN(_1940_));
 DFF_X1 \result[13]$_SDFF_PN0_  (.D(_0046_),
    .CK(clknet_4_15_0_clk),
    .Q(net61),
    .QN(_1939_));
 DFF_X1 \result[14]$_SDFF_PN0_  (.D(_0047_),
    .CK(clknet_4_15_0_clk),
    .Q(net62),
    .QN(_1938_));
 DFF_X1 \result[15]$_SDFF_PN0_  (.D(_0048_),
    .CK(clknet_4_15_0_clk),
    .Q(net63),
    .QN(_1937_));
 DFF_X1 \result[16]$_SDFF_PN0_  (.D(_0049_),
    .CK(clknet_4_13_0_clk),
    .Q(net64),
    .QN(_1936_));
 DFF_X1 \result[17]$_SDFF_PN0_  (.D(_0050_),
    .CK(clknet_4_13_0_clk),
    .Q(net65),
    .QN(_1935_));
 DFF_X1 \result[18]$_SDFF_PN0_  (.D(_0051_),
    .CK(clknet_4_13_0_clk),
    .Q(net66),
    .QN(_1934_));
 DFF_X1 \result[19]$_SDFF_PN0_  (.D(_0052_),
    .CK(clknet_4_15_0_clk),
    .Q(net67),
    .QN(_1933_));
 DFF_X1 \result[1]$_SDFF_PN0_  (.D(_0053_),
    .CK(clknet_4_15_0_clk),
    .Q(net68),
    .QN(_1932_));
 DFF_X1 \result[20]$_SDFF_PN0_  (.D(_0054_),
    .CK(clknet_4_13_0_clk),
    .Q(net69),
    .QN(_1931_));
 DFF_X1 \result[21]$_SDFF_PN0_  (.D(_0055_),
    .CK(clknet_4_13_0_clk),
    .Q(net70),
    .QN(_1930_));
 DFF_X1 \result[22]$_SDFF_PN0_  (.D(_0056_),
    .CK(clknet_4_15_0_clk),
    .Q(net71),
    .QN(_1929_));
 DFF_X1 \result[23]$_SDFF_PN0_  (.D(_0057_),
    .CK(clknet_4_1_0_clk),
    .Q(net72),
    .QN(_1928_));
 DFF_X1 \result[24]$_SDFF_PN0_  (.D(_0058_),
    .CK(clknet_4_5_0_clk),
    .Q(net73),
    .QN(_1927_));
 DFF_X1 \result[25]$_SDFF_PN0_  (.D(_0059_),
    .CK(clknet_4_1_0_clk),
    .Q(net74),
    .QN(_1926_));
 DFF_X1 \result[26]$_SDFF_PN0_  (.D(_0060_),
    .CK(clknet_4_1_0_clk),
    .Q(net75),
    .QN(_1925_));
 DFF_X1 \result[27]$_SDFF_PN0_  (.D(_0061_),
    .CK(clknet_4_1_0_clk),
    .Q(net76),
    .QN(_1924_));
 DFF_X1 \result[28]$_SDFF_PN0_  (.D(_0062_),
    .CK(clknet_4_1_0_clk),
    .Q(net77),
    .QN(_1923_));
 DFF_X1 \result[29]$_SDFF_PN0_  (.D(_0063_),
    .CK(clknet_4_5_0_clk),
    .Q(net78),
    .QN(_1922_));
 DFF_X1 \result[2]$_SDFF_PN0_  (.D(_0064_),
    .CK(clknet_4_15_0_clk),
    .Q(net79),
    .QN(_1921_));
 DFF_X1 \result[30]$_SDFF_PN0_  (.D(_0065_),
    .CK(clknet_4_5_0_clk),
    .Q(net80),
    .QN(_1920_));
 DFF_X1 \result[31]$_SDFF_PN0_  (.D(_0066_),
    .CK(clknet_4_1_0_clk),
    .Q(net81),
    .QN(_1919_));
 DFF_X1 \result[3]$_SDFF_PN0_  (.D(_0067_),
    .CK(clknet_4_14_0_clk),
    .Q(net82),
    .QN(_1918_));
 DFF_X1 \result[4]$_SDFF_PN0_  (.D(_0068_),
    .CK(clknet_4_15_0_clk),
    .Q(net83),
    .QN(_1917_));
 DFF_X1 \result[5]$_SDFF_PN0_  (.D(_0069_),
    .CK(clknet_4_14_0_clk),
    .Q(net84),
    .QN(_1916_));
 DFF_X1 \result[6]$_SDFF_PN0_  (.D(_0070_),
    .CK(clknet_4_15_0_clk),
    .Q(net85),
    .QN(_1915_));
 DFF_X1 \result[7]$_SDFF_PN0_  (.D(_0071_),
    .CK(clknet_4_7_0_clk),
    .Q(net86),
    .QN(_1914_));
 DFF_X1 \result[8]$_SDFF_PN0_  (.D(_0072_),
    .CK(clknet_4_0_0_clk),
    .Q(net87),
    .QN(_1913_));
 DFF_X1 \result[9]$_SDFF_PN0_  (.D(_0073_),
    .CK(clknet_4_15_0_clk),
    .Q(net88),
    .QN(_1912_));
 DFF_X2 \result_exp_stage2[0]$_SDFF_PN0_  (.D(_0074_),
    .CK(clknet_4_6_0_clk),
    .Q(\result_exp_stage2[0] ),
    .QN(_2124_));
 DFF_X2 \result_exp_stage2[1]$_SDFF_PN0_  (.D(_0075_),
    .CK(clknet_4_6_0_clk),
    .Q(\result_exp_stage2[1] ),
    .QN(_2002_));
 DFF_X2 \result_exp_stage2[2]$_SDFF_PN0_  (.D(_0076_),
    .CK(clknet_4_4_0_clk),
    .Q(\result_exp_stage2[2] ),
    .QN(_2135_));
 DFF_X1 \result_exp_stage2[3]$_SDFF_PN0_  (.D(_0077_),
    .CK(clknet_4_4_0_clk),
    .Q(\result_exp_stage2[3] ),
    .QN(_0024_));
 DFF_X1 \result_exp_stage2[4]$_SDFF_PN0_  (.D(_0078_),
    .CK(clknet_4_0_0_clk),
    .Q(\result_exp_stage2[4] ),
    .QN(_1911_));
 DFF_X1 \result_exp_stage2[5]$_SDFF_PN0_  (.D(_0079_),
    .CK(clknet_4_1_0_clk),
    .Q(\result_exp_stage2[5] ),
    .QN(_1910_));
 DFF_X1 \result_exp_stage2[6]$_SDFF_PN0_  (.D(_0080_),
    .CK(clknet_4_0_0_clk),
    .Q(\result_exp_stage2[6] ),
    .QN(_1909_));
 DFF_X1 \result_exp_stage2[7]$_SDFF_PN0_  (.D(_0081_),
    .CK(clknet_4_4_0_clk),
    .Q(\result_exp_stage2[7] ),
    .QN(_1908_));
 DFF_X1 \result_sign_stage2$_SDFF_PP0_  (.D(_0082_),
    .CK(clknet_4_1_0_clk),
    .Q(result_sign_stage2),
    .QN(_1907_));
 DFF_X1 \underflow$_SDFF_PP0_  (.D(_0083_),
    .CK(clknet_4_7_0_clk),
    .Q(net89),
    .QN(_1906_));
 DFF_X1 \valid_out$_SDFF_PN0_  (.D(_0084_),
    .CK(clknet_4_0_0_clk),
    .Q(net90),
    .QN(_1905_));
 DFF_X1 \valid_stage1$_SDFF_PN0_  (.D(_0085_),
    .CK(clknet_4_1_0_clk),
    .Q(valid_stage1),
    .QN(_1904_));
 DFF_X1 \valid_stage2$_SDFF_PN0_  (.D(_0086_),
    .CK(clknet_4_1_0_clk),
    .Q(valid_stage2),
    .QN(_1903_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_113 ();
 BUF_X1 input1 (.A(a[0]),
    .Z(net1));
 BUF_X1 input2 (.A(a[10]),
    .Z(net2));
 BUF_X1 input3 (.A(a[11]),
    .Z(net3));
 BUF_X1 input4 (.A(a[12]),
    .Z(net4));
 BUF_X1 input5 (.A(a[13]),
    .Z(net5));
 BUF_X1 input6 (.A(a[14]),
    .Z(net6));
 BUF_X1 input7 (.A(a[15]),
    .Z(net7));
 BUF_X1 input8 (.A(a[16]),
    .Z(net8));
 CLKBUF_X2 input9 (.A(a[17]),
    .Z(net9));
 CLKBUF_X2 input10 (.A(a[18]),
    .Z(net10));
 BUF_X2 input11 (.A(a[19]),
    .Z(net11));
 BUF_X2 input12 (.A(a[1]),
    .Z(net12));
 BUF_X1 input13 (.A(a[20]),
    .Z(net13));
 BUF_X2 input14 (.A(a[21]),
    .Z(net14));
 BUF_X2 input15 (.A(a[22]),
    .Z(net15));
 BUF_X2 input16 (.A(a[23]),
    .Z(net16));
 BUF_X2 input17 (.A(a[24]),
    .Z(net17));
 BUF_X2 input18 (.A(a[25]),
    .Z(net18));
 BUF_X2 input19 (.A(a[26]),
    .Z(net19));
 CLKBUF_X2 input20 (.A(a[27]),
    .Z(net20));
 CLKBUF_X2 input21 (.A(a[28]),
    .Z(net21));
 CLKBUF_X2 input22 (.A(a[29]),
    .Z(net22));
 BUF_X2 input23 (.A(a[2]),
    .Z(net23));
 CLKBUF_X2 input24 (.A(a[30]),
    .Z(net24));
 BUF_X1 input25 (.A(a[31]),
    .Z(net25));
 BUF_X2 input26 (.A(a[3]),
    .Z(net26));
 BUF_X1 input27 (.A(a[4]),
    .Z(net27));
 CLKBUF_X2 input28 (.A(a[5]),
    .Z(net28));
 BUF_X2 input29 (.A(a[6]),
    .Z(net29));
 BUF_X1 input30 (.A(a[7]),
    .Z(net30));
 BUF_X1 input31 (.A(a[8]),
    .Z(net31));
 BUF_X1 input32 (.A(a[9]),
    .Z(net32));
 BUF_X2 input33 (.A(b[0]),
    .Z(net33));
 BUF_X1 input34 (.A(b[10]),
    .Z(net34));
 BUF_X1 input35 (.A(b[11]),
    .Z(net35));
 BUF_X1 input36 (.A(b[12]),
    .Z(net36));
 BUF_X1 input37 (.A(b[15]),
    .Z(net37));
 BUF_X2 input38 (.A(b[1]),
    .Z(net38));
 CLKBUF_X2 input39 (.A(b[20]),
    .Z(net39));
 BUF_X2 input40 (.A(b[23]),
    .Z(net40));
 BUF_X2 input41 (.A(b[24]),
    .Z(net41));
 BUF_X2 input42 (.A(b[25]),
    .Z(net42));
 BUF_X2 input43 (.A(b[26]),
    .Z(net43));
 BUF_X2 input44 (.A(b[27]),
    .Z(net44));
 BUF_X2 input45 (.A(b[28]),
    .Z(net45));
 BUF_X2 input46 (.A(b[29]),
    .Z(net46));
 BUF_X1 input47 (.A(b[2]),
    .Z(net47));
 BUF_X2 input48 (.A(b[30]),
    .Z(net48));
 BUF_X1 input49 (.A(b[31]),
    .Z(net49));
 CLKBUF_X2 input50 (.A(b[3]),
    .Z(net50));
 BUF_X1 input51 (.A(b[4]),
    .Z(net51));
 BUF_X1 input52 (.A(b[5]),
    .Z(net52));
 BUF_X1 input53 (.A(valid_in),
    .Z(net53));
 BUF_X1 output54 (.A(net54),
    .Z(inexact));
 BUF_X1 output55 (.A(net55),
    .Z(invalid_op));
 BUF_X1 output56 (.A(net56),
    .Z(overflow));
 BUF_X1 output57 (.A(net57),
    .Z(result[0]));
 BUF_X1 output58 (.A(net58),
    .Z(result[10]));
 BUF_X1 output59 (.A(net59),
    .Z(result[11]));
 BUF_X1 output60 (.A(net60),
    .Z(result[12]));
 BUF_X1 output61 (.A(net61),
    .Z(result[13]));
 BUF_X1 output62 (.A(net62),
    .Z(result[14]));
 BUF_X1 output63 (.A(net63),
    .Z(result[15]));
 BUF_X1 output64 (.A(net64),
    .Z(result[16]));
 BUF_X1 output65 (.A(net65),
    .Z(result[17]));
 BUF_X1 output66 (.A(net66),
    .Z(result[18]));
 BUF_X1 output67 (.A(net67),
    .Z(result[19]));
 BUF_X1 output68 (.A(net68),
    .Z(result[1]));
 BUF_X1 output69 (.A(net69),
    .Z(result[20]));
 BUF_X1 output70 (.A(net70),
    .Z(result[21]));
 BUF_X1 output71 (.A(net71),
    .Z(result[22]));
 BUF_X1 output72 (.A(net72),
    .Z(result[23]));
 BUF_X1 output73 (.A(net73),
    .Z(result[24]));
 BUF_X1 output74 (.A(net74),
    .Z(result[25]));
 BUF_X1 output75 (.A(net75),
    .Z(result[26]));
 BUF_X1 output76 (.A(net76),
    .Z(result[27]));
 BUF_X1 output77 (.A(net77),
    .Z(result[28]));
 BUF_X1 output78 (.A(net78),
    .Z(result[29]));
 BUF_X1 output79 (.A(net79),
    .Z(result[2]));
 BUF_X1 output80 (.A(net80),
    .Z(result[30]));
 BUF_X1 output81 (.A(net81),
    .Z(result[31]));
 BUF_X1 output82 (.A(net82),
    .Z(result[3]));
 BUF_X1 output83 (.A(net83),
    .Z(result[4]));
 BUF_X1 output84 (.A(net84),
    .Z(result[5]));
 BUF_X1 output85 (.A(net85),
    .Z(result[6]));
 BUF_X1 output86 (.A(net86),
    .Z(result[7]));
 BUF_X1 output87 (.A(net87),
    .Z(result[8]));
 BUF_X1 output88 (.A(net88),
    .Z(result[9]));
 BUF_X1 output89 (.A(net89),
    .Z(underflow));
 BUF_X1 output90 (.A(net90),
    .Z(valid_out));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X8 clkload0 (.A(clknet_4_0_0_clk));
 INV_X4 clkload1 (.A(clknet_4_1_0_clk));
 INV_X8 clkload2 (.A(clknet_4_2_0_clk));
 INV_X8 clkload3 (.A(clknet_4_3_0_clk));
 INV_X8 clkload4 (.A(clknet_4_4_0_clk));
 INV_X8 clkload5 (.A(clknet_4_5_0_clk));
 INV_X8 clkload6 (.A(clknet_4_6_0_clk));
 INV_X8 clkload7 (.A(clknet_4_7_0_clk));
 INV_X4 clkload8 (.A(clknet_4_8_0_clk));
 INV_X8 clkload9 (.A(clknet_4_9_0_clk));
 INV_X8 clkload10 (.A(clknet_4_10_0_clk));
 INV_X4 clkload11 (.A(clknet_4_11_0_clk));
 INV_X4 clkload12 (.A(clknet_4_12_0_clk));
 INV_X2 clkload13 (.A(clknet_4_13_0_clk));
 INV_X4 clkload14 (.A(clknet_4_14_0_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X4 FILLER_0_65 ();
 FILLCELL_X2 FILLER_0_69 ();
 FILLCELL_X4 FILLER_0_75 ();
 FILLCELL_X1 FILLER_0_79 ();
 FILLCELL_X1 FILLER_0_104 ();
 FILLCELL_X2 FILLER_0_117 ();
 FILLCELL_X8 FILLER_0_127 ();
 FILLCELL_X4 FILLER_0_135 ();
 FILLCELL_X2 FILLER_0_139 ();
 FILLCELL_X1 FILLER_0_161 ();
 FILLCELL_X2 FILLER_0_165 ();
 FILLCELL_X1 FILLER_0_167 ();
 FILLCELL_X4 FILLER_0_171 ();
 FILLCELL_X2 FILLER_0_175 ();
 FILLCELL_X8 FILLER_0_183 ();
 FILLCELL_X2 FILLER_0_191 ();
 FILLCELL_X32 FILLER_0_222 ();
 FILLCELL_X8 FILLER_0_254 ();
 FILLCELL_X4 FILLER_0_262 ();
 FILLCELL_X2 FILLER_0_266 ();
 FILLCELL_X1 FILLER_0_268 ();
 FILLCELL_X8 FILLER_0_272 ();
 FILLCELL_X1 FILLER_0_280 ();
 FILLCELL_X16 FILLER_0_301 ();
 FILLCELL_X8 FILLER_0_317 ();
 FILLCELL_X2 FILLER_0_325 ();
 FILLCELL_X32 FILLER_0_330 ();
 FILLCELL_X32 FILLER_0_362 ();
 FILLCELL_X32 FILLER_0_394 ();
 FILLCELL_X1 FILLER_0_426 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X4 FILLER_1_65 ();
 FILLCELL_X8 FILLER_1_73 ();
 FILLCELL_X4 FILLER_1_81 ();
 FILLCELL_X1 FILLER_1_85 ();
 FILLCELL_X2 FILLER_1_90 ();
 FILLCELL_X1 FILLER_1_92 ();
 FILLCELL_X2 FILLER_1_109 ();
 FILLCELL_X4 FILLER_1_125 ();
 FILLCELL_X1 FILLER_1_129 ();
 FILLCELL_X4 FILLER_1_151 ();
 FILLCELL_X2 FILLER_1_155 ();
 FILLCELL_X2 FILLER_1_160 ();
 FILLCELL_X8 FILLER_1_183 ();
 FILLCELL_X4 FILLER_1_191 ();
 FILLCELL_X2 FILLER_1_195 ();
 FILLCELL_X16 FILLER_1_239 ();
 FILLCELL_X1 FILLER_1_255 ();
 FILLCELL_X8 FILLER_1_273 ();
 FILLCELL_X2 FILLER_1_298 ();
 FILLCELL_X8 FILLER_1_303 ();
 FILLCELL_X1 FILLER_1_311 ();
 FILLCELL_X32 FILLER_1_329 ();
 FILLCELL_X32 FILLER_1_361 ();
 FILLCELL_X32 FILLER_1_393 ();
 FILLCELL_X2 FILLER_1_425 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X16 FILLER_2_65 ();
 FILLCELL_X2 FILLER_2_81 ();
 FILLCELL_X16 FILLER_2_124 ();
 FILLCELL_X4 FILLER_2_140 ();
 FILLCELL_X1 FILLER_2_144 ();
 FILLCELL_X1 FILLER_2_183 ();
 FILLCELL_X1 FILLER_2_207 ();
 FILLCELL_X2 FILLER_2_211 ();
 FILLCELL_X8 FILLER_2_232 ();
 FILLCELL_X4 FILLER_2_240 ();
 FILLCELL_X2 FILLER_2_244 ();
 FILLCELL_X1 FILLER_2_246 ();
 FILLCELL_X4 FILLER_2_264 ();
 FILLCELL_X16 FILLER_2_293 ();
 FILLCELL_X4 FILLER_2_309 ();
 FILLCELL_X32 FILLER_2_317 ();
 FILLCELL_X32 FILLER_2_349 ();
 FILLCELL_X32 FILLER_2_381 ();
 FILLCELL_X8 FILLER_2_413 ();
 FILLCELL_X4 FILLER_2_421 ();
 FILLCELL_X2 FILLER_2_425 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_65 ();
 FILLCELL_X4 FILLER_3_73 ();
 FILLCELL_X2 FILLER_3_77 ();
 FILLCELL_X32 FILLER_3_103 ();
 FILLCELL_X8 FILLER_3_135 ();
 FILLCELL_X1 FILLER_3_143 ();
 FILLCELL_X16 FILLER_3_168 ();
 FILLCELL_X8 FILLER_3_184 ();
 FILLCELL_X2 FILLER_3_192 ();
 FILLCELL_X8 FILLER_3_211 ();
 FILLCELL_X4 FILLER_3_219 ();
 FILLCELL_X8 FILLER_3_235 ();
 FILLCELL_X4 FILLER_3_243 ();
 FILLCELL_X1 FILLER_3_247 ();
 FILLCELL_X4 FILLER_3_252 ();
 FILLCELL_X4 FILLER_3_282 ();
 FILLCELL_X2 FILLER_3_286 ();
 FILLCELL_X1 FILLER_3_297 ();
 FILLCELL_X32 FILLER_3_315 ();
 FILLCELL_X32 FILLER_3_347 ();
 FILLCELL_X32 FILLER_3_379 ();
 FILLCELL_X16 FILLER_3_411 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X16 FILLER_4_33 ();
 FILLCELL_X1 FILLER_4_49 ();
 FILLCELL_X16 FILLER_4_52 ();
 FILLCELL_X4 FILLER_4_68 ();
 FILLCELL_X1 FILLER_4_72 ();
 FILLCELL_X1 FILLER_4_77 ();
 FILLCELL_X2 FILLER_4_88 ();
 FILLCELL_X8 FILLER_4_106 ();
 FILLCELL_X4 FILLER_4_114 ();
 FILLCELL_X2 FILLER_4_121 ();
 FILLCELL_X1 FILLER_4_123 ();
 FILLCELL_X4 FILLER_4_141 ();
 FILLCELL_X1 FILLER_4_145 ();
 FILLCELL_X1 FILLER_4_150 ();
 FILLCELL_X8 FILLER_4_168 ();
 FILLCELL_X16 FILLER_4_183 ();
 FILLCELL_X1 FILLER_4_199 ();
 FILLCELL_X2 FILLER_4_203 ();
 FILLCELL_X1 FILLER_4_205 ();
 FILLCELL_X2 FILLER_4_229 ();
 FILLCELL_X1 FILLER_4_231 ();
 FILLCELL_X2 FILLER_4_235 ();
 FILLCELL_X1 FILLER_4_237 ();
 FILLCELL_X2 FILLER_4_244 ();
 FILLCELL_X4 FILLER_4_295 ();
 FILLCELL_X2 FILLER_4_299 ();
 FILLCELL_X2 FILLER_4_305 ();
 FILLCELL_X1 FILLER_4_307 ();
 FILLCELL_X16 FILLER_4_313 ();
 FILLCELL_X2 FILLER_4_341 ();
 FILLCELL_X1 FILLER_4_343 ();
 FILLCELL_X1 FILLER_4_357 ();
 FILLCELL_X2 FILLER_4_363 ();
 FILLCELL_X4 FILLER_4_368 ();
 FILLCELL_X2 FILLER_4_372 ();
 FILLCELL_X1 FILLER_4_374 ();
 FILLCELL_X1 FILLER_4_386 ();
 FILLCELL_X32 FILLER_4_392 ();
 FILLCELL_X2 FILLER_4_424 ();
 FILLCELL_X1 FILLER_4_426 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X16 FILLER_5_33 ();
 FILLCELL_X1 FILLER_5_49 ();
 FILLCELL_X8 FILLER_5_57 ();
 FILLCELL_X1 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_85 ();
 FILLCELL_X1 FILLER_5_100 ();
 FILLCELL_X2 FILLER_5_122 ();
 FILLCELL_X1 FILLER_5_127 ();
 FILLCELL_X8 FILLER_5_145 ();
 FILLCELL_X2 FILLER_5_153 ();
 FILLCELL_X8 FILLER_5_176 ();
 FILLCELL_X2 FILLER_5_184 ();
 FILLCELL_X1 FILLER_5_186 ();
 FILLCELL_X4 FILLER_5_213 ();
 FILLCELL_X1 FILLER_5_217 ();
 FILLCELL_X1 FILLER_5_224 ();
 FILLCELL_X1 FILLER_5_228 ();
 FILLCELL_X1 FILLER_5_246 ();
 FILLCELL_X1 FILLER_5_251 ();
 FILLCELL_X1 FILLER_5_275 ();
 FILLCELL_X1 FILLER_5_283 ();
 FILLCELL_X1 FILLER_5_304 ();
 FILLCELL_X1 FILLER_5_308 ();
 FILLCELL_X1 FILLER_5_319 ();
 FILLCELL_X4 FILLER_5_346 ();
 FILLCELL_X2 FILLER_5_350 ();
 FILLCELL_X1 FILLER_5_352 ();
 FILLCELL_X4 FILLER_5_368 ();
 FILLCELL_X2 FILLER_5_389 ();
 FILLCELL_X1 FILLER_5_391 ();
 FILLCELL_X16 FILLER_5_396 ();
 FILLCELL_X8 FILLER_5_412 ();
 FILLCELL_X4 FILLER_5_420 ();
 FILLCELL_X2 FILLER_5_424 ();
 FILLCELL_X1 FILLER_5_426 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X8 FILLER_6_33 ();
 FILLCELL_X4 FILLER_6_41 ();
 FILLCELL_X1 FILLER_6_45 ();
 FILLCELL_X8 FILLER_6_59 ();
 FILLCELL_X4 FILLER_6_67 ();
 FILLCELL_X1 FILLER_6_71 ();
 FILLCELL_X8 FILLER_6_82 ();
 FILLCELL_X4 FILLER_6_90 ();
 FILLCELL_X4 FILLER_6_113 ();
 FILLCELL_X2 FILLER_6_117 ();
 FILLCELL_X1 FILLER_6_119 ();
 FILLCELL_X4 FILLER_6_123 ();
 FILLCELL_X8 FILLER_6_144 ();
 FILLCELL_X2 FILLER_6_152 ();
 FILLCELL_X16 FILLER_6_158 ();
 FILLCELL_X8 FILLER_6_174 ();
 FILLCELL_X8 FILLER_6_202 ();
 FILLCELL_X4 FILLER_6_210 ();
 FILLCELL_X2 FILLER_6_214 ();
 FILLCELL_X2 FILLER_6_218 ();
 FILLCELL_X1 FILLER_6_223 ();
 FILLCELL_X2 FILLER_6_275 ();
 FILLCELL_X1 FILLER_6_302 ();
 FILLCELL_X2 FILLER_6_331 ();
 FILLCELL_X1 FILLER_6_333 ();
 FILLCELL_X4 FILLER_6_355 ();
 FILLCELL_X1 FILLER_6_371 ();
 FILLCELL_X1 FILLER_6_376 ();
 FILLCELL_X2 FILLER_6_380 ();
 FILLCELL_X1 FILLER_6_391 ();
 FILLCELL_X2 FILLER_6_396 ();
 FILLCELL_X1 FILLER_6_402 ();
 FILLCELL_X16 FILLER_6_408 ();
 FILLCELL_X2 FILLER_6_424 ();
 FILLCELL_X1 FILLER_6_426 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X8 FILLER_7_33 ();
 FILLCELL_X4 FILLER_7_41 ();
 FILLCELL_X2 FILLER_7_45 ();
 FILLCELL_X4 FILLER_7_64 ();
 FILLCELL_X2 FILLER_7_68 ();
 FILLCELL_X16 FILLER_7_90 ();
 FILLCELL_X4 FILLER_7_106 ();
 FILLCELL_X2 FILLER_7_110 ();
 FILLCELL_X1 FILLER_7_112 ();
 FILLCELL_X16 FILLER_7_125 ();
 FILLCELL_X8 FILLER_7_141 ();
 FILLCELL_X4 FILLER_7_149 ();
 FILLCELL_X1 FILLER_7_153 ();
 FILLCELL_X2 FILLER_7_171 ();
 FILLCELL_X1 FILLER_7_173 ();
 FILLCELL_X16 FILLER_7_181 ();
 FILLCELL_X2 FILLER_7_197 ();
 FILLCELL_X1 FILLER_7_199 ();
 FILLCELL_X8 FILLER_7_217 ();
 FILLCELL_X2 FILLER_7_225 ();
 FILLCELL_X4 FILLER_7_233 ();
 FILLCELL_X2 FILLER_7_237 ();
 FILLCELL_X2 FILLER_7_315 ();
 FILLCELL_X1 FILLER_7_317 ();
 FILLCELL_X2 FILLER_7_322 ();
 FILLCELL_X4 FILLER_7_341 ();
 FILLCELL_X2 FILLER_7_345 ();
 FILLCELL_X1 FILLER_7_351 ();
 FILLCELL_X4 FILLER_7_370 ();
 FILLCELL_X2 FILLER_7_374 ();
 FILLCELL_X16 FILLER_7_411 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X8 FILLER_8_33 ();
 FILLCELL_X4 FILLER_8_41 ();
 FILLCELL_X2 FILLER_8_45 ();
 FILLCELL_X4 FILLER_8_64 ();
 FILLCELL_X1 FILLER_8_68 ();
 FILLCELL_X1 FILLER_8_82 ();
 FILLCELL_X8 FILLER_8_87 ();
 FILLCELL_X8 FILLER_8_105 ();
 FILLCELL_X4 FILLER_8_113 ();
 FILLCELL_X1 FILLER_8_117 ();
 FILLCELL_X2 FILLER_8_130 ();
 FILLCELL_X8 FILLER_8_149 ();
 FILLCELL_X4 FILLER_8_157 ();
 FILLCELL_X16 FILLER_8_165 ();
 FILLCELL_X4 FILLER_8_217 ();
 FILLCELL_X2 FILLER_8_221 ();
 FILLCELL_X1 FILLER_8_229 ();
 FILLCELL_X2 FILLER_8_296 ();
 FILLCELL_X1 FILLER_8_298 ();
 FILLCELL_X2 FILLER_8_301 ();
 FILLCELL_X2 FILLER_8_313 ();
 FILLCELL_X4 FILLER_8_331 ();
 FILLCELL_X2 FILLER_8_364 ();
 FILLCELL_X2 FILLER_8_384 ();
 FILLCELL_X1 FILLER_8_408 ();
 FILLCELL_X8 FILLER_8_412 ();
 FILLCELL_X4 FILLER_8_420 ();
 FILLCELL_X2 FILLER_8_424 ();
 FILLCELL_X1 FILLER_8_426 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X8 FILLER_9_49 ();
 FILLCELL_X2 FILLER_9_84 ();
 FILLCELL_X4 FILLER_9_90 ();
 FILLCELL_X1 FILLER_9_94 ();
 FILLCELL_X2 FILLER_9_121 ();
 FILLCELL_X1 FILLER_9_123 ();
 FILLCELL_X2 FILLER_9_127 ();
 FILLCELL_X1 FILLER_9_129 ();
 FILLCELL_X16 FILLER_9_147 ();
 FILLCELL_X1 FILLER_9_167 ();
 FILLCELL_X4 FILLER_9_185 ();
 FILLCELL_X4 FILLER_9_206 ();
 FILLCELL_X2 FILLER_9_210 ();
 FILLCELL_X1 FILLER_9_212 ();
 FILLCELL_X1 FILLER_9_227 ();
 FILLCELL_X4 FILLER_9_319 ();
 FILLCELL_X2 FILLER_9_323 ();
 FILLCELL_X1 FILLER_9_325 ();
 FILLCELL_X2 FILLER_9_333 ();
 FILLCELL_X2 FILLER_9_410 ();
 FILLCELL_X8 FILLER_9_415 ();
 FILLCELL_X4 FILLER_9_423 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_33 ();
 FILLCELL_X2 FILLER_10_37 ();
 FILLCELL_X1 FILLER_10_70 ();
 FILLCELL_X8 FILLER_10_85 ();
 FILLCELL_X1 FILLER_10_93 ();
 FILLCELL_X1 FILLER_10_99 ();
 FILLCELL_X4 FILLER_10_110 ();
 FILLCELL_X32 FILLER_10_116 ();
 FILLCELL_X2 FILLER_10_148 ();
 FILLCELL_X1 FILLER_10_150 ();
 FILLCELL_X8 FILLER_10_172 ();
 FILLCELL_X2 FILLER_10_180 ();
 FILLCELL_X8 FILLER_10_192 ();
 FILLCELL_X4 FILLER_10_200 ();
 FILLCELL_X1 FILLER_10_257 ();
 FILLCELL_X1 FILLER_10_296 ();
 FILLCELL_X2 FILLER_10_316 ();
 FILLCELL_X1 FILLER_10_318 ();
 FILLCELL_X1 FILLER_10_334 ();
 FILLCELL_X2 FILLER_10_345 ();
 FILLCELL_X1 FILLER_10_350 ();
 FILLCELL_X2 FILLER_10_382 ();
 FILLCELL_X2 FILLER_10_394 ();
 FILLCELL_X1 FILLER_10_396 ();
 FILLCELL_X8 FILLER_10_415 ();
 FILLCELL_X4 FILLER_10_423 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X8 FILLER_11_33 ();
 FILLCELL_X4 FILLER_11_41 ();
 FILLCELL_X2 FILLER_11_45 ();
 FILLCELL_X2 FILLER_11_59 ();
 FILLCELL_X1 FILLER_11_61 ();
 FILLCELL_X4 FILLER_11_83 ();
 FILLCELL_X1 FILLER_11_87 ();
 FILLCELL_X2 FILLER_11_90 ();
 FILLCELL_X1 FILLER_11_92 ();
 FILLCELL_X1 FILLER_11_98 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X4 FILLER_11_161 ();
 FILLCELL_X2 FILLER_11_182 ();
 FILLCELL_X4 FILLER_11_194 ();
 FILLCELL_X2 FILLER_11_198 ();
 FILLCELL_X8 FILLER_11_204 ();
 FILLCELL_X2 FILLER_11_212 ();
 FILLCELL_X1 FILLER_11_254 ();
 FILLCELL_X4 FILLER_11_276 ();
 FILLCELL_X2 FILLER_11_280 ();
 FILLCELL_X8 FILLER_11_287 ();
 FILLCELL_X1 FILLER_11_295 ();
 FILLCELL_X1 FILLER_11_301 ();
 FILLCELL_X4 FILLER_11_321 ();
 FILLCELL_X1 FILLER_11_325 ();
 FILLCELL_X2 FILLER_11_410 ();
 FILLCELL_X1 FILLER_11_412 ();
 FILLCELL_X4 FILLER_11_420 ();
 FILLCELL_X2 FILLER_11_424 ();
 FILLCELL_X1 FILLER_11_426 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_17 ();
 FILLCELL_X1 FILLER_12_25 ();
 FILLCELL_X2 FILLER_12_44 ();
 FILLCELL_X1 FILLER_12_46 ();
 FILLCELL_X8 FILLER_12_56 ();
 FILLCELL_X2 FILLER_12_64 ();
 FILLCELL_X1 FILLER_12_66 ();
 FILLCELL_X1 FILLER_12_74 ();
 FILLCELL_X1 FILLER_12_79 ();
 FILLCELL_X1 FILLER_12_86 ();
 FILLCELL_X2 FILLER_12_96 ();
 FILLCELL_X4 FILLER_12_112 ();
 FILLCELL_X2 FILLER_12_116 ();
 FILLCELL_X8 FILLER_12_127 ();
 FILLCELL_X2 FILLER_12_135 ();
 FILLCELL_X1 FILLER_12_142 ();
 FILLCELL_X1 FILLER_12_147 ();
 FILLCELL_X2 FILLER_12_155 ();
 FILLCELL_X1 FILLER_12_157 ();
 FILLCELL_X1 FILLER_12_161 ();
 FILLCELL_X1 FILLER_12_166 ();
 FILLCELL_X2 FILLER_12_191 ();
 FILLCELL_X1 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_201 ();
 FILLCELL_X8 FILLER_12_233 ();
 FILLCELL_X4 FILLER_12_241 ();
 FILLCELL_X16 FILLER_12_254 ();
 FILLCELL_X2 FILLER_12_270 ();
 FILLCELL_X2 FILLER_12_295 ();
 FILLCELL_X1 FILLER_12_297 ();
 FILLCELL_X2 FILLER_12_321 ();
 FILLCELL_X2 FILLER_12_330 ();
 FILLCELL_X1 FILLER_12_332 ();
 FILLCELL_X4 FILLER_12_347 ();
 FILLCELL_X1 FILLER_12_351 ();
 FILLCELL_X2 FILLER_12_362 ();
 FILLCELL_X1 FILLER_12_364 ();
 FILLCELL_X8 FILLER_12_382 ();
 FILLCELL_X8 FILLER_12_394 ();
 FILLCELL_X16 FILLER_12_409 ();
 FILLCELL_X2 FILLER_12_425 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X8 FILLER_13_17 ();
 FILLCELL_X1 FILLER_13_25 ();
 FILLCELL_X1 FILLER_13_63 ();
 FILLCELL_X4 FILLER_13_89 ();
 FILLCELL_X2 FILLER_13_107 ();
 FILLCELL_X1 FILLER_13_109 ();
 FILLCELL_X4 FILLER_13_114 ();
 FILLCELL_X1 FILLER_13_118 ();
 FILLCELL_X8 FILLER_13_129 ();
 FILLCELL_X2 FILLER_13_137 ();
 FILLCELL_X1 FILLER_13_148 ();
 FILLCELL_X4 FILLER_13_207 ();
 FILLCELL_X1 FILLER_13_211 ();
 FILLCELL_X1 FILLER_13_231 ();
 FILLCELL_X1 FILLER_13_241 ();
 FILLCELL_X1 FILLER_13_260 ();
 FILLCELL_X4 FILLER_13_263 ();
 FILLCELL_X2 FILLER_13_267 ();
 FILLCELL_X8 FILLER_13_279 ();
 FILLCELL_X2 FILLER_13_287 ();
 FILLCELL_X1 FILLER_13_289 ();
 FILLCELL_X1 FILLER_13_297 ();
 FILLCELL_X2 FILLER_13_313 ();
 FILLCELL_X2 FILLER_13_318 ();
 FILLCELL_X2 FILLER_13_361 ();
 FILLCELL_X2 FILLER_13_374 ();
 FILLCELL_X4 FILLER_13_384 ();
 FILLCELL_X16 FILLER_13_409 ();
 FILLCELL_X2 FILLER_13_425 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_9 ();
 FILLCELL_X16 FILLER_14_14 ();
 FILLCELL_X1 FILLER_14_30 ();
 FILLCELL_X1 FILLER_14_66 ();
 FILLCELL_X2 FILLER_14_80 ();
 FILLCELL_X8 FILLER_14_128 ();
 FILLCELL_X2 FILLER_14_136 ();
 FILLCELL_X1 FILLER_14_138 ();
 FILLCELL_X16 FILLER_14_157 ();
 FILLCELL_X4 FILLER_14_173 ();
 FILLCELL_X4 FILLER_14_186 ();
 FILLCELL_X2 FILLER_14_190 ();
 FILLCELL_X1 FILLER_14_192 ();
 FILLCELL_X16 FILLER_14_212 ();
 FILLCELL_X2 FILLER_14_228 ();
 FILLCELL_X1 FILLER_14_230 ();
 FILLCELL_X2 FILLER_14_241 ();
 FILLCELL_X1 FILLER_14_246 ();
 FILLCELL_X4 FILLER_14_265 ();
 FILLCELL_X1 FILLER_14_269 ();
 FILLCELL_X4 FILLER_14_275 ();
 FILLCELL_X1 FILLER_14_279 ();
 FILLCELL_X4 FILLER_14_290 ();
 FILLCELL_X2 FILLER_14_294 ();
 FILLCELL_X1 FILLER_14_300 ();
 FILLCELL_X1 FILLER_14_305 ();
 FILLCELL_X2 FILLER_14_314 ();
 FILLCELL_X1 FILLER_14_316 ();
 FILLCELL_X2 FILLER_14_321 ();
 FILLCELL_X1 FILLER_14_323 ();
 FILLCELL_X2 FILLER_14_328 ();
 FILLCELL_X4 FILLER_14_335 ();
 FILLCELL_X2 FILLER_14_339 ();
 FILLCELL_X1 FILLER_14_341 ();
 FILLCELL_X1 FILLER_14_352 ();
 FILLCELL_X2 FILLER_14_355 ();
 FILLCELL_X1 FILLER_14_357 ();
 FILLCELL_X1 FILLER_14_384 ();
 FILLCELL_X8 FILLER_14_412 ();
 FILLCELL_X4 FILLER_14_420 ();
 FILLCELL_X2 FILLER_14_424 ();
 FILLCELL_X1 FILLER_14_426 ();
 FILLCELL_X8 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_9 ();
 FILLCELL_X8 FILLER_15_24 ();
 FILLCELL_X1 FILLER_15_32 ();
 FILLCELL_X2 FILLER_15_65 ();
 FILLCELL_X1 FILLER_15_84 ();
 FILLCELL_X1 FILLER_15_89 ();
 FILLCELL_X1 FILLER_15_95 ();
 FILLCELL_X1 FILLER_15_100 ();
 FILLCELL_X1 FILLER_15_119 ();
 FILLCELL_X8 FILLER_15_122 ();
 FILLCELL_X4 FILLER_15_130 ();
 FILLCELL_X2 FILLER_15_134 ();
 FILLCELL_X1 FILLER_15_136 ();
 FILLCELL_X1 FILLER_15_145 ();
 FILLCELL_X4 FILLER_15_149 ();
 FILLCELL_X1 FILLER_15_153 ();
 FILLCELL_X16 FILLER_15_162 ();
 FILLCELL_X8 FILLER_15_178 ();
 FILLCELL_X1 FILLER_15_186 ();
 FILLCELL_X2 FILLER_15_192 ();
 FILLCELL_X16 FILLER_15_225 ();
 FILLCELL_X4 FILLER_15_241 ();
 FILLCELL_X1 FILLER_15_245 ();
 FILLCELL_X8 FILLER_15_258 ();
 FILLCELL_X4 FILLER_15_266 ();
 FILLCELL_X2 FILLER_15_270 ();
 FILLCELL_X1 FILLER_15_272 ();
 FILLCELL_X4 FILLER_15_287 ();
 FILLCELL_X2 FILLER_15_291 ();
 FILLCELL_X1 FILLER_15_293 ();
 FILLCELL_X2 FILLER_15_322 ();
 FILLCELL_X4 FILLER_15_337 ();
 FILLCELL_X1 FILLER_15_341 ();
 FILLCELL_X4 FILLER_15_344 ();
 FILLCELL_X1 FILLER_15_348 ();
 FILLCELL_X4 FILLER_15_353 ();
 FILLCELL_X2 FILLER_15_357 ();
 FILLCELL_X2 FILLER_15_365 ();
 FILLCELL_X1 FILLER_15_367 ();
 FILLCELL_X8 FILLER_15_372 ();
 FILLCELL_X2 FILLER_15_391 ();
 FILLCELL_X1 FILLER_15_393 ();
 FILLCELL_X1 FILLER_15_401 ();
 FILLCELL_X8 FILLER_15_416 ();
 FILLCELL_X2 FILLER_15_424 ();
 FILLCELL_X1 FILLER_15_426 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_17 ();
 FILLCELL_X1 FILLER_16_57 ();
 FILLCELL_X2 FILLER_16_68 ();
 FILLCELL_X2 FILLER_16_73 ();
 FILLCELL_X2 FILLER_16_82 ();
 FILLCELL_X8 FILLER_16_111 ();
 FILLCELL_X4 FILLER_16_119 ();
 FILLCELL_X1 FILLER_16_123 ();
 FILLCELL_X8 FILLER_16_129 ();
 FILLCELL_X1 FILLER_16_137 ();
 FILLCELL_X16 FILLER_16_159 ();
 FILLCELL_X4 FILLER_16_175 ();
 FILLCELL_X4 FILLER_16_189 ();
 FILLCELL_X1 FILLER_16_193 ();
 FILLCELL_X16 FILLER_16_225 ();
 FILLCELL_X8 FILLER_16_241 ();
 FILLCELL_X1 FILLER_16_249 ();
 FILLCELL_X4 FILLER_16_272 ();
 FILLCELL_X1 FILLER_16_283 ();
 FILLCELL_X1 FILLER_16_309 ();
 FILLCELL_X1 FILLER_16_317 ();
 FILLCELL_X2 FILLER_16_337 ();
 FILLCELL_X1 FILLER_16_343 ();
 FILLCELL_X1 FILLER_16_348 ();
 FILLCELL_X1 FILLER_16_352 ();
 FILLCELL_X1 FILLER_16_362 ();
 FILLCELL_X1 FILLER_16_372 ();
 FILLCELL_X4 FILLER_16_377 ();
 FILLCELL_X2 FILLER_16_381 ();
 FILLCELL_X1 FILLER_16_387 ();
 FILLCELL_X16 FILLER_16_409 ();
 FILLCELL_X2 FILLER_16_425 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_5 ();
 FILLCELL_X1 FILLER_17_8 ();
 FILLCELL_X2 FILLER_17_49 ();
 FILLCELL_X8 FILLER_17_73 ();
 FILLCELL_X1 FILLER_17_81 ();
 FILLCELL_X2 FILLER_17_97 ();
 FILLCELL_X8 FILLER_17_110 ();
 FILLCELL_X4 FILLER_17_118 ();
 FILLCELL_X2 FILLER_17_122 ();
 FILLCELL_X2 FILLER_17_129 ();
 FILLCELL_X1 FILLER_17_131 ();
 FILLCELL_X8 FILLER_17_141 ();
 FILLCELL_X2 FILLER_17_149 ();
 FILLCELL_X1 FILLER_17_154 ();
 FILLCELL_X8 FILLER_17_187 ();
 FILLCELL_X8 FILLER_17_197 ();
 FILLCELL_X4 FILLER_17_205 ();
 FILLCELL_X2 FILLER_17_209 ();
 FILLCELL_X1 FILLER_17_211 ();
 FILLCELL_X2 FILLER_17_222 ();
 FILLCELL_X1 FILLER_17_230 ();
 FILLCELL_X1 FILLER_17_236 ();
 FILLCELL_X1 FILLER_17_262 ();
 FILLCELL_X4 FILLER_17_287 ();
 FILLCELL_X1 FILLER_17_294 ();
 FILLCELL_X1 FILLER_17_298 ();
 FILLCELL_X4 FILLER_17_321 ();
 FILLCELL_X1 FILLER_17_334 ();
 FILLCELL_X2 FILLER_17_351 ();
 FILLCELL_X4 FILLER_17_383 ();
 FILLCELL_X1 FILLER_17_387 ();
 FILLCELL_X1 FILLER_17_400 ();
 FILLCELL_X16 FILLER_17_408 ();
 FILLCELL_X2 FILLER_17_424 ();
 FILLCELL_X1 FILLER_17_426 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_9 ();
 FILLCELL_X2 FILLER_18_12 ();
 FILLCELL_X4 FILLER_18_29 ();
 FILLCELL_X2 FILLER_18_33 ();
 FILLCELL_X1 FILLER_18_35 ();
 FILLCELL_X8 FILLER_18_50 ();
 FILLCELL_X4 FILLER_18_58 ();
 FILLCELL_X8 FILLER_18_72 ();
 FILLCELL_X1 FILLER_18_95 ();
 FILLCELL_X2 FILLER_18_98 ();
 FILLCELL_X4 FILLER_18_113 ();
 FILLCELL_X4 FILLER_18_124 ();
 FILLCELL_X1 FILLER_18_128 ();
 FILLCELL_X4 FILLER_18_166 ();
 FILLCELL_X2 FILLER_18_170 ();
 FILLCELL_X4 FILLER_18_189 ();
 FILLCELL_X1 FILLER_18_203 ();
 FILLCELL_X4 FILLER_18_208 ();
 FILLCELL_X2 FILLER_18_212 ();
 FILLCELL_X2 FILLER_18_218 ();
 FILLCELL_X1 FILLER_18_235 ();
 FILLCELL_X2 FILLER_18_244 ();
 FILLCELL_X1 FILLER_18_246 ();
 FILLCELL_X1 FILLER_18_250 ();
 FILLCELL_X32 FILLER_18_263 ();
 FILLCELL_X2 FILLER_18_295 ();
 FILLCELL_X1 FILLER_18_297 ();
 FILLCELL_X2 FILLER_18_310 ();
 FILLCELL_X4 FILLER_18_314 ();
 FILLCELL_X2 FILLER_18_318 ();
 FILLCELL_X1 FILLER_18_320 ();
 FILLCELL_X2 FILLER_18_344 ();
 FILLCELL_X1 FILLER_18_346 ();
 FILLCELL_X4 FILLER_18_355 ();
 FILLCELL_X2 FILLER_18_359 ();
 FILLCELL_X1 FILLER_18_361 ();
 FILLCELL_X1 FILLER_18_381 ();
 FILLCELL_X1 FILLER_18_389 ();
 FILLCELL_X2 FILLER_18_424 ();
 FILLCELL_X1 FILLER_18_426 ();
 FILLCELL_X1 FILLER_19_4 ();
 FILLCELL_X4 FILLER_19_26 ();
 FILLCELL_X2 FILLER_19_30 ();
 FILLCELL_X16 FILLER_19_50 ();
 FILLCELL_X2 FILLER_19_66 ();
 FILLCELL_X1 FILLER_19_68 ();
 FILLCELL_X2 FILLER_19_130 ();
 FILLCELL_X1 FILLER_19_132 ();
 FILLCELL_X4 FILLER_19_164 ();
 FILLCELL_X1 FILLER_19_168 ();
 FILLCELL_X4 FILLER_19_178 ();
 FILLCELL_X1 FILLER_19_182 ();
 FILLCELL_X8 FILLER_19_193 ();
 FILLCELL_X4 FILLER_19_201 ();
 FILLCELL_X2 FILLER_19_205 ();
 FILLCELL_X2 FILLER_19_217 ();
 FILLCELL_X1 FILLER_19_219 ();
 FILLCELL_X2 FILLER_19_222 ();
 FILLCELL_X1 FILLER_19_255 ();
 FILLCELL_X2 FILLER_19_262 ();
 FILLCELL_X8 FILLER_19_275 ();
 FILLCELL_X4 FILLER_19_283 ();
 FILLCELL_X2 FILLER_19_287 ();
 FILLCELL_X1 FILLER_19_289 ();
 FILLCELL_X2 FILLER_19_344 ();
 FILLCELL_X1 FILLER_19_353 ();
 FILLCELL_X4 FILLER_19_361 ();
 FILLCELL_X2 FILLER_19_365 ();
 FILLCELL_X1 FILLER_19_374 ();
 FILLCELL_X2 FILLER_19_382 ();
 FILLCELL_X2 FILLER_19_387 ();
 FILLCELL_X16 FILLER_19_403 ();
 FILLCELL_X8 FILLER_19_419 ();
 FILLCELL_X2 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_31 ();
 FILLCELL_X16 FILLER_20_46 ();
 FILLCELL_X4 FILLER_20_62 ();
 FILLCELL_X2 FILLER_20_78 ();
 FILLCELL_X1 FILLER_20_93 ();
 FILLCELL_X1 FILLER_20_103 ();
 FILLCELL_X4 FILLER_20_117 ();
 FILLCELL_X16 FILLER_20_136 ();
 FILLCELL_X4 FILLER_20_152 ();
 FILLCELL_X1 FILLER_20_156 ();
 FILLCELL_X2 FILLER_20_193 ();
 FILLCELL_X1 FILLER_20_195 ();
 FILLCELL_X2 FILLER_20_200 ();
 FILLCELL_X1 FILLER_20_202 ();
 FILLCELL_X2 FILLER_20_207 ();
 FILLCELL_X1 FILLER_20_221 ();
 FILLCELL_X1 FILLER_20_230 ();
 FILLCELL_X1 FILLER_20_234 ();
 FILLCELL_X16 FILLER_20_238 ();
 FILLCELL_X2 FILLER_20_254 ();
 FILLCELL_X1 FILLER_20_258 ();
 FILLCELL_X1 FILLER_20_262 ();
 FILLCELL_X32 FILLER_20_268 ();
 FILLCELL_X2 FILLER_20_307 ();
 FILLCELL_X2 FILLER_20_325 ();
 FILLCELL_X8 FILLER_20_334 ();
 FILLCELL_X1 FILLER_20_342 ();
 FILLCELL_X1 FILLER_20_357 ();
 FILLCELL_X8 FILLER_20_369 ();
 FILLCELL_X4 FILLER_20_377 ();
 FILLCELL_X4 FILLER_20_392 ();
 FILLCELL_X2 FILLER_20_396 ();
 FILLCELL_X16 FILLER_20_405 ();
 FILLCELL_X4 FILLER_20_421 ();
 FILLCELL_X2 FILLER_20_425 ();
 FILLCELL_X1 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_6 ();
 FILLCELL_X2 FILLER_21_10 ();
 FILLCELL_X2 FILLER_21_14 ();
 FILLCELL_X1 FILLER_21_16 ();
 FILLCELL_X16 FILLER_21_21 ();
 FILLCELL_X2 FILLER_21_54 ();
 FILLCELL_X1 FILLER_21_56 ();
 FILLCELL_X2 FILLER_21_60 ();
 FILLCELL_X2 FILLER_21_98 ();
 FILLCELL_X1 FILLER_21_100 ();
 FILLCELL_X4 FILLER_21_104 ();
 FILLCELL_X1 FILLER_21_108 ();
 FILLCELL_X4 FILLER_21_114 ();
 FILLCELL_X1 FILLER_21_141 ();
 FILLCELL_X16 FILLER_21_146 ();
 FILLCELL_X1 FILLER_21_162 ();
 FILLCELL_X2 FILLER_21_204 ();
 FILLCELL_X1 FILLER_21_214 ();
 FILLCELL_X8 FILLER_21_223 ();
 FILLCELL_X4 FILLER_21_231 ();
 FILLCELL_X1 FILLER_21_265 ();
 FILLCELL_X16 FILLER_21_270 ();
 FILLCELL_X8 FILLER_21_286 ();
 FILLCELL_X2 FILLER_21_294 ();
 FILLCELL_X1 FILLER_21_296 ();
 FILLCELL_X2 FILLER_21_304 ();
 FILLCELL_X1 FILLER_21_306 ();
 FILLCELL_X4 FILLER_21_352 ();
 FILLCELL_X1 FILLER_21_377 ();
 FILLCELL_X4 FILLER_21_385 ();
 FILLCELL_X4 FILLER_21_399 ();
 FILLCELL_X16 FILLER_21_410 ();
 FILLCELL_X1 FILLER_21_426 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_17 ();
 FILLCELL_X2 FILLER_22_21 ();
 FILLCELL_X1 FILLER_22_23 ();
 FILLCELL_X2 FILLER_22_31 ();
 FILLCELL_X1 FILLER_22_33 ();
 FILLCELL_X4 FILLER_22_71 ();
 FILLCELL_X2 FILLER_22_108 ();
 FILLCELL_X2 FILLER_22_130 ();
 FILLCELL_X1 FILLER_22_132 ();
 FILLCELL_X2 FILLER_22_137 ();
 FILLCELL_X1 FILLER_22_139 ();
 FILLCELL_X2 FILLER_22_144 ();
 FILLCELL_X4 FILLER_22_168 ();
 FILLCELL_X2 FILLER_22_172 ();
 FILLCELL_X2 FILLER_22_184 ();
 FILLCELL_X2 FILLER_22_196 ();
 FILLCELL_X1 FILLER_22_198 ();
 FILLCELL_X2 FILLER_22_204 ();
 FILLCELL_X1 FILLER_22_206 ();
 FILLCELL_X2 FILLER_22_211 ();
 FILLCELL_X1 FILLER_22_213 ();
 FILLCELL_X2 FILLER_22_230 ();
 FILLCELL_X1 FILLER_22_232 ();
 FILLCELL_X4 FILLER_22_240 ();
 FILLCELL_X1 FILLER_22_244 ();
 FILLCELL_X2 FILLER_22_247 ();
 FILLCELL_X2 FILLER_22_271 ();
 FILLCELL_X16 FILLER_22_282 ();
 FILLCELL_X8 FILLER_22_298 ();
 FILLCELL_X2 FILLER_22_306 ();
 FILLCELL_X4 FILLER_22_311 ();
 FILLCELL_X2 FILLER_22_315 ();
 FILLCELL_X1 FILLER_22_329 ();
 FILLCELL_X4 FILLER_22_335 ();
 FILLCELL_X2 FILLER_22_339 ();
 FILLCELL_X8 FILLER_22_353 ();
 FILLCELL_X1 FILLER_22_361 ();
 FILLCELL_X4 FILLER_22_373 ();
 FILLCELL_X2 FILLER_22_382 ();
 FILLCELL_X8 FILLER_22_417 ();
 FILLCELL_X2 FILLER_22_425 ();
 FILLCELL_X16 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_17 ();
 FILLCELL_X1 FILLER_23_32 ();
 FILLCELL_X8 FILLER_23_42 ();
 FILLCELL_X4 FILLER_23_50 ();
 FILLCELL_X1 FILLER_23_58 ();
 FILLCELL_X1 FILLER_23_66 ();
 FILLCELL_X1 FILLER_23_69 ();
 FILLCELL_X1 FILLER_23_77 ();
 FILLCELL_X1 FILLER_23_81 ();
 FILLCELL_X2 FILLER_23_88 ();
 FILLCELL_X4 FILLER_23_118 ();
 FILLCELL_X1 FILLER_23_127 ();
 FILLCELL_X4 FILLER_23_132 ();
 FILLCELL_X2 FILLER_23_136 ();
 FILLCELL_X1 FILLER_23_138 ();
 FILLCELL_X2 FILLER_23_142 ();
 FILLCELL_X8 FILLER_23_148 ();
 FILLCELL_X1 FILLER_23_156 ();
 FILLCELL_X32 FILLER_23_184 ();
 FILLCELL_X2 FILLER_23_220 ();
 FILLCELL_X4 FILLER_23_234 ();
 FILLCELL_X1 FILLER_23_238 ();
 FILLCELL_X4 FILLER_23_243 ();
 FILLCELL_X4 FILLER_23_250 ();
 FILLCELL_X2 FILLER_23_254 ();
 FILLCELL_X1 FILLER_23_256 ();
 FILLCELL_X1 FILLER_23_283 ();
 FILLCELL_X1 FILLER_23_288 ();
 FILLCELL_X1 FILLER_23_306 ();
 FILLCELL_X1 FILLER_23_320 ();
 FILLCELL_X1 FILLER_23_328 ();
 FILLCELL_X1 FILLER_23_332 ();
 FILLCELL_X1 FILLER_23_336 ();
 FILLCELL_X4 FILLER_23_342 ();
 FILLCELL_X2 FILLER_23_346 ();
 FILLCELL_X1 FILLER_23_348 ();
 FILLCELL_X2 FILLER_23_379 ();
 FILLCELL_X4 FILLER_23_391 ();
 FILLCELL_X2 FILLER_23_395 ();
 FILLCELL_X1 FILLER_23_397 ();
 FILLCELL_X1 FILLER_23_402 ();
 FILLCELL_X1 FILLER_23_408 ();
 FILLCELL_X8 FILLER_23_413 ();
 FILLCELL_X4 FILLER_23_421 ();
 FILLCELL_X2 FILLER_23_425 ();
 FILLCELL_X1 FILLER_24_9 ();
 FILLCELL_X1 FILLER_24_20 ();
 FILLCELL_X1 FILLER_24_25 ();
 FILLCELL_X1 FILLER_24_29 ();
 FILLCELL_X1 FILLER_24_88 ();
 FILLCELL_X1 FILLER_24_94 ();
 FILLCELL_X4 FILLER_24_112 ();
 FILLCELL_X2 FILLER_24_120 ();
 FILLCELL_X1 FILLER_24_122 ();
 FILLCELL_X2 FILLER_24_128 ();
 FILLCELL_X2 FILLER_24_134 ();
 FILLCELL_X1 FILLER_24_139 ();
 FILLCELL_X4 FILLER_24_144 ();
 FILLCELL_X2 FILLER_24_148 ();
 FILLCELL_X8 FILLER_24_153 ();
 FILLCELL_X2 FILLER_24_161 ();
 FILLCELL_X1 FILLER_24_163 ();
 FILLCELL_X32 FILLER_24_171 ();
 FILLCELL_X4 FILLER_24_203 ();
 FILLCELL_X2 FILLER_24_207 ();
 FILLCELL_X1 FILLER_24_209 ();
 FILLCELL_X2 FILLER_24_214 ();
 FILLCELL_X1 FILLER_24_216 ();
 FILLCELL_X1 FILLER_24_221 ();
 FILLCELL_X4 FILLER_24_226 ();
 FILLCELL_X2 FILLER_24_230 ();
 FILLCELL_X2 FILLER_24_242 ();
 FILLCELL_X8 FILLER_24_253 ();
 FILLCELL_X2 FILLER_24_261 ();
 FILLCELL_X4 FILLER_24_267 ();
 FILLCELL_X16 FILLER_24_281 ();
 FILLCELL_X8 FILLER_24_297 ();
 FILLCELL_X2 FILLER_24_335 ();
 FILLCELL_X1 FILLER_24_337 ();
 FILLCELL_X4 FILLER_24_342 ();
 FILLCELL_X1 FILLER_24_353 ();
 FILLCELL_X8 FILLER_24_369 ();
 FILLCELL_X4 FILLER_24_377 ();
 FILLCELL_X2 FILLER_24_381 ();
 FILLCELL_X1 FILLER_24_383 ();
 FILLCELL_X1 FILLER_24_389 ();
 FILLCELL_X1 FILLER_24_393 ();
 FILLCELL_X2 FILLER_24_425 ();
 FILLCELL_X2 FILLER_25_1 ();
 FILLCELL_X8 FILLER_25_41 ();
 FILLCELL_X1 FILLER_25_49 ();
 FILLCELL_X1 FILLER_25_57 ();
 FILLCELL_X1 FILLER_25_69 ();
 FILLCELL_X4 FILLER_25_75 ();
 FILLCELL_X2 FILLER_25_79 ();
 FILLCELL_X1 FILLER_25_81 ();
 FILLCELL_X1 FILLER_25_93 ();
 FILLCELL_X2 FILLER_25_101 ();
 FILLCELL_X1 FILLER_25_106 ();
 FILLCELL_X2 FILLER_25_146 ();
 FILLCELL_X1 FILLER_25_148 ();
 FILLCELL_X16 FILLER_25_153 ();
 FILLCELL_X8 FILLER_25_169 ();
 FILLCELL_X2 FILLER_25_177 ();
 FILLCELL_X1 FILLER_25_179 ();
 FILLCELL_X2 FILLER_25_217 ();
 FILLCELL_X1 FILLER_25_219 ();
 FILLCELL_X2 FILLER_25_224 ();
 FILLCELL_X1 FILLER_25_228 ();
 FILLCELL_X1 FILLER_25_233 ();
 FILLCELL_X1 FILLER_25_238 ();
 FILLCELL_X4 FILLER_25_243 ();
 FILLCELL_X2 FILLER_25_252 ();
 FILLCELL_X1 FILLER_25_254 ();
 FILLCELL_X8 FILLER_25_277 ();
 FILLCELL_X2 FILLER_25_307 ();
 FILLCELL_X1 FILLER_25_309 ();
 FILLCELL_X2 FILLER_25_342 ();
 FILLCELL_X8 FILLER_25_352 ();
 FILLCELL_X2 FILLER_25_360 ();
 FILLCELL_X1 FILLER_25_362 ();
 FILLCELL_X4 FILLER_25_367 ();
 FILLCELL_X2 FILLER_25_371 ();
 FILLCELL_X2 FILLER_25_376 ();
 FILLCELL_X2 FILLER_25_382 ();
 FILLCELL_X4 FILLER_25_391 ();
 FILLCELL_X8 FILLER_25_417 ();
 FILLCELL_X2 FILLER_25_425 ();
 FILLCELL_X4 FILLER_26_7 ();
 FILLCELL_X1 FILLER_26_11 ();
 FILLCELL_X4 FILLER_26_28 ();
 FILLCELL_X2 FILLER_26_32 ();
 FILLCELL_X2 FILLER_26_41 ();
 FILLCELL_X1 FILLER_26_43 ();
 FILLCELL_X1 FILLER_26_79 ();
 FILLCELL_X2 FILLER_26_147 ();
 FILLCELL_X1 FILLER_26_166 ();
 FILLCELL_X8 FILLER_26_204 ();
 FILLCELL_X4 FILLER_26_212 ();
 FILLCELL_X2 FILLER_26_216 ();
 FILLCELL_X4 FILLER_26_228 ();
 FILLCELL_X1 FILLER_26_232 ();
 FILLCELL_X8 FILLER_26_240 ();
 FILLCELL_X4 FILLER_26_248 ();
 FILLCELL_X8 FILLER_26_274 ();
 FILLCELL_X2 FILLER_26_282 ();
 FILLCELL_X4 FILLER_26_292 ();
 FILLCELL_X1 FILLER_26_296 ();
 FILLCELL_X2 FILLER_26_345 ();
 FILLCELL_X4 FILLER_26_375 ();
 FILLCELL_X2 FILLER_26_379 ();
 FILLCELL_X16 FILLER_26_388 ();
 FILLCELL_X4 FILLER_26_404 ();
 FILLCELL_X2 FILLER_26_408 ();
 FILLCELL_X8 FILLER_26_414 ();
 FILLCELL_X4 FILLER_26_422 ();
 FILLCELL_X1 FILLER_26_426 ();
 FILLCELL_X2 FILLER_27_1 ();
 FILLCELL_X1 FILLER_27_3 ();
 FILLCELL_X4 FILLER_27_12 ();
 FILLCELL_X2 FILLER_27_16 ();
 FILLCELL_X8 FILLER_27_22 ();
 FILLCELL_X4 FILLER_27_39 ();
 FILLCELL_X2 FILLER_27_43 ();
 FILLCELL_X1 FILLER_27_45 ();
 FILLCELL_X2 FILLER_27_84 ();
 FILLCELL_X8 FILLER_27_100 ();
 FILLCELL_X4 FILLER_27_108 ();
 FILLCELL_X2 FILLER_27_112 ();
 FILLCELL_X2 FILLER_27_143 ();
 FILLCELL_X1 FILLER_27_149 ();
 FILLCELL_X2 FILLER_27_177 ();
 FILLCELL_X1 FILLER_27_183 ();
 FILLCELL_X1 FILLER_27_201 ();
 FILLCELL_X4 FILLER_27_212 ();
 FILLCELL_X1 FILLER_27_218 ();
 FILLCELL_X2 FILLER_27_237 ();
 FILLCELL_X2 FILLER_27_245 ();
 FILLCELL_X1 FILLER_27_247 ();
 FILLCELL_X1 FILLER_27_266 ();
 FILLCELL_X1 FILLER_27_275 ();
 FILLCELL_X16 FILLER_27_286 ();
 FILLCELL_X8 FILLER_27_302 ();
 FILLCELL_X4 FILLER_27_310 ();
 FILLCELL_X8 FILLER_27_318 ();
 FILLCELL_X2 FILLER_27_326 ();
 FILLCELL_X1 FILLER_27_348 ();
 FILLCELL_X2 FILLER_27_377 ();
 FILLCELL_X8 FILLER_27_383 ();
 FILLCELL_X2 FILLER_27_391 ();
 FILLCELL_X8 FILLER_27_402 ();
 FILLCELL_X4 FILLER_28_5 ();
 FILLCELL_X1 FILLER_28_11 ();
 FILLCELL_X8 FILLER_28_23 ();
 FILLCELL_X8 FILLER_28_47 ();
 FILLCELL_X1 FILLER_28_55 ();
 FILLCELL_X4 FILLER_28_72 ();
 FILLCELL_X2 FILLER_28_76 ();
 FILLCELL_X2 FILLER_28_85 ();
 FILLCELL_X4 FILLER_28_91 ();
 FILLCELL_X4 FILLER_28_121 ();
 FILLCELL_X2 FILLER_28_136 ();
 FILLCELL_X8 FILLER_28_143 ();
 FILLCELL_X2 FILLER_28_151 ();
 FILLCELL_X8 FILLER_28_156 ();
 FILLCELL_X1 FILLER_28_164 ();
 FILLCELL_X4 FILLER_28_175 ();
 FILLCELL_X2 FILLER_28_179 ();
 FILLCELL_X1 FILLER_28_181 ();
 FILLCELL_X1 FILLER_28_199 ();
 FILLCELL_X1 FILLER_28_224 ();
 FILLCELL_X8 FILLER_28_244 ();
 FILLCELL_X2 FILLER_28_252 ();
 FILLCELL_X2 FILLER_28_258 ();
 FILLCELL_X1 FILLER_28_260 ();
 FILLCELL_X4 FILLER_28_263 ();
 FILLCELL_X2 FILLER_28_279 ();
 FILLCELL_X2 FILLER_28_287 ();
 FILLCELL_X1 FILLER_28_289 ();
 FILLCELL_X8 FILLER_28_295 ();
 FILLCELL_X2 FILLER_28_303 ();
 FILLCELL_X4 FILLER_28_322 ();
 FILLCELL_X1 FILLER_28_326 ();
 FILLCELL_X4 FILLER_28_348 ();
 FILLCELL_X2 FILLER_28_376 ();
 FILLCELL_X1 FILLER_28_378 ();
 FILLCELL_X8 FILLER_28_388 ();
 FILLCELL_X2 FILLER_28_396 ();
 FILLCELL_X1 FILLER_28_398 ();
 FILLCELL_X8 FILLER_28_416 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X2 FILLER_29_9 ();
 FILLCELL_X1 FILLER_29_11 ();
 FILLCELL_X1 FILLER_29_25 ();
 FILLCELL_X2 FILLER_29_35 ();
 FILLCELL_X1 FILLER_29_37 ();
 FILLCELL_X2 FILLER_29_41 ();
 FILLCELL_X4 FILLER_29_50 ();
 FILLCELL_X1 FILLER_29_54 ();
 FILLCELL_X1 FILLER_29_79 ();
 FILLCELL_X4 FILLER_29_90 ();
 FILLCELL_X1 FILLER_29_94 ();
 FILLCELL_X2 FILLER_29_98 ();
 FILLCELL_X4 FILLER_29_116 ();
 FILLCELL_X1 FILLER_29_123 ();
 FILLCELL_X2 FILLER_29_127 ();
 FILLCELL_X4 FILLER_29_135 ();
 FILLCELL_X2 FILLER_29_139 ();
 FILLCELL_X32 FILLER_29_145 ();
 FILLCELL_X32 FILLER_29_177 ();
 FILLCELL_X2 FILLER_29_209 ();
 FILLCELL_X1 FILLER_29_211 ();
 FILLCELL_X2 FILLER_29_217 ();
 FILLCELL_X8 FILLER_29_223 ();
 FILLCELL_X2 FILLER_29_241 ();
 FILLCELL_X4 FILLER_29_245 ();
 FILLCELL_X2 FILLER_29_249 ();
 FILLCELL_X8 FILLER_29_279 ();
 FILLCELL_X4 FILLER_29_287 ();
 FILLCELL_X2 FILLER_29_291 ();
 FILLCELL_X1 FILLER_29_293 ();
 FILLCELL_X1 FILLER_29_297 ();
 FILLCELL_X1 FILLER_29_315 ();
 FILLCELL_X1 FILLER_29_335 ();
 FILLCELL_X4 FILLER_29_362 ();
 FILLCELL_X1 FILLER_29_366 ();
 FILLCELL_X2 FILLER_29_371 ();
 FILLCELL_X1 FILLER_29_373 ();
 FILLCELL_X1 FILLER_29_383 ();
 FILLCELL_X4 FILLER_29_401 ();
 FILLCELL_X2 FILLER_29_405 ();
 FILLCELL_X2 FILLER_30_5 ();
 FILLCELL_X4 FILLER_30_13 ();
 FILLCELL_X4 FILLER_30_37 ();
 FILLCELL_X1 FILLER_30_41 ();
 FILLCELL_X4 FILLER_30_52 ();
 FILLCELL_X4 FILLER_30_84 ();
 FILLCELL_X4 FILLER_30_101 ();
 FILLCELL_X1 FILLER_30_105 ();
 FILLCELL_X1 FILLER_30_126 ();
 FILLCELL_X16 FILLER_30_135 ();
 FILLCELL_X1 FILLER_30_151 ();
 FILLCELL_X8 FILLER_30_189 ();
 FILLCELL_X4 FILLER_30_197 ();
 FILLCELL_X2 FILLER_30_201 ();
 FILLCELL_X1 FILLER_30_203 ();
 FILLCELL_X16 FILLER_30_206 ();
 FILLCELL_X4 FILLER_30_226 ();
 FILLCELL_X2 FILLER_30_230 ();
 FILLCELL_X1 FILLER_30_232 ();
 FILLCELL_X8 FILLER_30_239 ();
 FILLCELL_X2 FILLER_30_247 ();
 FILLCELL_X1 FILLER_30_268 ();
 FILLCELL_X8 FILLER_30_286 ();
 FILLCELL_X4 FILLER_30_294 ();
 FILLCELL_X2 FILLER_30_298 ();
 FILLCELL_X16 FILLER_30_308 ();
 FILLCELL_X4 FILLER_30_324 ();
 FILLCELL_X2 FILLER_30_328 ();
 FILLCELL_X2 FILLER_30_337 ();
 FILLCELL_X4 FILLER_30_352 ();
 FILLCELL_X2 FILLER_30_356 ();
 FILLCELL_X1 FILLER_30_358 ();
 FILLCELL_X1 FILLER_30_383 ();
 FILLCELL_X16 FILLER_30_390 ();
 FILLCELL_X4 FILLER_30_406 ();
 FILLCELL_X8 FILLER_30_414 ();
 FILLCELL_X4 FILLER_30_422 ();
 FILLCELL_X1 FILLER_30_426 ();
 FILLCELL_X4 FILLER_31_1 ();
 FILLCELL_X2 FILLER_31_5 ();
 FILLCELL_X2 FILLER_31_20 ();
 FILLCELL_X2 FILLER_31_38 ();
 FILLCELL_X8 FILLER_31_47 ();
 FILLCELL_X4 FILLER_31_86 ();
 FILLCELL_X1 FILLER_31_90 ();
 FILLCELL_X16 FILLER_31_105 ();
 FILLCELL_X1 FILLER_31_121 ();
 FILLCELL_X1 FILLER_31_137 ();
 FILLCELL_X4 FILLER_31_151 ();
 FILLCELL_X1 FILLER_31_172 ();
 FILLCELL_X2 FILLER_31_183 ();
 FILLCELL_X1 FILLER_31_190 ();
 FILLCELL_X4 FILLER_31_218 ();
 FILLCELL_X1 FILLER_31_228 ();
 FILLCELL_X8 FILLER_31_240 ();
 FILLCELL_X1 FILLER_31_248 ();
 FILLCELL_X1 FILLER_31_258 ();
 FILLCELL_X1 FILLER_31_263 ();
 FILLCELL_X1 FILLER_31_268 ();
 FILLCELL_X2 FILLER_31_274 ();
 FILLCELL_X1 FILLER_31_276 ();
 FILLCELL_X4 FILLER_31_281 ();
 FILLCELL_X1 FILLER_31_285 ();
 FILLCELL_X1 FILLER_31_292 ();
 FILLCELL_X8 FILLER_31_296 ();
 FILLCELL_X8 FILLER_31_307 ();
 FILLCELL_X4 FILLER_31_315 ();
 FILLCELL_X2 FILLER_31_319 ();
 FILLCELL_X2 FILLER_31_365 ();
 FILLCELL_X1 FILLER_31_367 ();
 FILLCELL_X4 FILLER_31_371 ();
 FILLCELL_X2 FILLER_31_375 ();
 FILLCELL_X1 FILLER_31_394 ();
 FILLCELL_X8 FILLER_31_400 ();
 FILLCELL_X2 FILLER_31_408 ();
 FILLCELL_X1 FILLER_32_1 ();
 FILLCELL_X4 FILLER_32_5 ();
 FILLCELL_X2 FILLER_32_9 ();
 FILLCELL_X1 FILLER_32_11 ();
 FILLCELL_X4 FILLER_32_32 ();
 FILLCELL_X2 FILLER_32_36 ();
 FILLCELL_X1 FILLER_32_38 ();
 FILLCELL_X4 FILLER_32_46 ();
 FILLCELL_X1 FILLER_32_50 ();
 FILLCELL_X8 FILLER_32_77 ();
 FILLCELL_X4 FILLER_32_85 ();
 FILLCELL_X1 FILLER_32_89 ();
 FILLCELL_X1 FILLER_32_101 ();
 FILLCELL_X8 FILLER_32_112 ();
 FILLCELL_X2 FILLER_32_136 ();
 FILLCELL_X1 FILLER_32_138 ();
 FILLCELL_X32 FILLER_32_147 ();
 FILLCELL_X4 FILLER_32_179 ();
 FILLCELL_X2 FILLER_32_183 ();
 FILLCELL_X2 FILLER_32_222 ();
 FILLCELL_X1 FILLER_32_224 ();
 FILLCELL_X4 FILLER_32_229 ();
 FILLCELL_X2 FILLER_32_233 ();
 FILLCELL_X4 FILLER_32_239 ();
 FILLCELL_X1 FILLER_32_243 ();
 FILLCELL_X1 FILLER_32_251 ();
 FILLCELL_X1 FILLER_32_256 ();
 FILLCELL_X4 FILLER_32_268 ();
 FILLCELL_X1 FILLER_32_282 ();
 FILLCELL_X4 FILLER_32_337 ();
 FILLCELL_X16 FILLER_32_367 ();
 FILLCELL_X4 FILLER_32_383 ();
 FILLCELL_X4 FILLER_32_404 ();
 FILLCELL_X8 FILLER_32_412 ();
 FILLCELL_X4 FILLER_32_420 ();
 FILLCELL_X16 FILLER_33_5 ();
 FILLCELL_X2 FILLER_33_21 ();
 FILLCELL_X4 FILLER_33_32 ();
 FILLCELL_X16 FILLER_33_43 ();
 FILLCELL_X4 FILLER_33_59 ();
 FILLCELL_X1 FILLER_33_85 ();
 FILLCELL_X4 FILLER_33_105 ();
 FILLCELL_X2 FILLER_33_116 ();
 FILLCELL_X4 FILLER_33_121 ();
 FILLCELL_X1 FILLER_33_129 ();
 FILLCELL_X2 FILLER_33_133 ();
 FILLCELL_X1 FILLER_33_135 ();
 FILLCELL_X32 FILLER_33_139 ();
 FILLCELL_X32 FILLER_33_171 ();
 FILLCELL_X8 FILLER_33_203 ();
 FILLCELL_X4 FILLER_33_211 ();
 FILLCELL_X2 FILLER_33_215 ();
 FILLCELL_X1 FILLER_33_217 ();
 FILLCELL_X1 FILLER_33_257 ();
 FILLCELL_X1 FILLER_33_269 ();
 FILLCELL_X2 FILLER_33_277 ();
 FILLCELL_X4 FILLER_33_285 ();
 FILLCELL_X2 FILLER_33_292 ();
 FILLCELL_X1 FILLER_33_294 ();
 FILLCELL_X2 FILLER_33_301 ();
 FILLCELL_X1 FILLER_33_303 ();
 FILLCELL_X2 FILLER_33_308 ();
 FILLCELL_X1 FILLER_33_328 ();
 FILLCELL_X2 FILLER_33_338 ();
 FILLCELL_X2 FILLER_33_345 ();
 FILLCELL_X2 FILLER_33_358 ();
 FILLCELL_X1 FILLER_33_360 ();
 FILLCELL_X4 FILLER_33_385 ();
 FILLCELL_X4 FILLER_33_406 ();
 FILLCELL_X2 FILLER_34_1 ();
 FILLCELL_X4 FILLER_34_28 ();
 FILLCELL_X1 FILLER_34_32 ();
 FILLCELL_X1 FILLER_34_40 ();
 FILLCELL_X4 FILLER_34_48 ();
 FILLCELL_X2 FILLER_34_52 ();
 FILLCELL_X1 FILLER_34_66 ();
 FILLCELL_X1 FILLER_34_75 ();
 FILLCELL_X1 FILLER_34_80 ();
 FILLCELL_X2 FILLER_34_88 ();
 FILLCELL_X1 FILLER_34_90 ();
 FILLCELL_X4 FILLER_34_94 ();
 FILLCELL_X1 FILLER_34_98 ();
 FILLCELL_X4 FILLER_34_103 ();
 FILLCELL_X2 FILLER_34_107 ();
 FILLCELL_X1 FILLER_34_114 ();
 FILLCELL_X1 FILLER_34_126 ();
 FILLCELL_X8 FILLER_34_150 ();
 FILLCELL_X4 FILLER_34_158 ();
 FILLCELL_X2 FILLER_34_162 ();
 FILLCELL_X1 FILLER_34_164 ();
 FILLCELL_X4 FILLER_34_192 ();
 FILLCELL_X1 FILLER_34_206 ();
 FILLCELL_X2 FILLER_34_217 ();
 FILLCELL_X1 FILLER_34_219 ();
 FILLCELL_X4 FILLER_34_233 ();
 FILLCELL_X8 FILLER_34_239 ();
 FILLCELL_X16 FILLER_34_254 ();
 FILLCELL_X2 FILLER_34_270 ();
 FILLCELL_X1 FILLER_34_277 ();
 FILLCELL_X8 FILLER_34_282 ();
 FILLCELL_X8 FILLER_34_307 ();
 FILLCELL_X4 FILLER_34_315 ();
 FILLCELL_X1 FILLER_34_319 ();
 FILLCELL_X2 FILLER_34_324 ();
 FILLCELL_X1 FILLER_34_326 ();
 FILLCELL_X8 FILLER_34_390 ();
 FILLCELL_X4 FILLER_34_398 ();
 FILLCELL_X2 FILLER_34_402 ();
 FILLCELL_X16 FILLER_34_408 ();
 FILLCELL_X4 FILLER_35_1 ();
 FILLCELL_X1 FILLER_35_5 ();
 FILLCELL_X2 FILLER_35_8 ();
 FILLCELL_X1 FILLER_35_10 ();
 FILLCELL_X4 FILLER_35_20 ();
 FILLCELL_X1 FILLER_35_24 ();
 FILLCELL_X4 FILLER_35_32 ();
 FILLCELL_X2 FILLER_35_50 ();
 FILLCELL_X2 FILLER_35_72 ();
 FILLCELL_X1 FILLER_35_74 ();
 FILLCELL_X4 FILLER_35_79 ();
 FILLCELL_X4 FILLER_35_86 ();
 FILLCELL_X1 FILLER_35_90 ();
 FILLCELL_X4 FILLER_35_104 ();
 FILLCELL_X1 FILLER_35_113 ();
 FILLCELL_X1 FILLER_35_118 ();
 FILLCELL_X2 FILLER_35_123 ();
 FILLCELL_X2 FILLER_35_146 ();
 FILLCELL_X1 FILLER_35_148 ();
 FILLCELL_X8 FILLER_35_156 ();
 FILLCELL_X2 FILLER_35_164 ();
 FILLCELL_X1 FILLER_35_166 ();
 FILLCELL_X32 FILLER_35_184 ();
 FILLCELL_X8 FILLER_35_216 ();
 FILLCELL_X2 FILLER_35_224 ();
 FILLCELL_X1 FILLER_35_226 ();
 FILLCELL_X2 FILLER_35_241 ();
 FILLCELL_X1 FILLER_35_243 ();
 FILLCELL_X2 FILLER_35_262 ();
 FILLCELL_X1 FILLER_35_264 ();
 FILLCELL_X32 FILLER_35_274 ();
 FILLCELL_X2 FILLER_35_306 ();
 FILLCELL_X2 FILLER_35_331 ();
 FILLCELL_X2 FILLER_35_361 ();
 FILLCELL_X1 FILLER_35_363 ();
 FILLCELL_X2 FILLER_35_368 ();
 FILLCELL_X1 FILLER_35_370 ();
 FILLCELL_X16 FILLER_35_385 ();
 FILLCELL_X2 FILLER_35_401 ();
 FILLCELL_X2 FILLER_35_407 ();
 FILLCELL_X1 FILLER_35_426 ();
 FILLCELL_X4 FILLER_36_1 ();
 FILLCELL_X1 FILLER_36_19 ();
 FILLCELL_X1 FILLER_36_59 ();
 FILLCELL_X1 FILLER_36_65 ();
 FILLCELL_X16 FILLER_36_72 ();
 FILLCELL_X1 FILLER_36_88 ();
 FILLCELL_X2 FILLER_36_107 ();
 FILLCELL_X4 FILLER_36_132 ();
 FILLCELL_X2 FILLER_36_136 ();
 FILLCELL_X1 FILLER_36_138 ();
 FILLCELL_X2 FILLER_36_143 ();
 FILLCELL_X1 FILLER_36_145 ();
 FILLCELL_X8 FILLER_36_150 ();
 FILLCELL_X4 FILLER_36_158 ();
 FILLCELL_X2 FILLER_36_162 ();
 FILLCELL_X4 FILLER_36_181 ();
 FILLCELL_X2 FILLER_36_185 ();
 FILLCELL_X2 FILLER_36_197 ();
 FILLCELL_X2 FILLER_36_216 ();
 FILLCELL_X2 FILLER_36_228 ();
 FILLCELL_X8 FILLER_36_238 ();
 FILLCELL_X1 FILLER_36_250 ();
 FILLCELL_X1 FILLER_36_255 ();
 FILLCELL_X4 FILLER_36_259 ();
 FILLCELL_X1 FILLER_36_271 ();
 FILLCELL_X4 FILLER_36_281 ();
 FILLCELL_X2 FILLER_36_285 ();
 FILLCELL_X1 FILLER_36_287 ();
 FILLCELL_X2 FILLER_36_294 ();
 FILLCELL_X1 FILLER_36_296 ();
 FILLCELL_X8 FILLER_36_303 ();
 FILLCELL_X1 FILLER_36_311 ();
 FILLCELL_X4 FILLER_36_348 ();
 FILLCELL_X4 FILLER_36_369 ();
 FILLCELL_X1 FILLER_36_384 ();
 FILLCELL_X2 FILLER_36_422 ();
 FILLCELL_X2 FILLER_37_11 ();
 FILLCELL_X2 FILLER_37_22 ();
 FILLCELL_X2 FILLER_37_31 ();
 FILLCELL_X1 FILLER_37_33 ();
 FILLCELL_X1 FILLER_37_41 ();
 FILLCELL_X2 FILLER_37_49 ();
 FILLCELL_X1 FILLER_37_51 ();
 FILLCELL_X2 FILLER_37_57 ();
 FILLCELL_X1 FILLER_37_59 ();
 FILLCELL_X2 FILLER_37_78 ();
 FILLCELL_X2 FILLER_37_96 ();
 FILLCELL_X8 FILLER_37_107 ();
 FILLCELL_X2 FILLER_37_115 ();
 FILLCELL_X2 FILLER_37_129 ();
 FILLCELL_X1 FILLER_37_131 ();
 FILLCELL_X2 FILLER_37_144 ();
 FILLCELL_X16 FILLER_37_150 ();
 FILLCELL_X2 FILLER_37_166 ();
 FILLCELL_X4 FILLER_37_195 ();
 FILLCELL_X2 FILLER_37_199 ();
 FILLCELL_X4 FILLER_37_238 ();
 FILLCELL_X2 FILLER_37_242 ();
 FILLCELL_X1 FILLER_37_254 ();
 FILLCELL_X2 FILLER_37_273 ();
 FILLCELL_X1 FILLER_37_275 ();
 FILLCELL_X8 FILLER_37_291 ();
 FILLCELL_X1 FILLER_37_302 ();
 FILLCELL_X16 FILLER_37_306 ();
 FILLCELL_X8 FILLER_37_322 ();
 FILLCELL_X1 FILLER_37_330 ();
 FILLCELL_X2 FILLER_37_348 ();
 FILLCELL_X1 FILLER_37_350 ();
 FILLCELL_X2 FILLER_37_355 ();
 FILLCELL_X1 FILLER_37_357 ();
 FILLCELL_X8 FILLER_37_361 ();
 FILLCELL_X1 FILLER_37_369 ();
 FILLCELL_X16 FILLER_37_387 ();
 FILLCELL_X1 FILLER_37_403 ();
 FILLCELL_X8 FILLER_37_408 ();
 FILLCELL_X4 FILLER_37_416 ();
 FILLCELL_X1 FILLER_37_420 ();
 FILLCELL_X2 FILLER_37_424 ();
 FILLCELL_X1 FILLER_37_426 ();
 FILLCELL_X8 FILLER_38_1 ();
 FILLCELL_X4 FILLER_38_9 ();
 FILLCELL_X2 FILLER_38_33 ();
 FILLCELL_X8 FILLER_38_42 ();
 FILLCELL_X1 FILLER_38_50 ();
 FILLCELL_X1 FILLER_38_62 ();
 FILLCELL_X2 FILLER_38_66 ();
 FILLCELL_X2 FILLER_38_72 ();
 FILLCELL_X2 FILLER_38_79 ();
 FILLCELL_X1 FILLER_38_81 ();
 FILLCELL_X4 FILLER_38_117 ();
 FILLCELL_X1 FILLER_38_121 ();
 FILLCELL_X2 FILLER_38_130 ();
 FILLCELL_X1 FILLER_38_132 ();
 FILLCELL_X16 FILLER_38_154 ();
 FILLCELL_X8 FILLER_38_170 ();
 FILLCELL_X4 FILLER_38_178 ();
 FILLCELL_X1 FILLER_38_182 ();
 FILLCELL_X1 FILLER_38_193 ();
 FILLCELL_X16 FILLER_38_209 ();
 FILLCELL_X4 FILLER_38_225 ();
 FILLCELL_X2 FILLER_38_229 ();
 FILLCELL_X1 FILLER_38_231 ();
 FILLCELL_X1 FILLER_38_254 ();
 FILLCELL_X4 FILLER_38_262 ();
 FILLCELL_X1 FILLER_38_266 ();
 FILLCELL_X1 FILLER_38_280 ();
 FILLCELL_X1 FILLER_38_284 ();
 FILLCELL_X1 FILLER_38_289 ();
 FILLCELL_X2 FILLER_38_299 ();
 FILLCELL_X8 FILLER_38_304 ();
 FILLCELL_X4 FILLER_38_312 ();
 FILLCELL_X2 FILLER_38_339 ();
 FILLCELL_X1 FILLER_38_341 ();
 FILLCELL_X4 FILLER_38_361 ();
 FILLCELL_X1 FILLER_38_365 ();
 FILLCELL_X2 FILLER_38_383 ();
 FILLCELL_X1 FILLER_38_385 ();
 FILLCELL_X4 FILLER_38_393 ();
 FILLCELL_X2 FILLER_38_397 ();
 FILLCELL_X2 FILLER_38_420 ();
 FILLCELL_X1 FILLER_38_422 ();
 FILLCELL_X1 FILLER_38_426 ();
 FILLCELL_X16 FILLER_39_1 ();
 FILLCELL_X2 FILLER_39_17 ();
 FILLCELL_X2 FILLER_39_26 ();
 FILLCELL_X2 FILLER_39_41 ();
 FILLCELL_X1 FILLER_39_43 ();
 FILLCELL_X1 FILLER_39_78 ();
 FILLCELL_X1 FILLER_39_109 ();
 FILLCELL_X1 FILLER_39_114 ();
 FILLCELL_X4 FILLER_39_119 ();
 FILLCELL_X1 FILLER_39_123 ();
 FILLCELL_X4 FILLER_39_128 ();
 FILLCELL_X2 FILLER_39_132 ();
 FILLCELL_X8 FILLER_39_151 ();
 FILLCELL_X32 FILLER_39_162 ();
 FILLCELL_X32 FILLER_39_194 ();
 FILLCELL_X16 FILLER_39_226 ();
 FILLCELL_X1 FILLER_39_242 ();
 FILLCELL_X1 FILLER_39_251 ();
 FILLCELL_X1 FILLER_39_265 ();
 FILLCELL_X1 FILLER_39_280 ();
 FILLCELL_X4 FILLER_39_285 ();
 FILLCELL_X1 FILLER_39_289 ();
 FILLCELL_X2 FILLER_39_293 ();
 FILLCELL_X1 FILLER_39_295 ();
 FILLCELL_X8 FILLER_39_302 ();
 FILLCELL_X2 FILLER_39_310 ();
 FILLCELL_X2 FILLER_39_348 ();
 FILLCELL_X1 FILLER_39_350 ();
 FILLCELL_X4 FILLER_39_354 ();
 FILLCELL_X1 FILLER_39_358 ();
 FILLCELL_X4 FILLER_39_366 ();
 FILLCELL_X2 FILLER_39_370 ();
 FILLCELL_X1 FILLER_39_396 ();
 FILLCELL_X8 FILLER_39_414 ();
 FILLCELL_X4 FILLER_39_422 ();
 FILLCELL_X1 FILLER_39_426 ();
 FILLCELL_X4 FILLER_40_1 ();
 FILLCELL_X1 FILLER_40_5 ();
 FILLCELL_X8 FILLER_40_10 ();
 FILLCELL_X2 FILLER_40_18 ();
 FILLCELL_X4 FILLER_40_29 ();
 FILLCELL_X1 FILLER_40_33 ();
 FILLCELL_X1 FILLER_40_41 ();
 FILLCELL_X2 FILLER_40_49 ();
 FILLCELL_X1 FILLER_40_51 ();
 FILLCELL_X1 FILLER_40_64 ();
 FILLCELL_X2 FILLER_40_76 ();
 FILLCELL_X4 FILLER_40_85 ();
 FILLCELL_X2 FILLER_40_89 ();
 FILLCELL_X1 FILLER_40_91 ();
 FILLCELL_X4 FILLER_40_102 ();
 FILLCELL_X1 FILLER_40_137 ();
 FILLCELL_X1 FILLER_40_148 ();
 FILLCELL_X32 FILLER_40_152 ();
 FILLCELL_X2 FILLER_40_184 ();
 FILLCELL_X1 FILLER_40_186 ();
 FILLCELL_X4 FILLER_40_262 ();
 FILLCELL_X2 FILLER_40_266 ();
 FILLCELL_X1 FILLER_40_268 ();
 FILLCELL_X2 FILLER_40_272 ();
 FILLCELL_X4 FILLER_40_286 ();
 FILLCELL_X1 FILLER_40_290 ();
 FILLCELL_X1 FILLER_40_297 ();
 FILLCELL_X1 FILLER_40_304 ();
 FILLCELL_X16 FILLER_40_322 ();
 FILLCELL_X8 FILLER_40_338 ();
 FILLCELL_X8 FILLER_40_351 ();
 FILLCELL_X4 FILLER_40_359 ();
 FILLCELL_X1 FILLER_40_363 ();
 FILLCELL_X16 FILLER_40_386 ();
 FILLCELL_X2 FILLER_40_419 ();
 FILLCELL_X2 FILLER_40_424 ();
 FILLCELL_X1 FILLER_40_426 ();
 FILLCELL_X2 FILLER_41_1 ();
 FILLCELL_X8 FILLER_41_6 ();
 FILLCELL_X4 FILLER_41_14 ();
 FILLCELL_X2 FILLER_41_18 ();
 FILLCELL_X1 FILLER_41_20 ();
 FILLCELL_X1 FILLER_41_28 ();
 FILLCELL_X1 FILLER_41_36 ();
 FILLCELL_X1 FILLER_41_44 ();
 FILLCELL_X4 FILLER_41_54 ();
 FILLCELL_X1 FILLER_41_58 ();
 FILLCELL_X1 FILLER_41_69 ();
 FILLCELL_X8 FILLER_41_87 ();
 FILLCELL_X8 FILLER_41_100 ();
 FILLCELL_X1 FILLER_41_108 ();
 FILLCELL_X2 FILLER_41_141 ();
 FILLCELL_X2 FILLER_41_146 ();
 FILLCELL_X8 FILLER_41_150 ();
 FILLCELL_X4 FILLER_41_158 ();
 FILLCELL_X1 FILLER_41_162 ();
 FILLCELL_X1 FILLER_41_190 ();
 FILLCELL_X2 FILLER_41_201 ();
 FILLCELL_X2 FILLER_41_213 ();
 FILLCELL_X1 FILLER_41_215 ();
 FILLCELL_X4 FILLER_41_226 ();
 FILLCELL_X2 FILLER_41_230 ();
 FILLCELL_X1 FILLER_41_232 ();
 FILLCELL_X4 FILLER_41_240 ();
 FILLCELL_X1 FILLER_41_244 ();
 FILLCELL_X16 FILLER_41_255 ();
 FILLCELL_X1 FILLER_41_271 ();
 FILLCELL_X1 FILLER_41_297 ();
 FILLCELL_X1 FILLER_41_302 ();
 FILLCELL_X16 FILLER_41_306 ();
 FILLCELL_X8 FILLER_41_322 ();
 FILLCELL_X2 FILLER_41_330 ();
 FILLCELL_X1 FILLER_41_332 ();
 FILLCELL_X32 FILLER_41_364 ();
 FILLCELL_X16 FILLER_41_400 ();
 FILLCELL_X8 FILLER_41_419 ();
 FILLCELL_X2 FILLER_42_1 ();
 FILLCELL_X1 FILLER_42_3 ();
 FILLCELL_X4 FILLER_42_34 ();
 FILLCELL_X1 FILLER_42_38 ();
 FILLCELL_X1 FILLER_42_64 ();
 FILLCELL_X2 FILLER_42_69 ();
 FILLCELL_X2 FILLER_42_85 ();
 FILLCELL_X2 FILLER_42_96 ();
 FILLCELL_X1 FILLER_42_98 ();
 FILLCELL_X1 FILLER_42_103 ();
 FILLCELL_X4 FILLER_42_124 ();
 FILLCELL_X4 FILLER_42_131 ();
 FILLCELL_X1 FILLER_42_148 ();
 FILLCELL_X8 FILLER_42_155 ();
 FILLCELL_X4 FILLER_42_163 ();
 FILLCELL_X2 FILLER_42_167 ();
 FILLCELL_X1 FILLER_42_169 ();
 FILLCELL_X4 FILLER_42_187 ();
 FILLCELL_X1 FILLER_42_191 ();
 FILLCELL_X2 FILLER_42_209 ();
 FILLCELL_X1 FILLER_42_211 ();
 FILLCELL_X4 FILLER_42_235 ();
 FILLCELL_X2 FILLER_42_239 ();
 FILLCELL_X1 FILLER_42_241 ();
 FILLCELL_X16 FILLER_42_254 ();
 FILLCELL_X4 FILLER_42_270 ();
 FILLCELL_X1 FILLER_42_274 ();
 FILLCELL_X16 FILLER_42_301 ();
 FILLCELL_X8 FILLER_42_317 ();
 FILLCELL_X2 FILLER_42_325 ();
 FILLCELL_X4 FILLER_42_331 ();
 FILLCELL_X1 FILLER_42_335 ();
 FILLCELL_X8 FILLER_42_338 ();
 FILLCELL_X1 FILLER_42_370 ();
 FILLCELL_X1 FILLER_42_388 ();
 FILLCELL_X8 FILLER_42_396 ();
 FILLCELL_X2 FILLER_42_404 ();
 FILLCELL_X1 FILLER_42_426 ();
 FILLCELL_X8 FILLER_43_7 ();
 FILLCELL_X1 FILLER_43_15 ();
 FILLCELL_X4 FILLER_43_23 ();
 FILLCELL_X1 FILLER_43_27 ();
 FILLCELL_X8 FILLER_43_30 ();
 FILLCELL_X4 FILLER_43_42 ();
 FILLCELL_X2 FILLER_43_46 ();
 FILLCELL_X1 FILLER_43_48 ();
 FILLCELL_X2 FILLER_43_83 ();
 FILLCELL_X1 FILLER_43_85 ();
 FILLCELL_X2 FILLER_43_104 ();
 FILLCELL_X1 FILLER_43_109 ();
 FILLCELL_X8 FILLER_43_120 ();
 FILLCELL_X1 FILLER_43_128 ();
 FILLCELL_X16 FILLER_43_157 ();
 FILLCELL_X2 FILLER_43_173 ();
 FILLCELL_X4 FILLER_43_185 ();
 FILLCELL_X1 FILLER_43_189 ();
 FILLCELL_X2 FILLER_43_212 ();
 FILLCELL_X1 FILLER_43_214 ();
 FILLCELL_X4 FILLER_43_237 ();
 FILLCELL_X1 FILLER_43_241 ();
 FILLCELL_X2 FILLER_43_250 ();
 FILLCELL_X4 FILLER_43_265 ();
 FILLCELL_X2 FILLER_43_269 ();
 FILLCELL_X1 FILLER_43_276 ();
 FILLCELL_X2 FILLER_43_281 ();
 FILLCELL_X1 FILLER_43_283 ();
 FILLCELL_X2 FILLER_43_289 ();
 FILLCELL_X1 FILLER_43_301 ();
 FILLCELL_X8 FILLER_43_308 ();
 FILLCELL_X2 FILLER_43_320 ();
 FILLCELL_X1 FILLER_43_322 ();
 FILLCELL_X4 FILLER_43_351 ();
 FILLCELL_X2 FILLER_43_355 ();
 FILLCELL_X1 FILLER_43_357 ();
 FILLCELL_X1 FILLER_43_362 ();
 FILLCELL_X8 FILLER_43_365 ();
 FILLCELL_X8 FILLER_43_397 ();
 FILLCELL_X4 FILLER_43_405 ();
 FILLCELL_X1 FILLER_43_409 ();
 FILLCELL_X4 FILLER_44_1 ();
 FILLCELL_X2 FILLER_44_8 ();
 FILLCELL_X1 FILLER_44_18 ();
 FILLCELL_X1 FILLER_44_26 ();
 FILLCELL_X1 FILLER_44_31 ();
 FILLCELL_X1 FILLER_44_41 ();
 FILLCELL_X2 FILLER_44_46 ();
 FILLCELL_X1 FILLER_44_48 ();
 FILLCELL_X4 FILLER_44_56 ();
 FILLCELL_X2 FILLER_44_60 ();
 FILLCELL_X1 FILLER_44_62 ();
 FILLCELL_X2 FILLER_44_74 ();
 FILLCELL_X2 FILLER_44_81 ();
 FILLCELL_X1 FILLER_44_83 ();
 FILLCELL_X4 FILLER_44_87 ();
 FILLCELL_X2 FILLER_44_91 ();
 FILLCELL_X1 FILLER_44_93 ();
 FILLCELL_X2 FILLER_44_133 ();
 FILLCELL_X8 FILLER_44_146 ();
 FILLCELL_X2 FILLER_44_158 ();
 FILLCELL_X4 FILLER_44_187 ();
 FILLCELL_X2 FILLER_44_191 ();
 FILLCELL_X8 FILLER_44_218 ();
 FILLCELL_X1 FILLER_44_226 ();
 FILLCELL_X4 FILLER_44_235 ();
 FILLCELL_X2 FILLER_44_239 ();
 FILLCELL_X2 FILLER_44_257 ();
 FILLCELL_X1 FILLER_44_263 ();
 FILLCELL_X4 FILLER_44_271 ();
 FILLCELL_X1 FILLER_44_275 ();
 FILLCELL_X1 FILLER_44_297 ();
 FILLCELL_X2 FILLER_44_301 ();
 FILLCELL_X4 FILLER_44_320 ();
 FILLCELL_X2 FILLER_44_324 ();
 FILLCELL_X4 FILLER_44_330 ();
 FILLCELL_X1 FILLER_44_334 ();
 FILLCELL_X1 FILLER_44_337 ();
 FILLCELL_X2 FILLER_44_372 ();
 FILLCELL_X8 FILLER_44_391 ();
 FILLCELL_X4 FILLER_44_399 ();
 FILLCELL_X1 FILLER_44_403 ();
 FILLCELL_X8 FILLER_44_408 ();
 FILLCELL_X4 FILLER_44_416 ();
 FILLCELL_X1 FILLER_44_420 ();
 FILLCELL_X2 FILLER_45_4 ();
 FILLCELL_X1 FILLER_45_13 ();
 FILLCELL_X4 FILLER_45_28 ();
 FILLCELL_X2 FILLER_45_32 ();
 FILLCELL_X1 FILLER_45_34 ();
 FILLCELL_X2 FILLER_45_80 ();
 FILLCELL_X1 FILLER_45_82 ();
 FILLCELL_X2 FILLER_45_90 ();
 FILLCELL_X8 FILLER_45_101 ();
 FILLCELL_X1 FILLER_45_128 ();
 FILLCELL_X16 FILLER_45_136 ();
 FILLCELL_X2 FILLER_45_152 ();
 FILLCELL_X1 FILLER_45_154 ();
 FILLCELL_X1 FILLER_45_182 ();
 FILLCELL_X2 FILLER_45_210 ();
 FILLCELL_X2 FILLER_45_222 ();
 FILLCELL_X2 FILLER_45_236 ();
 FILLCELL_X1 FILLER_45_242 ();
 FILLCELL_X1 FILLER_45_262 ();
 FILLCELL_X1 FILLER_45_266 ();
 FILLCELL_X1 FILLER_45_272 ();
 FILLCELL_X8 FILLER_45_304 ();
 FILLCELL_X4 FILLER_45_312 ();
 FILLCELL_X16 FILLER_45_337 ();
 FILLCELL_X8 FILLER_45_361 ();
 FILLCELL_X4 FILLER_45_371 ();
 FILLCELL_X16 FILLER_45_382 ();
 FILLCELL_X8 FILLER_45_398 ();
 FILLCELL_X1 FILLER_45_406 ();
 FILLCELL_X2 FILLER_46_1 ();
 FILLCELL_X1 FILLER_46_6 ();
 FILLCELL_X4 FILLER_46_28 ();
 FILLCELL_X2 FILLER_46_46 ();
 FILLCELL_X4 FILLER_46_60 ();
 FILLCELL_X2 FILLER_46_64 ();
 FILLCELL_X1 FILLER_46_66 ();
 FILLCELL_X4 FILLER_46_74 ();
 FILLCELL_X1 FILLER_46_78 ();
 FILLCELL_X16 FILLER_46_84 ();
 FILLCELL_X8 FILLER_46_100 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X8 FILLER_46_161 ();
 FILLCELL_X4 FILLER_46_169 ();
 FILLCELL_X2 FILLER_46_173 ();
 FILLCELL_X1 FILLER_46_175 ();
 FILLCELL_X8 FILLER_46_203 ();
 FILLCELL_X2 FILLER_46_211 ();
 FILLCELL_X1 FILLER_46_217 ();
 FILLCELL_X2 FILLER_46_226 ();
 FILLCELL_X1 FILLER_46_235 ();
 FILLCELL_X1 FILLER_46_240 ();
 FILLCELL_X1 FILLER_46_249 ();
 FILLCELL_X8 FILLER_46_260 ();
 FILLCELL_X8 FILLER_46_302 ();
 FILLCELL_X4 FILLER_46_329 ();
 FILLCELL_X2 FILLER_46_333 ();
 FILLCELL_X1 FILLER_46_335 ();
 FILLCELL_X2 FILLER_46_344 ();
 FILLCELL_X4 FILLER_46_348 ();
 FILLCELL_X2 FILLER_46_352 ();
 FILLCELL_X2 FILLER_46_375 ();
 FILLCELL_X4 FILLER_46_398 ();
 FILLCELL_X1 FILLER_46_423 ();
 FILLCELL_X4 FILLER_47_5 ();
 FILLCELL_X1 FILLER_47_9 ();
 FILLCELL_X2 FILLER_47_17 ();
 FILLCELL_X1 FILLER_47_42 ();
 FILLCELL_X2 FILLER_47_50 ();
 FILLCELL_X2 FILLER_47_66 ();
 FILLCELL_X2 FILLER_47_89 ();
 FILLCELL_X1 FILLER_47_91 ();
 FILLCELL_X8 FILLER_47_126 ();
 FILLCELL_X4 FILLER_47_134 ();
 FILLCELL_X8 FILLER_47_155 ();
 FILLCELL_X4 FILLER_47_163 ();
 FILLCELL_X2 FILLER_47_167 ();
 FILLCELL_X1 FILLER_47_169 ();
 FILLCELL_X32 FILLER_47_180 ();
 FILLCELL_X16 FILLER_47_212 ();
 FILLCELL_X8 FILLER_47_228 ();
 FILLCELL_X2 FILLER_47_236 ();
 FILLCELL_X1 FILLER_47_238 ();
 FILLCELL_X2 FILLER_47_263 ();
 FILLCELL_X2 FILLER_47_282 ();
 FILLCELL_X2 FILLER_47_294 ();
 FILLCELL_X1 FILLER_47_296 ();
 FILLCELL_X16 FILLER_47_303 ();
 FILLCELL_X4 FILLER_47_319 ();
 FILLCELL_X1 FILLER_47_323 ();
 FILLCELL_X4 FILLER_47_328 ();
 FILLCELL_X1 FILLER_47_332 ();
 FILLCELL_X16 FILLER_47_354 ();
 FILLCELL_X8 FILLER_47_370 ();
 FILLCELL_X2 FILLER_47_378 ();
 FILLCELL_X8 FILLER_47_397 ();
 FILLCELL_X2 FILLER_47_405 ();
 FILLCELL_X1 FILLER_48_4 ();
 FILLCELL_X1 FILLER_48_9 ();
 FILLCELL_X16 FILLER_48_14 ();
 FILLCELL_X1 FILLER_48_30 ();
 FILLCELL_X1 FILLER_48_38 ();
 FILLCELL_X1 FILLER_48_46 ();
 FILLCELL_X1 FILLER_48_54 ();
 FILLCELL_X2 FILLER_48_60 ();
 FILLCELL_X1 FILLER_48_70 ();
 FILLCELL_X1 FILLER_48_76 ();
 FILLCELL_X2 FILLER_48_89 ();
 FILLCELL_X2 FILLER_48_95 ();
 FILLCELL_X1 FILLER_48_97 ();
 FILLCELL_X1 FILLER_48_107 ();
 FILLCELL_X2 FILLER_48_115 ();
 FILLCELL_X1 FILLER_48_117 ();
 FILLCELL_X8 FILLER_48_132 ();
 FILLCELL_X1 FILLER_48_140 ();
 FILLCELL_X2 FILLER_48_158 ();
 FILLCELL_X4 FILLER_48_170 ();
 FILLCELL_X16 FILLER_48_177 ();
 FILLCELL_X4 FILLER_48_193 ();
 FILLCELL_X2 FILLER_48_197 ();
 FILLCELL_X1 FILLER_48_199 ();
 FILLCELL_X2 FILLER_48_227 ();
 FILLCELL_X8 FILLER_48_243 ();
 FILLCELL_X16 FILLER_48_262 ();
 FILLCELL_X2 FILLER_48_278 ();
 FILLCELL_X1 FILLER_48_280 ();
 FILLCELL_X1 FILLER_48_294 ();
 FILLCELL_X16 FILLER_48_302 ();
 FILLCELL_X4 FILLER_48_318 ();
 FILLCELL_X1 FILLER_48_322 ();
 FILLCELL_X16 FILLER_48_340 ();
 FILLCELL_X8 FILLER_48_356 ();
 FILLCELL_X2 FILLER_48_364 ();
 FILLCELL_X1 FILLER_48_366 ();
 FILLCELL_X16 FILLER_48_384 ();
 FILLCELL_X1 FILLER_48_400 ();
 FILLCELL_X2 FILLER_48_424 ();
 FILLCELL_X1 FILLER_48_426 ();
 FILLCELL_X1 FILLER_49_1 ();
 FILLCELL_X8 FILLER_49_30 ();
 FILLCELL_X2 FILLER_49_38 ();
 FILLCELL_X2 FILLER_49_67 ();
 FILLCELL_X1 FILLER_49_69 ();
 FILLCELL_X16 FILLER_49_75 ();
 FILLCELL_X4 FILLER_49_91 ();
 FILLCELL_X1 FILLER_49_99 ();
 FILLCELL_X2 FILLER_49_104 ();
 FILLCELL_X2 FILLER_49_113 ();
 FILLCELL_X2 FILLER_49_122 ();
 FILLCELL_X16 FILLER_49_131 ();
 FILLCELL_X8 FILLER_49_147 ();
 FILLCELL_X2 FILLER_49_165 ();
 FILLCELL_X8 FILLER_49_184 ();
 FILLCELL_X2 FILLER_49_192 ();
 FILLCELL_X4 FILLER_49_211 ();
 FILLCELL_X1 FILLER_49_215 ();
 FILLCELL_X1 FILLER_49_230 ();
 FILLCELL_X1 FILLER_49_235 ();
 FILLCELL_X1 FILLER_49_240 ();
 FILLCELL_X2 FILLER_49_248 ();
 FILLCELL_X1 FILLER_49_254 ();
 FILLCELL_X4 FILLER_49_260 ();
 FILLCELL_X1 FILLER_49_264 ();
 FILLCELL_X1 FILLER_49_275 ();
 FILLCELL_X32 FILLER_49_306 ();
 FILLCELL_X32 FILLER_49_338 ();
 FILLCELL_X16 FILLER_49_370 ();
 FILLCELL_X2 FILLER_49_386 ();
 FILLCELL_X1 FILLER_49_388 ();
 FILLCELL_X32 FILLER_49_392 ();
 FILLCELL_X2 FILLER_49_424 ();
 FILLCELL_X1 FILLER_49_426 ();
 FILLCELL_X1 FILLER_50_13 ();
 FILLCELL_X4 FILLER_50_31 ();
 FILLCELL_X2 FILLER_50_35 ();
 FILLCELL_X1 FILLER_50_37 ();
 FILLCELL_X2 FILLER_50_52 ();
 FILLCELL_X1 FILLER_50_54 ();
 FILLCELL_X8 FILLER_50_60 ();
 FILLCELL_X4 FILLER_50_68 ();
 FILLCELL_X1 FILLER_50_72 ();
 FILLCELL_X8 FILLER_50_83 ();
 FILLCELL_X2 FILLER_50_91 ();
 FILLCELL_X8 FILLER_50_114 ();
 FILLCELL_X4 FILLER_50_122 ();
 FILLCELL_X2 FILLER_50_126 ();
 FILLCELL_X32 FILLER_50_130 ();
 FILLCELL_X1 FILLER_50_179 ();
 FILLCELL_X1 FILLER_50_210 ();
 FILLCELL_X8 FILLER_50_226 ();
 FILLCELL_X1 FILLER_50_234 ();
 FILLCELL_X2 FILLER_50_241 ();
 FILLCELL_X1 FILLER_50_243 ();
 FILLCELL_X1 FILLER_50_246 ();
 FILLCELL_X4 FILLER_50_251 ();
 FILLCELL_X1 FILLER_50_255 ();
 FILLCELL_X1 FILLER_50_260 ();
 FILLCELL_X8 FILLER_50_269 ();
 FILLCELL_X2 FILLER_50_277 ();
 FILLCELL_X32 FILLER_50_300 ();
 FILLCELL_X8 FILLER_50_332 ();
 FILLCELL_X4 FILLER_50_340 ();
 FILLCELL_X32 FILLER_50_361 ();
 FILLCELL_X32 FILLER_50_393 ();
 FILLCELL_X2 FILLER_50_425 ();
 FILLCELL_X4 FILLER_51_1 ();
 FILLCELL_X2 FILLER_51_17 ();
 FILLCELL_X1 FILLER_51_28 ();
 FILLCELL_X16 FILLER_51_47 ();
 FILLCELL_X16 FILLER_51_83 ();
 FILLCELL_X2 FILLER_51_99 ();
 FILLCELL_X1 FILLER_51_101 ();
 FILLCELL_X4 FILLER_51_109 ();
 FILLCELL_X1 FILLER_51_113 ();
 FILLCELL_X8 FILLER_51_127 ();
 FILLCELL_X4 FILLER_51_135 ();
 FILLCELL_X1 FILLER_51_139 ();
 FILLCELL_X2 FILLER_51_162 ();
 FILLCELL_X32 FILLER_51_174 ();
 FILLCELL_X16 FILLER_51_206 ();
 FILLCELL_X4 FILLER_51_222 ();
 FILLCELL_X2 FILLER_51_237 ();
 FILLCELL_X2 FILLER_51_246 ();
 FILLCELL_X2 FILLER_51_250 ();
 FILLCELL_X2 FILLER_51_264 ();
 FILLCELL_X1 FILLER_51_266 ();
 FILLCELL_X2 FILLER_51_277 ();
 FILLCELL_X32 FILLER_51_285 ();
 FILLCELL_X32 FILLER_51_317 ();
 FILLCELL_X32 FILLER_51_349 ();
 FILLCELL_X32 FILLER_51_381 ();
 FILLCELL_X8 FILLER_51_413 ();
 FILLCELL_X4 FILLER_51_421 ();
 FILLCELL_X2 FILLER_51_425 ();
 FILLCELL_X2 FILLER_52_1 ();
 FILLCELL_X1 FILLER_52_3 ();
 FILLCELL_X16 FILLER_52_25 ();
 FILLCELL_X4 FILLER_52_41 ();
 FILLCELL_X4 FILLER_52_54 ();
 FILLCELL_X4 FILLER_52_60 ();
 FILLCELL_X2 FILLER_52_66 ();
 FILLCELL_X1 FILLER_52_75 ();
 FILLCELL_X16 FILLER_52_80 ();
 FILLCELL_X4 FILLER_52_96 ();
 FILLCELL_X8 FILLER_52_104 ();
 FILLCELL_X2 FILLER_52_112 ();
 FILLCELL_X1 FILLER_52_114 ();
 FILLCELL_X1 FILLER_52_132 ();
 FILLCELL_X2 FILLER_52_152 ();
 FILLCELL_X1 FILLER_52_174 ();
 FILLCELL_X2 FILLER_52_178 ();
 FILLCELL_X1 FILLER_52_180 ();
 FILLCELL_X1 FILLER_52_183 ();
 FILLCELL_X2 FILLER_52_194 ();
 FILLCELL_X1 FILLER_52_202 ();
 FILLCELL_X1 FILLER_52_207 ();
 FILLCELL_X8 FILLER_52_224 ();
 FILLCELL_X4 FILLER_52_232 ();
 FILLCELL_X1 FILLER_52_236 ();
 FILLCELL_X2 FILLER_52_256 ();
 FILLCELL_X1 FILLER_52_258 ();
 FILLCELL_X4 FILLER_52_262 ();
 FILLCELL_X2 FILLER_52_266 ();
 FILLCELL_X4 FILLER_52_277 ();
 FILLCELL_X2 FILLER_52_281 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X8 FILLER_52_417 ();
 FILLCELL_X2 FILLER_52_425 ();
 FILLCELL_X8 FILLER_53_1 ();
 FILLCELL_X4 FILLER_53_9 ();
 FILLCELL_X2 FILLER_53_13 ();
 FILLCELL_X1 FILLER_53_15 ();
 FILLCELL_X8 FILLER_53_51 ();
 FILLCELL_X4 FILLER_53_59 ();
 FILLCELL_X2 FILLER_53_63 ();
 FILLCELL_X1 FILLER_53_65 ();
 FILLCELL_X2 FILLER_53_86 ();
 FILLCELL_X1 FILLER_53_88 ();
 FILLCELL_X1 FILLER_53_93 ();
 FILLCELL_X4 FILLER_53_100 ();
 FILLCELL_X2 FILLER_53_104 ();
 FILLCELL_X2 FILLER_53_127 ();
 FILLCELL_X32 FILLER_53_132 ();
 FILLCELL_X4 FILLER_53_164 ();
 FILLCELL_X2 FILLER_53_182 ();
 FILLCELL_X2 FILLER_53_195 ();
 FILLCELL_X4 FILLER_53_206 ();
 FILLCELL_X2 FILLER_53_221 ();
 FILLCELL_X2 FILLER_53_229 ();
 FILLCELL_X1 FILLER_53_231 ();
 FILLCELL_X2 FILLER_53_239 ();
 FILLCELL_X1 FILLER_53_241 ();
 FILLCELL_X2 FILLER_53_246 ();
 FILLCELL_X1 FILLER_53_256 ();
 FILLCELL_X1 FILLER_53_261 ();
 FILLCELL_X2 FILLER_53_266 ();
 FILLCELL_X2 FILLER_53_272 ();
 FILLCELL_X2 FILLER_53_280 ();
 FILLCELL_X32 FILLER_53_300 ();
 FILLCELL_X32 FILLER_53_332 ();
 FILLCELL_X32 FILLER_53_364 ();
 FILLCELL_X16 FILLER_53_396 ();
 FILLCELL_X8 FILLER_53_412 ();
 FILLCELL_X4 FILLER_53_420 ();
 FILLCELL_X2 FILLER_53_424 ();
 FILLCELL_X1 FILLER_53_426 ();
 FILLCELL_X16 FILLER_54_1 ();
 FILLCELL_X8 FILLER_54_17 ();
 FILLCELL_X4 FILLER_54_25 ();
 FILLCELL_X1 FILLER_54_29 ();
 FILLCELL_X1 FILLER_54_50 ();
 FILLCELL_X1 FILLER_54_61 ();
 FILLCELL_X2 FILLER_54_65 ();
 FILLCELL_X1 FILLER_54_73 ();
 FILLCELL_X1 FILLER_54_78 ();
 FILLCELL_X1 FILLER_54_89 ();
 FILLCELL_X2 FILLER_54_134 ();
 FILLCELL_X8 FILLER_54_173 ();
 FILLCELL_X4 FILLER_54_181 ();
 FILLCELL_X4 FILLER_54_218 ();
 FILLCELL_X1 FILLER_54_222 ();
 FILLCELL_X4 FILLER_54_233 ();
 FILLCELL_X1 FILLER_54_237 ();
 FILLCELL_X1 FILLER_54_245 ();
 FILLCELL_X1 FILLER_54_253 ();
 FILLCELL_X1 FILLER_54_262 ();
 FILLCELL_X1 FILLER_54_266 ();
 FILLCELL_X1 FILLER_54_270 ();
 FILLCELL_X1 FILLER_54_282 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X8 FILLER_54_417 ();
 FILLCELL_X2 FILLER_54_425 ();
 FILLCELL_X16 FILLER_55_1 ();
 FILLCELL_X8 FILLER_55_17 ();
 FILLCELL_X4 FILLER_55_25 ();
 FILLCELL_X2 FILLER_55_29 ();
 FILLCELL_X1 FILLER_55_31 ();
 FILLCELL_X2 FILLER_55_58 ();
 FILLCELL_X2 FILLER_55_77 ();
 FILLCELL_X16 FILLER_55_83 ();
 FILLCELL_X8 FILLER_55_99 ();
 FILLCELL_X1 FILLER_55_107 ();
 FILLCELL_X4 FILLER_55_125 ();
 FILLCELL_X8 FILLER_55_139 ();
 FILLCELL_X1 FILLER_55_147 ();
 FILLCELL_X1 FILLER_55_251 ();
 FILLCELL_X1 FILLER_55_254 ();
 FILLCELL_X1 FILLER_55_276 ();
 FILLCELL_X32 FILLER_55_281 ();
 FILLCELL_X32 FILLER_55_313 ();
 FILLCELL_X32 FILLER_55_345 ();
 FILLCELL_X32 FILLER_55_377 ();
 FILLCELL_X16 FILLER_55_409 ();
 FILLCELL_X2 FILLER_55_425 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X8 FILLER_56_33 ();
 FILLCELL_X16 FILLER_56_52 ();
 FILLCELL_X4 FILLER_56_68 ();
 FILLCELL_X1 FILLER_56_76 ();
 FILLCELL_X8 FILLER_56_80 ();
 FILLCELL_X1 FILLER_56_91 ();
 FILLCELL_X4 FILLER_56_98 ();
 FILLCELL_X8 FILLER_56_105 ();
 FILLCELL_X4 FILLER_56_113 ();
 FILLCELL_X1 FILLER_56_117 ();
 FILLCELL_X8 FILLER_56_122 ();
 FILLCELL_X4 FILLER_56_130 ();
 FILLCELL_X2 FILLER_56_134 ();
 FILLCELL_X2 FILLER_56_139 ();
 FILLCELL_X2 FILLER_56_149 ();
 FILLCELL_X1 FILLER_56_151 ();
 FILLCELL_X2 FILLER_56_156 ();
 FILLCELL_X1 FILLER_56_158 ();
 FILLCELL_X32 FILLER_56_169 ();
 FILLCELL_X32 FILLER_56_201 ();
 FILLCELL_X8 FILLER_56_233 ();
 FILLCELL_X4 FILLER_56_241 ();
 FILLCELL_X2 FILLER_56_245 ();
 FILLCELL_X1 FILLER_56_249 ();
 FILLCELL_X2 FILLER_56_254 ();
 FILLCELL_X1 FILLER_56_256 ();
 FILLCELL_X32 FILLER_56_267 ();
 FILLCELL_X32 FILLER_56_299 ();
 FILLCELL_X8 FILLER_56_331 ();
 FILLCELL_X2 FILLER_56_339 ();
 FILLCELL_X16 FILLER_56_344 ();
 FILLCELL_X1 FILLER_56_360 ();
 FILLCELL_X32 FILLER_56_364 ();
 FILLCELL_X16 FILLER_56_396 ();
 FILLCELL_X8 FILLER_56_412 ();
 FILLCELL_X4 FILLER_56_420 ();
 FILLCELL_X2 FILLER_56_424 ();
 FILLCELL_X1 FILLER_56_426 ();
endmodule
