module lfsr (bit_out,
    clk,
    enable,
    load,
    rst_n,
    lfsr_out,
    seed);
 output bit_out;
 input clk;
 input enable;
 input load;
 input rst_n;
 output [7:0] lfsr_out;
 input [7:0] seed;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net20;

 sky130_fd_sc_hd__clkbuf_2 _34_ (.A(net2),
    .X(_08_));
 sky130_fd_sc_hd__buf_2 _35_ (.A(_08_),
    .X(_09_));
 sky130_fd_sc_hd__buf_6 _36_ (.A(enable),
    .X(_10_));
 sky130_fd_sc_hd__mux2i_1 _37_ (.A0(net11),
    .A1(net13),
    .S(_10_),
    .Y(_11_));
 sky130_fd_sc_hd__nand2_1 _38_ (.A(_09_),
    .B(net3),
    .Y(_12_));
 sky130_fd_sc_hd__o21ai_0 _39_ (.A1(_09_),
    .A2(_11_),
    .B1(_12_),
    .Y(_00_));
 sky130_fd_sc_hd__mux2i_1 _40_ (.A0(net13),
    .A1(net14),
    .S(_10_),
    .Y(_13_));
 sky130_fd_sc_hd__nand2_1 _41_ (.A(_09_),
    .B(net4),
    .Y(_14_));
 sky130_fd_sc_hd__o21ai_0 _42_ (.A1(_09_),
    .A2(_13_),
    .B1(_14_),
    .Y(_01_));
 sky130_fd_sc_hd__mux2i_1 _43_ (.A0(net14),
    .A1(net15),
    .S(_10_),
    .Y(_15_));
 sky130_fd_sc_hd__nand2_1 _44_ (.A(_09_),
    .B(net5),
    .Y(_16_));
 sky130_fd_sc_hd__o21ai_0 _45_ (.A1(_09_),
    .A2(_15_),
    .B1(_16_),
    .Y(_02_));
 sky130_fd_sc_hd__mux2i_1 _46_ (.A0(net15),
    .A1(net16),
    .S(_10_),
    .Y(_17_));
 sky130_fd_sc_hd__nand2_1 _47_ (.A(_09_),
    .B(net6),
    .Y(_18_));
 sky130_fd_sc_hd__o21ai_0 _48_ (.A1(_08_),
    .A2(_17_),
    .B1(_18_),
    .Y(_03_));
 sky130_fd_sc_hd__mux2i_1 _49_ (.A0(net16),
    .A1(net17),
    .S(_10_),
    .Y(_19_));
 sky130_fd_sc_hd__nand2_1 _50_ (.A(_09_),
    .B(net7),
    .Y(_20_));
 sky130_fd_sc_hd__o21ai_0 _51_ (.A1(_08_),
    .A2(_19_),
    .B1(_20_),
    .Y(_04_));
 sky130_fd_sc_hd__mux2i_1 _52_ (.A0(net17),
    .A1(net18),
    .S(_10_),
    .Y(_21_));
 sky130_fd_sc_hd__nand2_1 _53_ (.A(_09_),
    .B(net8),
    .Y(_22_));
 sky130_fd_sc_hd__o21ai_0 _54_ (.A1(_08_),
    .A2(_21_),
    .B1(_22_),
    .Y(_05_));
 sky130_fd_sc_hd__mux2i_1 _55_ (.A0(net18),
    .A1(net19),
    .S(_10_),
    .Y(_23_));
 sky130_fd_sc_hd__nand2_1 _56_ (.A(_09_),
    .B(net9),
    .Y(_24_));
 sky130_fd_sc_hd__o21ai_0 _57_ (.A1(_08_),
    .A2(_23_),
    .B1(_24_),
    .Y(_06_));
 sky130_fd_sc_hd__or4b_1 _58_ (.A(net2),
    .B(net15),
    .C(net19),
    .D_N(_10_),
    .X(_25_));
 sky130_fd_sc_hd__nand3b_1 _59_ (.A_N(_08_),
    .B(net15),
    .C(net19),
    .Y(_26_));
 sky130_fd_sc_hd__xnor2_1 _60_ (.A(net16),
    .B(net17),
    .Y(_27_));
 sky130_fd_sc_hd__a21oi_1 _61_ (.A1(_25_),
    .A2(_26_),
    .B1(_27_),
    .Y(_28_));
 sky130_fd_sc_hd__nor4bb_1 _62_ (.A(_08_),
    .B(net19),
    .C_N(net15),
    .D_N(_10_),
    .Y(_29_));
 sky130_fd_sc_hd__nor3b_1 _63_ (.A(_08_),
    .B(net15),
    .C_N(net19),
    .Y(_30_));
 sky130_fd_sc_hd__o21ai_0 _64_ (.A1(_29_),
    .A2(_30_),
    .B1(_27_),
    .Y(_31_));
 sky130_fd_sc_hd__nor2_1 _65_ (.A(_08_),
    .B(_10_),
    .Y(_32_));
 sky130_fd_sc_hd__a22oi_1 _66_ (.A1(_08_),
    .A2(net10),
    .B1(_32_),
    .B2(net19),
    .Y(_33_));
 sky130_fd_sc_hd__nand3b_1 _67_ (.A_N(_28_),
    .B(_31_),
    .C(_33_),
    .Y(_07_));
 sky130_fd_sc_hd__clkbuf_1 _68_ (.A(net11),
    .X(net12));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[0]$_DFFE_PN0P_  (.D(_00_),
    .Q(net11),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[1]$_DFFE_PN0P_  (.D(_01_),
    .Q(net13),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[2]$_DFFE_PN0P_  (.D(_02_),
    .Q(net14),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \lfsr_reg[3]$_DFFE_PN0P_  (.D(_03_),
    .Q(net15),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[4]$_DFFE_PN0P_  (.D(_04_),
    .Q(net16),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[5]$_DFFE_PN0P_  (.D(_05_),
    .Q(net17),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[6]$_DFFE_PN0P_  (.D(_06_),
    .Q(net18),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \lfsr_reg[7]$_DFFE_PN0P_  (.D(_07_),
    .Q(net19),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__buf_2 hold1 (.A(net20),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_49 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(load),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(seed[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(seed[1]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(seed[2]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(seed[3]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(seed[4]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(seed[5]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(seed[6]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(seed[7]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net11),
    .X(bit_out));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net12),
    .X(lfsr_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(lfsr_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(lfsr_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(lfsr_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(lfsr_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(lfsr_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(lfsr_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(lfsr_out[7]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net20));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_137 ();
endmodule
