module clock_domain_crossing (dst_clk,
    dst_ready,
    dst_rst_n,
    dst_valid,
    src_clk,
    src_ready,
    src_rst_n,
    src_valid,
    dst_data,
    src_data);
 input dst_clk;
 input dst_ready;
 input dst_rst_n;
 output dst_valid;
 input src_clk;
 output src_ready;
 input src_rst_n;
 input src_valid;
 output [31:0] dst_data;
 input [31:0] src_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire dst_ack;
 wire dst_req_prev;
 wire \dst_req_sync[0] ;
 wire \dst_req_sync[1] ;
 wire src_ack;
 wire \src_ack_sync[0] ;
 wire \src_data_reg[0] ;
 wire \src_data_reg[10] ;
 wire \src_data_reg[11] ;
 wire \src_data_reg[12] ;
 wire \src_data_reg[13] ;
 wire \src_data_reg[14] ;
 wire \src_data_reg[15] ;
 wire \src_data_reg[16] ;
 wire \src_data_reg[17] ;
 wire \src_data_reg[18] ;
 wire \src_data_reg[19] ;
 wire \src_data_reg[1] ;
 wire \src_data_reg[20] ;
 wire \src_data_reg[21] ;
 wire \src_data_reg[22] ;
 wire \src_data_reg[23] ;
 wire \src_data_reg[24] ;
 wire \src_data_reg[25] ;
 wire \src_data_reg[26] ;
 wire \src_data_reg[27] ;
 wire \src_data_reg[28] ;
 wire \src_data_reg[29] ;
 wire \src_data_reg[2] ;
 wire \src_data_reg[30] ;
 wire \src_data_reg[31] ;
 wire \src_data_reg[3] ;
 wire \src_data_reg[4] ;
 wire \src_data_reg[5] ;
 wire \src_data_reg[6] ;
 wire \src_data_reg[7] ;
 wire \src_data_reg[8] ;
 wire \src_data_reg[9] ;
 wire src_req;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire clknet_0_src_clk;
 wire clknet_2_0__leaf_src_clk;
 wire clknet_2_1__leaf_src_clk;
 wire clknet_2_2__leaf_src_clk;
 wire clknet_2_3__leaf_src_clk;
 wire net72;

 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _082_ (.A1(src_req),
    .A2(src_ack),
    .ZN(net71));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _083_ (.A1(\dst_req_sync[1] ),
    .A2(net4),
    .B(dst_ack),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _084_ (.I(net4),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _085_ (.A1(\dst_req_sync[1] ),
    .A2(_068_),
    .B(dst_ack),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _086_ (.A1(dst_req_prev),
    .A2(_067_),
    .B(_069_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _087_ (.A1(dst_req_prev),
    .A2(\dst_req_sync[1] ),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _088_ (.I(_070_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _089_ (.I(_071_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _090_ (.I0(net38),
    .I1(\src_data_reg[0] ),
    .S(_072_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _091_ (.I0(net39),
    .I1(\src_data_reg[10] ),
    .S(_072_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _092_ (.I0(net40),
    .I1(\src_data_reg[11] ),
    .S(_072_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _093_ (.I0(net41),
    .I1(\src_data_reg[12] ),
    .S(_072_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _094_ (.I0(net42),
    .I1(\src_data_reg[13] ),
    .S(_072_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _095_ (.I0(net43),
    .I1(\src_data_reg[14] ),
    .S(_072_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _096_ (.I0(net44),
    .I1(\src_data_reg[15] ),
    .S(_072_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _097_ (.I0(net45),
    .I1(\src_data_reg[16] ),
    .S(_072_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _098_ (.I0(net46),
    .I1(\src_data_reg[17] ),
    .S(_072_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _099_ (.I(_071_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _100_ (.I0(net47),
    .I1(\src_data_reg[18] ),
    .S(_073_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _101_ (.I0(net48),
    .I1(\src_data_reg[19] ),
    .S(_073_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _102_ (.I0(net49),
    .I1(\src_data_reg[1] ),
    .S(_073_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _103_ (.I0(net50),
    .I1(\src_data_reg[20] ),
    .S(_073_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _104_ (.I0(net51),
    .I1(\src_data_reg[21] ),
    .S(_073_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _105_ (.I0(net52),
    .I1(\src_data_reg[22] ),
    .S(_073_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _106_ (.I0(net53),
    .I1(\src_data_reg[23] ),
    .S(_073_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _107_ (.I0(net54),
    .I1(\src_data_reg[24] ),
    .S(_073_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _108_ (.I0(net55),
    .I1(\src_data_reg[25] ),
    .S(_073_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _109_ (.I0(net56),
    .I1(\src_data_reg[26] ),
    .S(_073_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _110_ (.I(_071_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _111_ (.I0(net57),
    .I1(\src_data_reg[27] ),
    .S(_074_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _112_ (.I0(net58),
    .I1(\src_data_reg[28] ),
    .S(_074_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _113_ (.I0(net59),
    .I1(\src_data_reg[29] ),
    .S(_074_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _114_ (.I0(net60),
    .I1(\src_data_reg[2] ),
    .S(_074_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _115_ (.I0(net61),
    .I1(\src_data_reg[30] ),
    .S(_074_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _116_ (.I0(net62),
    .I1(\src_data_reg[31] ),
    .S(_074_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _117_ (.I0(net63),
    .I1(\src_data_reg[3] ),
    .S(_074_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _118_ (.I0(net64),
    .I1(\src_data_reg[4] ),
    .S(_074_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _119_ (.I0(net65),
    .I1(\src_data_reg[5] ),
    .S(_074_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _120_ (.I0(net66),
    .I1(\src_data_reg[6] ),
    .S(_074_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _121_ (.I0(net67),
    .I1(\src_data_reg[7] ),
    .S(_071_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _122_ (.I0(net68),
    .I1(\src_data_reg[8] ),
    .S(_071_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _123_ (.I0(net69),
    .I1(\src_data_reg[9] ),
    .S(_071_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _124_ (.I(net3),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _125_ (.A1(_075_),
    .A2(net70),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _126_ (.A1(_072_),
    .A2(_076_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _127_ (.A1(net37),
    .A2(net71),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _128_ (.I(_077_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _129_ (.I0(\src_data_reg[0] ),
    .I1(net5),
    .S(_078_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _130_ (.I0(\src_data_reg[10] ),
    .I1(net6),
    .S(_078_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _131_ (.I0(\src_data_reg[11] ),
    .I1(net7),
    .S(_078_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _132_ (.I0(\src_data_reg[12] ),
    .I1(net8),
    .S(_078_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _133_ (.I0(\src_data_reg[13] ),
    .I1(net9),
    .S(_078_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _134_ (.I0(\src_data_reg[14] ),
    .I1(net10),
    .S(_078_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _135_ (.I0(\src_data_reg[15] ),
    .I1(net11),
    .S(_078_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _136_ (.I0(\src_data_reg[16] ),
    .I1(net12),
    .S(_078_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _137_ (.I0(\src_data_reg[17] ),
    .I1(net13),
    .S(_078_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _138_ (.I0(\src_data_reg[18] ),
    .I1(net14),
    .S(_078_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _139_ (.I(_077_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _140_ (.I0(\src_data_reg[19] ),
    .I1(net15),
    .S(_079_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _141_ (.I0(\src_data_reg[1] ),
    .I1(net16),
    .S(_079_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _142_ (.I0(\src_data_reg[20] ),
    .I1(net17),
    .S(_079_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _143_ (.I0(\src_data_reg[21] ),
    .I1(net18),
    .S(_079_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _144_ (.I0(\src_data_reg[22] ),
    .I1(net19),
    .S(_079_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _145_ (.I0(\src_data_reg[23] ),
    .I1(net20),
    .S(_079_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _146_ (.I0(\src_data_reg[24] ),
    .I1(net21),
    .S(_079_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _147_ (.I0(\src_data_reg[25] ),
    .I1(net22),
    .S(_079_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _148_ (.I0(\src_data_reg[26] ),
    .I1(net23),
    .S(_079_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _149_ (.I0(\src_data_reg[27] ),
    .I1(net24),
    .S(_079_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _150_ (.I(_077_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _151_ (.I0(\src_data_reg[28] ),
    .I1(net25),
    .S(_080_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _152_ (.I0(\src_data_reg[29] ),
    .I1(net26),
    .S(_080_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _153_ (.I0(\src_data_reg[2] ),
    .I1(net27),
    .S(_080_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _154_ (.I0(\src_data_reg[30] ),
    .I1(net28),
    .S(_080_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _155_ (.I0(\src_data_reg[31] ),
    .I1(net29),
    .S(_080_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _156_ (.I0(\src_data_reg[3] ),
    .I1(net30),
    .S(_080_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _157_ (.I0(\src_data_reg[4] ),
    .I1(net31),
    .S(_080_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _158_ (.I0(\src_data_reg[5] ),
    .I1(net32),
    .S(_080_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _159_ (.I0(\src_data_reg[6] ),
    .I1(net33),
    .S(_080_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _160_ (.I0(\src_data_reg[7] ),
    .I1(net34),
    .S(_080_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _161_ (.I0(\src_data_reg[8] ),
    .I1(net35),
    .S(_077_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _162_ (.I0(\src_data_reg[9] ),
    .I1(net36),
    .S(_077_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _163_ (.I(src_ack),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _164_ (.I0(src_req),
    .I1(_081_),
    .S(net37),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dst_ack$_DFFE_PP_  (.D(_000_),
    .CLK(net2),
    .Q(dst_ack));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[0]$_DFFE_PN0P_  (.D(_001_),
    .RN(net4),
    .CLK(net2),
    .Q(net38));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[10]$_DFFE_PN0P_  (.D(_002_),
    .RN(net4),
    .CLK(net2),
    .Q(net39));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[11]$_DFFE_PN0P_  (.D(_003_),
    .RN(net4),
    .CLK(net2),
    .Q(net40));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[12]$_DFFE_PN0P_  (.D(_004_),
    .RN(net4),
    .CLK(net2),
    .Q(net41));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[13]$_DFFE_PN0P_  (.D(_005_),
    .RN(net4),
    .CLK(net2),
    .Q(net42));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[14]$_DFFE_PN0P_  (.D(_006_),
    .RN(net4),
    .CLK(net2),
    .Q(net43));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[15]$_DFFE_PN0P_  (.D(_007_),
    .RN(net4),
    .CLK(net2),
    .Q(net44));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[16]$_DFFE_PN0P_  (.D(_008_),
    .RN(net4),
    .CLK(net2),
    .Q(net45));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[17]$_DFFE_PN0P_  (.D(_009_),
    .RN(net4),
    .CLK(net2),
    .Q(net46));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[18]$_DFFE_PN0P_  (.D(_010_),
    .RN(net4),
    .CLK(net2),
    .Q(net47));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[19]$_DFFE_PN0P_  (.D(_011_),
    .RN(net4),
    .CLK(net2),
    .Q(net48));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[1]$_DFFE_PN0P_  (.D(_012_),
    .RN(net4),
    .CLK(net2),
    .Q(net49));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[20]$_DFFE_PN0P_  (.D(_013_),
    .RN(net4),
    .CLK(net2),
    .Q(net50));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[21]$_DFFE_PN0P_  (.D(_014_),
    .RN(net4),
    .CLK(net2),
    .Q(net51));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[22]$_DFFE_PN0P_  (.D(_015_),
    .RN(net4),
    .CLK(net2),
    .Q(net52));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[23]$_DFFE_PN0P_  (.D(_016_),
    .RN(net4),
    .CLK(net2),
    .Q(net53));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[24]$_DFFE_PN0P_  (.D(_017_),
    .RN(net4),
    .CLK(net2),
    .Q(net54));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[25]$_DFFE_PN0P_  (.D(_018_),
    .RN(net4),
    .CLK(net2),
    .Q(net55));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[26]$_DFFE_PN0P_  (.D(_019_),
    .RN(net4),
    .CLK(net2),
    .Q(net56));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[27]$_DFFE_PN0P_  (.D(_020_),
    .RN(net4),
    .CLK(net2),
    .Q(net57));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[28]$_DFFE_PN0P_  (.D(_021_),
    .RN(net4),
    .CLK(net2),
    .Q(net58));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[29]$_DFFE_PN0P_  (.D(_022_),
    .RN(net4),
    .CLK(net2),
    .Q(net59));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[2]$_DFFE_PN0P_  (.D(_023_),
    .RN(net4),
    .CLK(net2),
    .Q(net60));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[30]$_DFFE_PN0P_  (.D(_024_),
    .RN(net4),
    .CLK(net2),
    .Q(net61));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[31]$_DFFE_PN0P_  (.D(_025_),
    .RN(net4),
    .CLK(net2),
    .Q(net62));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[3]$_DFFE_PN0P_  (.D(_026_),
    .RN(net4),
    .CLK(net2),
    .Q(net63));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[4]$_DFFE_PN0P_  (.D(_027_),
    .RN(net4),
    .CLK(net2),
    .Q(net64));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[5]$_DFFE_PN0P_  (.D(_028_),
    .RN(net4),
    .CLK(net2),
    .Q(net65));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[6]$_DFFE_PN0P_  (.D(_029_),
    .RN(net4),
    .CLK(net2),
    .Q(net66));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[7]$_DFFE_PN0P_  (.D(_030_),
    .RN(net4),
    .CLK(net2),
    .Q(net67));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[8]$_DFFE_PN0P_  (.D(_031_),
    .RN(net4),
    .CLK(net2),
    .Q(net68));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_data[9]$_DFFE_PN0P_  (.D(_032_),
    .RN(net4),
    .CLK(net2),
    .Q(net69));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_req_prev$_DFF_PN0_  (.D(\dst_req_sync[1] ),
    .RN(net4),
    .CLK(net2),
    .Q(dst_req_prev));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_req_sync[0]$_DFF_PN0_  (.D(src_req),
    .RN(net4),
    .CLK(net2),
    .Q(\dst_req_sync[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_req_sync[1]$_DFF_PN0_  (.D(\dst_req_sync[0] ),
    .RN(net4),
    .CLK(net2),
    .Q(\dst_req_sync[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dst_valid$_DFFE_PN0P_  (.D(_033_),
    .RN(net4),
    .CLK(net2),
    .Q(net70));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_ack_sync[0]$_DFF_PN0_  (.D(dst_ack),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\src_ack_sync[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_ack_sync[1]$_DFF_PN0_  (.D(\src_ack_sync[0] ),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(src_ack));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[0]$_DFFE_PN0P_  (.D(_034_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[10]$_DFFE_PN0P_  (.D(_035_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[11]$_DFFE_PN0P_  (.D(_036_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[12]$_DFFE_PN0P_  (.D(_037_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[13]$_DFFE_PN0P_  (.D(_038_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[14]$_DFFE_PN0P_  (.D(_039_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[15]$_DFFE_PN0P_  (.D(_040_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[16]$_DFFE_PN0P_  (.D(_041_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[17]$_DFFE_PN0P_  (.D(_042_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[18]$_DFFE_PN0P_  (.D(_043_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_src_clk),
    .Q(\src_data_reg[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[19]$_DFFE_PN0P_  (.D(_044_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[1]$_DFFE_PN0P_  (.D(_045_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[20]$_DFFE_PN0P_  (.D(_046_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[21]$_DFFE_PN0P_  (.D(_047_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[22]$_DFFE_PN0P_  (.D(_048_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[23]$_DFFE_PN0P_  (.D(_049_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[24]$_DFFE_PN0P_  (.D(_050_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[25]$_DFFE_PN0P_  (.D(_051_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[26]$_DFFE_PN0P_  (.D(_052_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_src_clk),
    .Q(\src_data_reg[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[27]$_DFFE_PN0P_  (.D(_053_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[28]$_DFFE_PN0P_  (.D(_054_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[29]$_DFFE_PN0P_  (.D(_055_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[2]$_DFFE_PN0P_  (.D(_056_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[30]$_DFFE_PN0P_  (.D(_057_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[31]$_DFFE_PN0P_  (.D(_058_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[3]$_DFFE_PN0P_  (.D(_059_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[4]$_DFFE_PN0P_  (.D(_060_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[5]$_DFFE_PN0P_  (.D(_061_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[6]$_DFFE_PN0P_  (.D(_062_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[7]$_DFFE_PN0P_  (.D(_063_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_src_clk),
    .Q(\src_data_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[8]$_DFFE_PN0P_  (.D(_064_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_data_reg[9]$_DFFE_PN0P_  (.D(_065_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(\src_data_reg[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \src_req$_DFFE_PN0P_  (.D(_066_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_src_clk),
    .Q(src_req));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 hold1 (.I(net72),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_67 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_68 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_69 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_70 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_71 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_72 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_73 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_74 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_75 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_76 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_77 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input1 (.I(dst_clk),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(dst_ready),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 input3 (.I(dst_rst_n),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(src_data[0]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(src_data[10]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(src_data[11]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(src_data[12]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(src_data[13]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(src_data[14]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(src_data[15]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(src_data[16]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(src_data[17]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(src_data[18]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(src_data[19]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(src_data[1]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(src_data[20]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(src_data[21]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(src_data[22]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(src_data[23]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(src_data[24]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(src_data[25]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(src_data[26]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(src_data[27]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(src_data[28]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(src_data[29]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(src_data[2]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(src_data[30]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(src_data[31]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(src_data[3]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(src_data[4]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(src_data[5]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(src_data[6]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input33 (.I(src_data[7]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(src_data[8]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(src_data[9]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(src_valid),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output37 (.I(net38),
    .Z(dst_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output38 (.I(net39),
    .Z(dst_data[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net40),
    .Z(dst_data[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output40 (.I(net41),
    .Z(dst_data[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output41 (.I(net42),
    .Z(dst_data[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output42 (.I(net43),
    .Z(dst_data[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output43 (.I(net44),
    .Z(dst_data[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output44 (.I(net45),
    .Z(dst_data[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output45 (.I(net46),
    .Z(dst_data[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output46 (.I(net47),
    .Z(dst_data[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output47 (.I(net48),
    .Z(dst_data[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net49),
    .Z(dst_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net50),
    .Z(dst_data[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net51),
    .Z(dst_data[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output51 (.I(net52),
    .Z(dst_data[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output52 (.I(net53),
    .Z(dst_data[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output53 (.I(net54),
    .Z(dst_data[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output54 (.I(net55),
    .Z(dst_data[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output55 (.I(net56),
    .Z(dst_data[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output56 (.I(net57),
    .Z(dst_data[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output57 (.I(net58),
    .Z(dst_data[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output58 (.I(net59),
    .Z(dst_data[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output59 (.I(net60),
    .Z(dst_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output60 (.I(net61),
    .Z(dst_data[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output61 (.I(net62),
    .Z(dst_data[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net63),
    .Z(dst_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net64),
    .Z(dst_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net65),
    .Z(dst_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net66),
    .Z(dst_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net67),
    .Z(dst_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net68),
    .Z(dst_data[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net69),
    .Z(dst_data[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net70),
    .Z(dst_valid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net71),
    .Z(src_ready));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_src_clk (.I(src_clk),
    .Z(clknet_0_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_0__f_src_clk (.I(clknet_0_src_clk),
    .Z(clknet_2_0__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_1__f_src_clk (.I(clknet_0_src_clk),
    .Z(clknet_2_1__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_2__f_src_clk (.I(clknet_0_src_clk),
    .Z(clknet_2_2__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_3__f_src_clk (.I(clknet_0_src_clk),
    .Z(clknet_2_3__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload0 (.I(clknet_2_2__leaf_src_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(src_rst_n),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_270 ();
endmodule
