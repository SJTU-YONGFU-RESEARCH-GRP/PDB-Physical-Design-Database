module parameterized_uart_tx (clk,
    rst_n,
    tx,
    tx_busy,
    tx_start,
    data_in);
 input clk;
 input rst_n;
 output tx;
 output tx_busy;
 input tx_start;
 input [7:0] data_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire \bit_index[0] ;
 wire \bit_index[1] ;
 wire \bit_index[2] ;
 wire \clk_counter[0] ;
 wire \clk_counter[1] ;
 wire \clk_counter[2] ;
 wire \clk_counter[3] ;
 wire \clk_counter[4] ;
 wire \clk_counter[5] ;
 wire \data_reg[0] ;
 wire \data_reg[1] ;
 wire \data_reg[2] ;
 wire \data_reg[3] ;
 wire \data_reg[4] ;
 wire \data_reg[5] ;
 wire \data_reg[6] ;
 wire \data_reg[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _095_ (.I(\clk_counter[1] ),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _096_ (.I(\bit_index[0] ),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _097_ (.A1(\state[2] ),
    .A2(\state[0] ),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _098_ (.I(\state[2] ),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _099_ (.A1(_056_),
    .A2(\state[0] ),
    .A3(_088_),
    .A4(\bit_index[0] ),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _100_ (.A1(\clk_counter[3] ),
    .A2(\clk_counter[2] ),
    .A3(\clk_counter[1] ),
    .A4(_091_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _101_ (.A1(\clk_counter[5] ),
    .A2(\clk_counter[4] ),
    .A3(_058_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _102_ (.I(_059_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _103_ (.I0(_054_),
    .I1(_057_),
    .S(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _104_ (.I(\state[1] ),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _105_ (.A1(_054_),
    .A2(_055_),
    .B1(_061_),
    .B2(_062_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _106_ (.I(\bit_index[1] ),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _107_ (.A1(_087_),
    .A2(_055_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _108_ (.I0(_063_),
    .I1(_064_),
    .S(_059_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _109_ (.A1(_063_),
    .A2(_055_),
    .B1(_065_),
    .B2(_062_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _110_ (.I(\bit_index[2] ),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _111_ (.A1(_089_),
    .A2(_055_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _112_ (.I0(_066_),
    .I1(_067_),
    .S(_059_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _113_ (.A1(_066_),
    .A2(_055_),
    .B1(_068_),
    .B2(_062_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _114_ (.A1(\state[1] ),
    .A2(\state[0] ),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _115_ (.A1(\clk_counter[0] ),
    .A2(_069_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _116_ (.A1(\clk_counter[0] ),
    .A2(_069_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _117_ (.A1(_060_),
    .A2(_070_),
    .B(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _118_ (.A1(\state[1] ),
    .A2(\state[0] ),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _119_ (.A1(\clk_counter[0] ),
    .A2(_060_),
    .A3(_073_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _120_ (.I(\state[2] ),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _121_ (.I0(_072_),
    .I1(_074_),
    .S(_075_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _122_ (.A1(_092_),
    .A2(_060_),
    .A3(_073_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _123_ (.A1(\clk_counter[1] ),
    .A2(_069_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _124_ (.A1(_092_),
    .A2(_060_),
    .A3(_069_),
    .B(_077_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _125_ (.I0(_076_),
    .I1(_078_),
    .S(_056_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _126_ (.I(\clk_counter[2] ),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _127_ (.A1(\state[1] ),
    .A2(\state[0] ),
    .B(_056_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _128_ (.A1(_056_),
    .A2(_079_),
    .A3(_069_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _129_ (.A1(_075_),
    .A2(_073_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _130_ (.A1(\clk_counter[2] ),
    .A2(_093_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _131_ (.A1(_060_),
    .A2(_081_),
    .A3(_082_),
    .A4(_083_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _132_ (.A1(_079_),
    .A2(_080_),
    .B(_084_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _133_ (.I(\clk_counter[3] ),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _134_ (.A1(_056_),
    .A2(_085_),
    .A3(_069_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _135_ (.A1(\clk_counter[2] ),
    .A2(\clk_counter[1] ),
    .A3(\clk_counter[0] ),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _136_ (.A1(\clk_counter[3] ),
    .A2(_023_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _137_ (.A1(\clk_counter[3] ),
    .A2(\clk_counter[2] ),
    .A3(\clk_counter[1] ),
    .A4(\clk_counter[0] ),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _138_ (.A1(_082_),
    .A2(_022_),
    .A3(_024_),
    .A4(_025_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _139_ (.A1(_085_),
    .A2(_080_),
    .B1(_026_),
    .B2(_060_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _140_ (.A1(\clk_counter[3] ),
    .A2(\clk_counter[2] ),
    .A3(_093_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _141_ (.A1(\clk_counter[4] ),
    .A2(_027_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _142_ (.A1(\clk_counter[4] ),
    .A2(_027_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _143_ (.A1(_080_),
    .A2(_028_),
    .B(_029_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _144_ (.I(\clk_counter[4] ),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _145_ (.A1(_060_),
    .A2(_082_),
    .A3(_030_),
    .B1(_080_),
    .B2(_031_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _146_ (.A1(\clk_counter[5] ),
    .A2(\clk_counter[4] ),
    .A3(_058_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _147_ (.A1(_032_),
    .A2(_069_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _148_ (.A1(\clk_counter[4] ),
    .A2(_080_),
    .A3(_025_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _149_ (.A1(_032_),
    .A2(_069_),
    .B1(_034_),
    .B2(\clk_counter[5] ),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _150_ (.A1(_075_),
    .A2(_033_),
    .B(_035_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _151_ (.A1(_075_),
    .A2(net11),
    .A3(_073_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _152_ (.I0(\data_reg[0] ),
    .I1(net2),
    .S(_036_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _153_ (.I0(\data_reg[1] ),
    .I1(net3),
    .S(_036_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _154_ (.I0(\data_reg[2] ),
    .I1(net4),
    .S(_036_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _155_ (.I0(\data_reg[3] ),
    .I1(net5),
    .S(_036_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _156_ (.I0(\data_reg[4] ),
    .I1(net6),
    .S(_036_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _157_ (.I0(\data_reg[5] ),
    .I1(net7),
    .S(_036_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _158_ (.I0(\data_reg[6] ),
    .I1(net8),
    .S(_036_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _159_ (.I0(\data_reg[7] ),
    .I1(net9),
    .S(_036_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _160_ (.A1(\state[0] ),
    .A2(_032_),
    .B1(_073_),
    .B2(net11),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _161_ (.A1(_056_),
    .A2(_037_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _162_ (.A1(\state[0] ),
    .A2(_088_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _163_ (.A1(\clk_counter[5] ),
    .A2(\clk_counter[4] ),
    .A3(_058_),
    .A4(_038_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _164_ (.A1(_062_),
    .A2(\state[0] ),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _165_ (.A1(\state[1] ),
    .A2(_039_),
    .B1(_040_),
    .B2(_060_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _166_ (.A1(_056_),
    .A2(_041_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _167_ (.A1(_056_),
    .A2(_062_),
    .A3(_039_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _168_ (.A1(_075_),
    .A2(_060_),
    .A3(_069_),
    .B(_042_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _169_ (.I0(\data_reg[2] ),
    .I1(\data_reg[3] ),
    .I2(\data_reg[6] ),
    .I3(\data_reg[7] ),
    .S0(\bit_index[0] ),
    .S1(\bit_index[2] ),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _170_ (.A1(_063_),
    .A2(_043_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _171_ (.I0(\data_reg[4] ),
    .I1(\data_reg[5] ),
    .S(\bit_index[0] ),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _172_ (.A1(\bit_index[1] ),
    .A2(_066_),
    .A3(_045_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _173_ (.I0(\data_reg[0] ),
    .I1(\data_reg[1] ),
    .S(\bit_index[0] ),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _174_ (.A1(\bit_index[1] ),
    .A2(\bit_index[2] ),
    .A3(_047_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _175_ (.A1(_055_),
    .A2(_044_),
    .A3(_046_),
    .A4(_048_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _176_ (.A1(_056_),
    .A2(net12),
    .Z(_050_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _177_ (.A1(_073_),
    .A2(_049_),
    .A3(_050_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _178_ (.I0(net11),
    .I1(net13),
    .S(_069_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _179_ (.A1(_075_),
    .A2(_051_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _180_ (.A1(_056_),
    .A2(net13),
    .A3(_032_),
    .A4(_073_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _181_ (.A1(_052_),
    .A2(_053_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _182_ (.A(\bit_index[0] ),
    .B(\bit_index[1] ),
    .CO(_086_),
    .S(_087_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _183_ (.A(\bit_index[2] ),
    .B(_086_),
    .CO(_088_),
    .S(_089_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _184_ (.A(\clk_counter[0] ),
    .B(_090_),
    .CO(_091_),
    .S(_092_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _185_ (.A(\clk_counter[0] ),
    .B(\clk_counter[1] ),
    .CO(_093_),
    .S(_094_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_index[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\bit_index[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_index[1]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\bit_index[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_index[2]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\bit_index[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[0]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\clk_counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[1]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\clk_counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[2]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\clk_counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[3]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\clk_counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[4]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\clk_counter[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \clk_counter[5]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\clk_counter[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[0]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\data_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[1]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\data_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[2]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\data_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[3]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\data_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[4]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\data_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[5]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\data_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[6]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\data_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \data_reg[7]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\data_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[0]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[1]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[2]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \tx$_DFFE_PN1P_  (.D(_020_),
    .SETN(net10),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net12));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_busy$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 hold1 (.I(net10),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_44 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_55 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(data_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(data_in[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(data_in[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(data_in[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(data_in[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(data_in[5]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(data_in[6]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(data_in[7]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input9 (.I(rst_n),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(tx_start),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output11 (.I(net12),
    .Z(tx));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(tx_busy));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload0 (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_208 ();
endmodule
