module configurable_carry_lookahead_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 INV_X16 _070_ (.A(net65),
    .ZN(_000_));
 INV_X1 _071_ (.A(net25),
    .ZN(_052_));
 INV_X16 _072_ (.A(net1),
    .ZN(_001_));
 INV_X1 _073_ (.A(net57),
    .ZN(_053_));
 INV_X4 _074_ (.A(net33),
    .ZN(_002_));
 INV_X1 _075_ (.A(_006_),
    .ZN(net68));
 INV_X1 _076_ (.A(_008_),
    .ZN(net69));
 INV_X1 _077_ (.A(_010_),
    .ZN(net70));
 INV_X1 _078_ (.A(_012_),
    .ZN(net71));
 INV_X1 _079_ (.A(_014_),
    .ZN(net72));
 INV_X1 _080_ (.A(_016_),
    .ZN(net73));
 INV_X1 _081_ (.A(_018_),
    .ZN(net74));
 INV_X1 _082_ (.A(_020_),
    .ZN(net75));
 INV_X1 _083_ (.A(_022_),
    .ZN(net76));
 INV_X1 _084_ (.A(_024_),
    .ZN(net77));
 INV_X1 _085_ (.A(_027_),
    .ZN(net78));
 INV_X1 _086_ (.A(_029_),
    .ZN(net79));
 INV_X1 _087_ (.A(_031_),
    .ZN(net80));
 INV_X1 _088_ (.A(_033_),
    .ZN(net81));
 INV_X1 _089_ (.A(_035_),
    .ZN(net82));
 INV_X1 _090_ (.A(_037_),
    .ZN(net83));
 INV_X1 _091_ (.A(_039_),
    .ZN(net84));
 INV_X1 _092_ (.A(_041_),
    .ZN(net85));
 INV_X1 _093_ (.A(_043_),
    .ZN(net86));
 INV_X1 _094_ (.A(_045_),
    .ZN(net87));
 INV_X1 _095_ (.A(_047_),
    .ZN(net88));
 INV_X1 _096_ (.A(_049_),
    .ZN(net89));
 INV_X1 _097_ (.A(_051_),
    .ZN(net90));
 INV_X1 _098_ (.A(_056_),
    .ZN(net91));
 INV_X1 _099_ (.A(_058_),
    .ZN(net92));
 INV_X1 _100_ (.A(_060_),
    .ZN(net93));
 INV_X1 _101_ (.A(_062_),
    .ZN(net94));
 INV_X1 _102_ (.A(_064_),
    .ZN(net95));
 INV_X1 _103_ (.A(_066_),
    .ZN(net96));
 INV_X1 _104_ (.A(_068_),
    .ZN(net97));
 INV_X1 _105_ (.A(_069_),
    .ZN(net98));
 INV_X2 _106_ (.A(_050_),
    .ZN(_054_));
 INV_X1 _107_ (.A(_055_),
    .ZN(net66));
 INV_X2 _108_ (.A(_003_),
    .ZN(_025_));
 FA_X1 _109_ (.A(_000_),
    .B(_001_),
    .CI(_002_),
    .CO(_003_),
    .S(net67));
 FA_X1 _110_ (.A(net2),
    .B(net34),
    .CI(_004_),
    .CO(_005_),
    .S(_006_));
 FA_X1 _111_ (.A(net3),
    .B(net35),
    .CI(_005_),
    .CO(_007_),
    .S(_008_));
 FA_X1 _112_ (.A(net4),
    .B(net36),
    .CI(_007_),
    .CO(_009_),
    .S(_010_));
 FA_X1 _113_ (.A(net5),
    .B(net37),
    .CI(_009_),
    .CO(_011_),
    .S(_012_));
 FA_X1 _114_ (.A(net6),
    .B(net38),
    .CI(_011_),
    .CO(_013_),
    .S(_014_));
 FA_X1 _115_ (.A(net7),
    .B(net39),
    .CI(_013_),
    .CO(_015_),
    .S(_016_));
 FA_X1 _116_ (.A(net8),
    .B(net40),
    .CI(_015_),
    .CO(_017_),
    .S(_018_));
 FA_X1 _117_ (.A(net9),
    .B(net41),
    .CI(_017_),
    .CO(_019_),
    .S(_020_));
 FA_X1 _118_ (.A(net10),
    .B(net42),
    .CI(_019_),
    .CO(_021_),
    .S(_022_));
 FA_X1 _119_ (.A(net11),
    .B(net43),
    .CI(_021_),
    .CO(_023_),
    .S(_024_));
 FA_X1 _120_ (.A(net12),
    .B(net44),
    .CI(_025_),
    .CO(_026_),
    .S(_027_));
 FA_X1 _121_ (.A(net13),
    .B(net45),
    .CI(_023_),
    .CO(_028_),
    .S(_029_));
 FA_X1 _122_ (.A(net14),
    .B(net46),
    .CI(_028_),
    .CO(_030_),
    .S(_031_));
 FA_X1 _123_ (.A(net15),
    .B(net47),
    .CI(_030_),
    .CO(_032_),
    .S(_033_));
 FA_X1 _124_ (.A(net16),
    .B(net48),
    .CI(_032_),
    .CO(_034_),
    .S(_035_));
 FA_X1 _125_ (.A(net17),
    .B(net49),
    .CI(_034_),
    .CO(_036_),
    .S(_037_));
 FA_X1 _126_ (.A(net18),
    .B(net50),
    .CI(_036_),
    .CO(_038_),
    .S(_039_));
 FA_X1 _127_ (.A(net19),
    .B(net51),
    .CI(_038_),
    .CO(_040_),
    .S(_041_));
 FA_X1 _128_ (.A(net20),
    .B(net52),
    .CI(_040_),
    .CO(_042_),
    .S(_043_));
 FA_X1 _129_ (.A(net21),
    .B(net53),
    .CI(_042_),
    .CO(_044_),
    .S(_045_));
 FA_X1 _130_ (.A(net22),
    .B(net54),
    .CI(_044_),
    .CO(_046_),
    .S(_047_));
 FA_X1 _131_ (.A(net23),
    .B(net55),
    .CI(_026_),
    .CO(_048_),
    .S(_049_));
 FA_X1 _132_ (.A(net24),
    .B(net56),
    .CI(_046_),
    .CO(_050_),
    .S(_051_));
 FA_X1 _133_ (.A(_052_),
    .B(_053_),
    .CI(_054_),
    .CO(_055_),
    .S(_056_));
 FA_X1 _134_ (.A(net26),
    .B(net58),
    .CI(_048_),
    .CO(_057_),
    .S(_058_));
 FA_X1 _135_ (.A(net27),
    .B(net59),
    .CI(_057_),
    .CO(_059_),
    .S(_060_));
 FA_X1 _136_ (.A(net28),
    .B(net60),
    .CI(_059_),
    .CO(_061_),
    .S(_062_));
 FA_X1 _137_ (.A(net29),
    .B(net61),
    .CI(_061_),
    .CO(_063_),
    .S(_064_));
 FA_X1 _138_ (.A(net30),
    .B(net62),
    .CI(_063_),
    .CO(_065_),
    .S(_066_));
 FA_X1 _139_ (.A(net31),
    .B(net63),
    .CI(_065_),
    .CO(_067_),
    .S(_068_));
 FA_X1 _140_ (.A(net32),
    .B(net64),
    .CI(_067_),
    .CO(_004_),
    .S(_069_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_43 ();
 BUF_X32 input1 (.A(a[0]),
    .Z(net1));
 BUF_X1 input2 (.A(a[10]),
    .Z(net2));
 BUF_X1 input3 (.A(a[11]),
    .Z(net3));
 BUF_X1 input4 (.A(a[12]),
    .Z(net4));
 BUF_X1 input5 (.A(a[13]),
    .Z(net5));
 BUF_X1 input6 (.A(a[14]),
    .Z(net6));
 BUF_X1 input7 (.A(a[15]),
    .Z(net7));
 BUF_X1 input8 (.A(a[16]),
    .Z(net8));
 BUF_X1 input9 (.A(a[17]),
    .Z(net9));
 BUF_X1 input10 (.A(a[18]),
    .Z(net10));
 BUF_X1 input11 (.A(a[19]),
    .Z(net11));
 BUF_X1 input12 (.A(a[1]),
    .Z(net12));
 BUF_X1 input13 (.A(a[20]),
    .Z(net13));
 BUF_X1 input14 (.A(a[21]),
    .Z(net14));
 BUF_X1 input15 (.A(a[22]),
    .Z(net15));
 BUF_X1 input16 (.A(a[23]),
    .Z(net16));
 BUF_X1 input17 (.A(a[24]),
    .Z(net17));
 BUF_X1 input18 (.A(a[25]),
    .Z(net18));
 BUF_X1 input19 (.A(a[26]),
    .Z(net19));
 BUF_X1 input20 (.A(a[27]),
    .Z(net20));
 BUF_X1 input21 (.A(a[28]),
    .Z(net21));
 BUF_X1 input22 (.A(a[29]),
    .Z(net22));
 BUF_X1 input23 (.A(a[2]),
    .Z(net23));
 BUF_X1 input24 (.A(a[30]),
    .Z(net24));
 BUF_X1 input25 (.A(a[31]),
    .Z(net25));
 BUF_X1 input26 (.A(a[3]),
    .Z(net26));
 BUF_X1 input27 (.A(a[4]),
    .Z(net27));
 BUF_X1 input28 (.A(a[5]),
    .Z(net28));
 BUF_X1 input29 (.A(a[6]),
    .Z(net29));
 BUF_X1 input30 (.A(a[7]),
    .Z(net30));
 BUF_X1 input31 (.A(a[8]),
    .Z(net31));
 BUF_X1 input32 (.A(a[9]),
    .Z(net32));
 BUF_X4 input33 (.A(b[0]),
    .Z(net33));
 BUF_X1 input34 (.A(b[10]),
    .Z(net34));
 BUF_X1 input35 (.A(b[11]),
    .Z(net35));
 BUF_X1 input36 (.A(b[12]),
    .Z(net36));
 BUF_X1 input37 (.A(b[13]),
    .Z(net37));
 BUF_X1 input38 (.A(b[14]),
    .Z(net38));
 BUF_X1 input39 (.A(b[15]),
    .Z(net39));
 BUF_X1 input40 (.A(b[16]),
    .Z(net40));
 BUF_X1 input41 (.A(b[17]),
    .Z(net41));
 BUF_X1 input42 (.A(b[18]),
    .Z(net42));
 BUF_X1 input43 (.A(b[19]),
    .Z(net43));
 BUF_X1 input44 (.A(b[1]),
    .Z(net44));
 BUF_X1 input45 (.A(b[20]),
    .Z(net45));
 BUF_X1 input46 (.A(b[21]),
    .Z(net46));
 BUF_X1 input47 (.A(b[22]),
    .Z(net47));
 BUF_X1 input48 (.A(b[23]),
    .Z(net48));
 BUF_X1 input49 (.A(b[24]),
    .Z(net49));
 BUF_X1 input50 (.A(b[25]),
    .Z(net50));
 BUF_X1 input51 (.A(b[26]),
    .Z(net51));
 BUF_X1 input52 (.A(b[27]),
    .Z(net52));
 BUF_X1 input53 (.A(b[28]),
    .Z(net53));
 BUF_X1 input54 (.A(b[29]),
    .Z(net54));
 BUF_X1 input55 (.A(b[2]),
    .Z(net55));
 BUF_X1 input56 (.A(b[30]),
    .Z(net56));
 BUF_X1 input57 (.A(b[31]),
    .Z(net57));
 BUF_X1 input58 (.A(b[3]),
    .Z(net58));
 BUF_X1 input59 (.A(b[4]),
    .Z(net59));
 BUF_X1 input60 (.A(b[5]),
    .Z(net60));
 BUF_X1 input61 (.A(b[6]),
    .Z(net61));
 BUF_X1 input62 (.A(b[7]),
    .Z(net62));
 BUF_X1 input63 (.A(b[8]),
    .Z(net63));
 BUF_X1 input64 (.A(b[9]),
    .Z(net64));
 BUF_X32 input65 (.A(cin),
    .Z(net65));
 BUF_X1 output66 (.A(net66),
    .Z(cout));
 BUF_X1 output67 (.A(net67),
    .Z(sum[0]));
 BUF_X1 output68 (.A(net68),
    .Z(sum[10]));
 BUF_X1 output69 (.A(net69),
    .Z(sum[11]));
 BUF_X1 output70 (.A(net70),
    .Z(sum[12]));
 BUF_X1 output71 (.A(net71),
    .Z(sum[13]));
 BUF_X1 output72 (.A(net72),
    .Z(sum[14]));
 BUF_X1 output73 (.A(net73),
    .Z(sum[15]));
 BUF_X1 output74 (.A(net74),
    .Z(sum[16]));
 BUF_X2 output75 (.A(net75),
    .Z(sum[17]));
 BUF_X1 output76 (.A(net76),
    .Z(sum[18]));
 BUF_X1 output77 (.A(net77),
    .Z(sum[19]));
 BUF_X1 output78 (.A(net78),
    .Z(sum[1]));
 BUF_X1 output79 (.A(net79),
    .Z(sum[20]));
 BUF_X2 output80 (.A(net80),
    .Z(sum[21]));
 BUF_X2 output81 (.A(net81),
    .Z(sum[22]));
 BUF_X1 output82 (.A(net82),
    .Z(sum[23]));
 BUF_X1 output83 (.A(net83),
    .Z(sum[24]));
 BUF_X1 output84 (.A(net84),
    .Z(sum[25]));
 BUF_X1 output85 (.A(net85),
    .Z(sum[26]));
 BUF_X1 output86 (.A(net86),
    .Z(sum[27]));
 BUF_X1 output87 (.A(net87),
    .Z(sum[28]));
 BUF_X1 output88 (.A(net88),
    .Z(sum[29]));
 BUF_X1 output89 (.A(net89),
    .Z(sum[2]));
 BUF_X1 output90 (.A(net90),
    .Z(sum[30]));
 BUF_X1 output91 (.A(net91),
    .Z(sum[31]));
 BUF_X1 output92 (.A(net92),
    .Z(sum[3]));
 BUF_X1 output93 (.A(net93),
    .Z(sum[4]));
 BUF_X1 output94 (.A(net94),
    .Z(sum[5]));
 BUF_X1 output95 (.A(net95),
    .Z(sum[6]));
 BUF_X1 output96 (.A(net96),
    .Z(sum[7]));
 BUF_X1 output97 (.A(net97),
    .Z(sum[8]));
 BUF_X1 output98 (.A(net98),
    .Z(sum[9]));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X4 FILLER_0_65 ();
 FILLCELL_X16 FILLER_0_72 ();
 FILLCELL_X2 FILLER_0_88 ();
 FILLCELL_X16 FILLER_0_96 ();
 FILLCELL_X4 FILLER_0_112 ();
 FILLCELL_X2 FILLER_0_116 ();
 FILLCELL_X1 FILLER_0_118 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X4 FILLER_1_129 ();
 FILLCELL_X1 FILLER_1_133 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X16 FILLER_2_129 ();
 FILLCELL_X1 FILLER_2_145 ();
 FILLCELL_X1 FILLER_2_162 ();
 FILLCELL_X2 FILLER_2_166 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X16 FILLER_3_97 ();
 FILLCELL_X4 FILLER_3_113 ();
 FILLCELL_X2 FILLER_3_117 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X16 FILLER_4_129 ();
 FILLCELL_X2 FILLER_4_145 ();
 FILLCELL_X1 FILLER_4_147 ();
 FILLCELL_X1 FILLER_4_151 ();
 FILLCELL_X1 FILLER_4_160 ();
 FILLCELL_X1 FILLER_5_22 ();
 FILLCELL_X32 FILLER_5_26 ();
 FILLCELL_X32 FILLER_5_58 ();
 FILLCELL_X32 FILLER_5_90 ();
 FILLCELL_X16 FILLER_5_122 ();
 FILLCELL_X4 FILLER_5_138 ();
 FILLCELL_X1 FILLER_5_161 ();
 FILLCELL_X2 FILLER_6_19 ();
 FILLCELL_X1 FILLER_6_21 ();
 FILLCELL_X16 FILLER_6_30 ();
 FILLCELL_X8 FILLER_6_46 ();
 FILLCELL_X4 FILLER_6_54 ();
 FILLCELL_X32 FILLER_6_60 ();
 FILLCELL_X32 FILLER_6_92 ();
 FILLCELL_X16 FILLER_6_124 ();
 FILLCELL_X2 FILLER_6_140 ();
 FILLCELL_X1 FILLER_6_142 ();
 FILLCELL_X32 FILLER_7_32 ();
 FILLCELL_X16 FILLER_7_64 ();
 FILLCELL_X4 FILLER_7_80 ();
 FILLCELL_X2 FILLER_7_84 ();
 FILLCELL_X1 FILLER_7_86 ();
 FILLCELL_X16 FILLER_7_103 ();
 FILLCELL_X4 FILLER_7_119 ();
 FILLCELL_X2 FILLER_7_123 ();
 FILLCELL_X4 FILLER_7_127 ();
 FILLCELL_X2 FILLER_7_131 ();
 FILLCELL_X1 FILLER_7_133 ();
 FILLCELL_X1 FILLER_7_156 ();
 FILLCELL_X1 FILLER_7_161 ();
 FILLCELL_X1 FILLER_7_167 ();
 FILLCELL_X1 FILLER_8_22 ();
 FILLCELL_X2 FILLER_8_26 ();
 FILLCELL_X8 FILLER_8_30 ();
 FILLCELL_X2 FILLER_8_38 ();
 FILLCELL_X1 FILLER_8_40 ();
 FILLCELL_X32 FILLER_8_57 ();
 FILLCELL_X32 FILLER_8_89 ();
 FILLCELL_X8 FILLER_8_121 ();
 FILLCELL_X2 FILLER_8_129 ();
 FILLCELL_X4 FILLER_8_135 ();
 FILLCELL_X2 FILLER_8_139 ();
 FILLCELL_X1 FILLER_8_141 ();
 FILLCELL_X2 FILLER_8_166 ();
 FILLCELL_X4 FILLER_9_4 ();
 FILLCELL_X4 FILLER_9_10 ();
 FILLCELL_X1 FILLER_9_17 ();
 FILLCELL_X32 FILLER_9_37 ();
 FILLCELL_X32 FILLER_9_69 ();
 FILLCELL_X32 FILLER_9_101 ();
 FILLCELL_X8 FILLER_9_133 ();
 FILLCELL_X2 FILLER_9_141 ();
 FILLCELL_X1 FILLER_9_164 ();
 FILLCELL_X4 FILLER_10_1 ();
 FILLCELL_X2 FILLER_10_8 ();
 FILLCELL_X1 FILLER_10_10 ();
 FILLCELL_X16 FILLER_10_14 ();
 FILLCELL_X2 FILLER_10_30 ();
 FILLCELL_X32 FILLER_10_35 ();
 FILLCELL_X32 FILLER_10_67 ();
 FILLCELL_X32 FILLER_10_99 ();
 FILLCELL_X16 FILLER_10_131 ();
 FILLCELL_X4 FILLER_10_147 ();
 FILLCELL_X2 FILLER_10_151 ();
 FILLCELL_X8 FILLER_10_156 ();
 FILLCELL_X1 FILLER_10_164 ();
 FILLCELL_X1 FILLER_11_4 ();
 FILLCELL_X32 FILLER_11_23 ();
 FILLCELL_X32 FILLER_11_55 ();
 FILLCELL_X32 FILLER_11_87 ();
 FILLCELL_X16 FILLER_11_119 ();
 FILLCELL_X4 FILLER_11_135 ();
 FILLCELL_X1 FILLER_11_139 ();
 FILLCELL_X1 FILLER_11_164 ();
 FILLCELL_X1 FILLER_12_7 ();
 FILLCELL_X32 FILLER_12_24 ();
 FILLCELL_X32 FILLER_12_56 ();
 FILLCELL_X32 FILLER_12_88 ();
 FILLCELL_X16 FILLER_12_120 ();
 FILLCELL_X8 FILLER_12_136 ();
 FILLCELL_X2 FILLER_13_10 ();
 FILLCELL_X1 FILLER_13_12 ();
 FILLCELL_X1 FILLER_13_18 ();
 FILLCELL_X32 FILLER_13_21 ();
 FILLCELL_X32 FILLER_13_53 ();
 FILLCELL_X32 FILLER_13_85 ();
 FILLCELL_X16 FILLER_13_117 ();
 FILLCELL_X8 FILLER_13_133 ();
 FILLCELL_X2 FILLER_13_163 ();
 FILLCELL_X4 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_5 ();
 FILLCELL_X1 FILLER_14_7 ();
 FILLCELL_X32 FILLER_14_27 ();
 FILLCELL_X32 FILLER_14_59 ();
 FILLCELL_X32 FILLER_14_91 ();
 FILLCELL_X8 FILLER_14_123 ();
 FILLCELL_X8 FILLER_14_147 ();
 FILLCELL_X32 FILLER_15_28 ();
 FILLCELL_X32 FILLER_15_60 ();
 FILLCELL_X32 FILLER_15_92 ();
 FILLCELL_X16 FILLER_15_124 ();
 FILLCELL_X4 FILLER_15_140 ();
 FILLCELL_X4 FILLER_16_4 ();
 FILLCELL_X32 FILLER_16_16 ();
 FILLCELL_X32 FILLER_16_48 ();
 FILLCELL_X32 FILLER_16_80 ();
 FILLCELL_X32 FILLER_16_112 ();
 FILLCELL_X8 FILLER_16_144 ();
 FILLCELL_X4 FILLER_16_152 ();
 FILLCELL_X4 FILLER_16_161 ();
 FILLCELL_X32 FILLER_17_17 ();
 FILLCELL_X32 FILLER_17_49 ();
 FILLCELL_X32 FILLER_17_81 ();
 FILLCELL_X16 FILLER_17_113 ();
 FILLCELL_X8 FILLER_17_129 ();
 FILLCELL_X4 FILLER_17_137 ();
 FILLCELL_X2 FILLER_17_141 ();
 FILLCELL_X2 FILLER_17_165 ();
 FILLCELL_X1 FILLER_17_167 ();
 FILLCELL_X4 FILLER_18_4 ();
 FILLCELL_X4 FILLER_18_11 ();
 FILLCELL_X1 FILLER_18_18 ();
 FILLCELL_X32 FILLER_18_35 ();
 FILLCELL_X32 FILLER_18_67 ();
 FILLCELL_X32 FILLER_18_99 ();
 FILLCELL_X8 FILLER_18_131 ();
 FILLCELL_X1 FILLER_18_139 ();
 FILLCELL_X1 FILLER_18_164 ();
 FILLCELL_X1 FILLER_19_9 ();
 FILLCELL_X2 FILLER_19_32 ();
 FILLCELL_X32 FILLER_19_36 ();
 FILLCELL_X16 FILLER_19_68 ();
 FILLCELL_X4 FILLER_19_84 ();
 FILLCELL_X8 FILLER_19_108 ();
 FILLCELL_X2 FILLER_19_116 ();
 FILLCELL_X32 FILLER_19_134 ();
 FILLCELL_X2 FILLER_19_166 ();
 FILLCELL_X1 FILLER_20_9 ();
 FILLCELL_X32 FILLER_20_32 ();
 FILLCELL_X16 FILLER_20_64 ();
 FILLCELL_X8 FILLER_20_80 ();
 FILLCELL_X2 FILLER_20_88 ();
 FILLCELL_X1 FILLER_20_90 ();
 FILLCELL_X4 FILLER_20_125 ();
 FILLCELL_X1 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_132 ();
 FILLCELL_X4 FILLER_20_164 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_17 ();
 FILLCELL_X2 FILLER_21_25 ();
 FILLCELL_X1 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_37 ();
 FILLCELL_X16 FILLER_21_69 ();
 FILLCELL_X4 FILLER_21_85 ();
 FILLCELL_X2 FILLER_21_89 ();
 FILLCELL_X1 FILLER_21_91 ();
 FILLCELL_X4 FILLER_21_116 ();
 FILLCELL_X1 FILLER_21_120 ();
 FILLCELL_X32 FILLER_21_133 ();
 FILLCELL_X2 FILLER_21_165 ();
 FILLCELL_X1 FILLER_21_167 ();
endmodule
