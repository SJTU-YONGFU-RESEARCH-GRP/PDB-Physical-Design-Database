module performance_counter (clear,
    clk,
    enable,
    rst_n,
    all_counts,
    count_value,
    counter_sel,
    event_inc);
 input clear;
 input clk;
 input enable;
 input rst_n;
 output [255:0] all_counts;
 output [31:0] count_value;
 input [7:0] counter_sel;
 input [7:0] event_inc;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire \prev_event_inc[0] ;
 wire \prev_event_inc[1] ;
 wire \prev_event_inc[2] ;
 wire \prev_event_inc[3] ;
 wire \prev_event_inc[4] ;
 wire \prev_event_inc[5] ;
 wire \prev_event_inc[6] ;
 wire \prev_event_inc[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 AOI21_X1 _1933_ (.A(_1197_),
    .B1(net223),
    .B2(_1198_),
    .ZN(_1268_));
 NAND2_X1 _1934_ (.A1(_1222_),
    .A2(net188),
    .ZN(_1269_));
 OAI21_X2 _1935_ (.A(_1268_),
    .B1(_1269_),
    .B2(_1224_),
    .ZN(_1270_));
 AOI21_X1 _1936_ (.A(_1169_),
    .B1(_0952_),
    .B2(_1227_),
    .ZN(_1271_));
 AOI221_X2 _1937_ (.A(_1209_),
    .B1(_1270_),
    .B2(_1271_),
    .C1(net38),
    .C2(_1229_),
    .ZN(_1272_));
 NOR2_X1 _1938_ (.A1(_1244_),
    .A2(net73),
    .ZN(_1273_));
 OR3_X1 _1939_ (.A1(_1196_),
    .A2(_1272_),
    .A3(_1273_),
    .ZN(_1274_));
 INV_X1 _1940_ (.A(net180),
    .ZN(_1275_));
 AOI221_X1 _1941_ (.A(_1266_),
    .B1(_1267_),
    .B2(_1274_),
    .C1(_1275_),
    .C2(_1234_),
    .ZN(net288));
 NOR3_X1 _1942_ (.A1(_1235_),
    .A2(net113),
    .A3(_0978_),
    .ZN(_1276_));
 AOI21_X2 _1943_ (.A(_1218_),
    .B1(_1660_),
    .B2(_1219_),
    .ZN(_1277_));
 AOI21_X1 _1944_ (.A(_1197_),
    .B1(_0700_),
    .B2(_1198_),
    .ZN(_1278_));
 NAND2_X1 _1945_ (.A1(_1222_),
    .A2(_1414_),
    .ZN(_1279_));
 OAI21_X1 _1946_ (.A(_1278_),
    .B1(_1279_),
    .B2(_1224_),
    .ZN(_1280_));
 INV_X1 _1947_ (.A(_0834_),
    .ZN(_1281_));
 AOI21_X1 _1948_ (.A(_1000_),
    .B1(_1281_),
    .B2(_1227_),
    .ZN(_1282_));
 AOI221_X2 _1949_ (.A(_1209_),
    .B1(_1280_),
    .B2(_1282_),
    .C1(_1359_),
    .C2(_1229_),
    .ZN(_1283_));
 NOR2_X1 _1950_ (.A1(_1244_),
    .A2(net43),
    .ZN(_1284_));
 OR3_X1 _1951_ (.A1(_1196_),
    .A2(_1283_),
    .A3(_1284_),
    .ZN(_1285_));
 AOI221_X2 _1952_ (.A(_1276_),
    .B1(_1277_),
    .B2(_1285_),
    .C1(_0532_),
    .C2(_1234_),
    .ZN(net289));
 NOR3_X1 _1953_ (.A1(_1235_),
    .A2(_0403_),
    .A3(_0978_),
    .ZN(_1286_));
 AOI21_X2 _1954_ (.A(_1218_),
    .B1(net79),
    .B2(_1219_),
    .ZN(_1287_));
 AOI21_X1 _1955_ (.A(_1197_),
    .B1(_0707_),
    .B2(_1198_),
    .ZN(_1288_));
 NAND2_X1 _1956_ (.A1(_1222_),
    .A2(_1415_),
    .ZN(_1289_));
 OAI21_X1 _1957_ (.A(_1288_),
    .B1(_1289_),
    .B2(_1224_),
    .ZN(_1290_));
 AOI21_X1 _1958_ (.A(_1000_),
    .B1(_0843_),
    .B2(_1227_),
    .ZN(_1291_));
 AOI221_X2 _1959_ (.A(_1209_),
    .B1(_1290_),
    .B2(_1291_),
    .C1(_1358_),
    .C2(_1229_),
    .ZN(_1292_));
 NOR2_X1 _1960_ (.A1(_1244_),
    .A2(net44),
    .ZN(_1293_));
 OR3_X1 _1961_ (.A1(_1196_),
    .A2(_1292_),
    .A3(_1293_),
    .ZN(_1294_));
 AOI221_X2 _1962_ (.A(_1286_),
    .B1(_1287_),
    .B2(_1294_),
    .C1(_0544_),
    .C2(_1234_),
    .ZN(net290));
 NOR3_X1 _1963_ (.A1(_1235_),
    .A2(net115),
    .A3(_0978_),
    .ZN(_1295_));
 AOI21_X2 _1964_ (.A(_1218_),
    .B1(net80),
    .B2(_1219_),
    .ZN(_1296_));
 AOI21_X1 _1965_ (.A(_1197_),
    .B1(_0712_),
    .B2(_1198_),
    .ZN(_1297_));
 NAND2_X1 _1966_ (.A1(_1222_),
    .A2(net219),
    .ZN(_1298_));
 OAI21_X1 _1967_ (.A(_1297_),
    .B1(_1298_),
    .B2(_1224_),
    .ZN(_1299_));
 INV_X1 _1968_ (.A(net229),
    .ZN(_1300_));
 AOI21_X1 _1969_ (.A(_1000_),
    .B1(_1300_),
    .B2(_1227_),
    .ZN(_1301_));
 AOI221_X2 _1970_ (.A(_1209_),
    .B1(_1299_),
    .B2(_1301_),
    .C1(_1368_),
    .C2(_1229_),
    .ZN(_1302_));
 NOR2_X1 _1971_ (.A1(_1244_),
    .A2(net45),
    .ZN(_1303_));
 OR3_X1 _1972_ (.A1(_1196_),
    .A2(_1302_),
    .A3(_1303_),
    .ZN(_1304_));
 AOI221_X2 _1973_ (.A(_1295_),
    .B1(_1296_),
    .B2(_1304_),
    .C1(_0546_),
    .C2(_1234_),
    .ZN(net291));
 NOR3_X2 _1974_ (.A1(_1235_),
    .A2(net116),
    .A3(_0978_),
    .ZN(_1305_));
 AOI21_X2 _1975_ (.A(_1218_),
    .B1(_0282_),
    .B2(_1219_),
    .ZN(_1306_));
 AOI21_X1 _1976_ (.A(_0990_),
    .B1(_0716_),
    .B2(_0992_),
    .ZN(_1307_));
 NAND2_X1 _1977_ (.A1(_1222_),
    .A2(_1419_),
    .ZN(_1308_));
 OAI21_X1 _1978_ (.A(_1307_),
    .B1(_1308_),
    .B2(_1224_),
    .ZN(_1309_));
 AOI21_X1 _1979_ (.A(_1000_),
    .B1(_0853_),
    .B2(_1227_),
    .ZN(_1310_));
 AOI221_X2 _1980_ (.A(_1209_),
    .B1(_1309_),
    .B2(_1310_),
    .C1(_1376_),
    .C2(_1229_),
    .ZN(_1311_));
 NOR2_X1 _1981_ (.A1(_1244_),
    .A2(_1539_),
    .ZN(_1312_));
 OR3_X1 _1982_ (.A1(_0984_),
    .A2(_1311_),
    .A3(_1312_),
    .ZN(_1313_));
 AOI221_X2 _1983_ (.A(_1305_),
    .B1(_1306_),
    .B2(_1313_),
    .C1(_0552_),
    .C2(_1234_),
    .ZN(net292));
 NOR3_X2 _1984_ (.A1(_1235_),
    .A2(_0412_),
    .A3(_0978_),
    .ZN(_1314_));
 AOI21_X2 _1985_ (.A(_1218_),
    .B1(_0288_),
    .B2(_1219_),
    .ZN(_1315_));
 AOI21_X1 _1986_ (.A(_0990_),
    .B1(_0720_),
    .B2(_0992_),
    .ZN(_1316_));
 NAND2_X1 _1987_ (.A1(_1222_),
    .A2(_1420_),
    .ZN(_1317_));
 OAI21_X1 _1988_ (.A(_1316_),
    .B1(_1317_),
    .B2(_1224_),
    .ZN(_1318_));
 INV_X1 _1989_ (.A(_0852_),
    .ZN(_1319_));
 AOI21_X1 _1990_ (.A(_1000_),
    .B1(_1319_),
    .B2(_1227_),
    .ZN(_1320_));
 AOI221_X2 _1991_ (.A(_0988_),
    .B1(_1318_),
    .B2(_1320_),
    .C1(_1380_),
    .C2(_1229_),
    .ZN(_1321_));
 NOR2_X1 _1992_ (.A1(_1244_),
    .A2(_1544_),
    .ZN(_1322_));
 OR3_X1 _1993_ (.A1(_0984_),
    .A2(_1321_),
    .A3(_1322_),
    .ZN(_1323_));
 AOI221_X2 _1994_ (.A(_1314_),
    .B1(_1315_),
    .B2(_1323_),
    .C1(_0555_),
    .C2(_1234_),
    .ZN(net293));
 NOR3_X2 _1995_ (.A1(_1235_),
    .A2(_0422_),
    .A3(_0978_),
    .ZN(_1324_));
 AOI21_X1 _1996_ (.A(_0982_),
    .B1(net83),
    .B2(_0987_),
    .ZN(_1325_));
 AOI21_X1 _1997_ (.A(_0990_),
    .B1(_0727_),
    .B2(_0992_),
    .ZN(_1326_));
 NAND2_X1 _1998_ (.A1(_0995_),
    .A2(net252),
    .ZN(_1327_));
 OAI21_X1 _1999_ (.A(_1326_),
    .B1(_1327_),
    .B2(_0993_),
    .ZN(_1328_));
 AOI21_X1 _2000_ (.A(_1000_),
    .B1(_0856_),
    .B2(_0991_),
    .ZN(_1329_));
 AOI221_X2 _2001_ (.A(_0988_),
    .B1(_1328_),
    .B2(_1329_),
    .C1(_1385_),
    .C2(_1001_),
    .ZN(_1330_));
 NOR2_X1 _2002_ (.A1(_1244_),
    .A2(_1549_),
    .ZN(_1331_));
 OR3_X1 _2003_ (.A1(_0984_),
    .A2(_1330_),
    .A3(_1331_),
    .ZN(_1332_));
 INV_X1 _2004_ (.A(_0558_),
    .ZN(_1333_));
 AOI221_X2 _2005_ (.A(_1324_),
    .B1(_1325_),
    .B2(_1332_),
    .C1(_1333_),
    .C2(_0979_),
    .ZN(net294));
 NOR3_X2 _2006_ (.A1(_0977_),
    .A2(net121),
    .A3(_0978_),
    .ZN(_1334_));
 AOI21_X1 _2007_ (.A(_0982_),
    .B1(net84),
    .B2(_0987_),
    .ZN(_1335_));
 AOI21_X1 _2008_ (.A(_0990_),
    .B1(_0731_),
    .B2(_0992_),
    .ZN(_1336_));
 NAND2_X1 _2009_ (.A1(_0995_),
    .A2(net263),
    .ZN(_1337_));
 OAI21_X1 _2010_ (.A(_1336_),
    .B1(_1337_),
    .B2(_0993_),
    .ZN(_1338_));
 INV_X1 _2011_ (.A(net234),
    .ZN(_1339_));
 AOI21_X1 _2012_ (.A(_1000_),
    .B1(_1339_),
    .B2(_0991_),
    .ZN(_1340_));
 AOI221_X2 _2013_ (.A(_0988_),
    .B1(_1338_),
    .B2(_1340_),
    .C1(_1389_),
    .C2(_1001_),
    .ZN(_1341_));
 NOR2_X1 _2014_ (.A1(_1007_),
    .A2(_1552_),
    .ZN(_1342_));
 OR3_X1 _2015_ (.A1(_0984_),
    .A2(_1341_),
    .A3(_1342_),
    .ZN(_1343_));
 AOI221_X2 _2016_ (.A(_1334_),
    .B1(_1335_),
    .B2(_1343_),
    .C1(_0563_),
    .C2(_0979_),
    .ZN(net295));
 BUF_X4 _2017_ (.A(clear),
    .Z(_1344_));
 INV_X4 _2018_ (.A(net7),
    .ZN(_1345_));
 NOR2_X1 _2019_ (.A1(_1344_),
    .A2(_1345_),
    .ZN(_1346_));
 BUF_X2 _2020_ (.A(_1346_),
    .Z(_1347_));
 CLKBUF_X3 _2021_ (.A(_1347_),
    .Z(_1348_));
 INV_X1 _2022_ (.A(\prev_event_inc[0] ),
    .ZN(_1349_));
 BUF_X4 _2023_ (.A(enable),
    .Z(_1350_));
 BUF_X8 _2024_ (.A(_1350_),
    .Z(_1351_));
 NAND3_X2 _2025_ (.A1(_1349_),
    .A2(net3),
    .A3(_1351_),
    .ZN(_1352_));
 MUX2_X1 _2026_ (.A(_0014_),
    .B(net8),
    .S(_1352_),
    .Z(_1353_));
 AND2_X1 _2027_ (.A1(_1348_),
    .A2(_1353_),
    .ZN(_0016_));
 INV_X4 _2028_ (.A(_1344_),
    .ZN(_1354_));
 NAND2_X2 _2029_ (.A1(_1354_),
    .A2(net7),
    .ZN(_1355_));
 BUF_X4 _2030_ (.A(_1355_),
    .Z(_1356_));
 CLKBUF_X3 _2031_ (.A(_1356_),
    .Z(_1357_));
 BUF_X2 _2032_ (.A(net9),
    .Z(_1358_));
 BUF_X2 _2033_ (.A(net262),
    .Z(_1359_));
 INV_X1 _2034_ (.A(_1359_),
    .ZN(_1360_));
 INV_X2 _2035_ (.A(\prev_event_inc[3] ),
    .ZN(_1361_));
 CLKBUF_X3 _2036_ (.A(event_inc[3]),
    .Z(_1362_));
 BUF_X2 _2037_ (.A(net261),
    .Z(_1363_));
 AND2_X1 _2038_ (.A1(_1363_),
    .A2(_1926_),
    .ZN(_1364_));
 NAND4_X4 _2039_ (.A1(_1351_),
    .A2(_1361_),
    .A3(_1362_),
    .A4(_1364_),
    .ZN(_1365_));
 NOR2_X1 _2040_ (.A1(_1360_),
    .A2(_1365_),
    .ZN(_1366_));
 XNOR2_X1 _2041_ (.A(_1358_),
    .B(_1366_),
    .ZN(_1367_));
 NOR2_X1 _2042_ (.A1(_1357_),
    .A2(_1367_),
    .ZN(_0017_));
 BUF_X2 _2043_ (.A(net10),
    .Z(_1368_));
 INV_X8 _2044_ (.A(_1350_),
    .ZN(_1369_));
 CLKBUF_X2 _2045_ (.A(net260),
    .Z(_1370_));
 NAND2_X1 _2046_ (.A1(_1370_),
    .A2(_1363_),
    .ZN(_1371_));
 NAND2_X2 _2047_ (.A1(_1362_),
    .A2(net259),
    .ZN(_1372_));
 NOR4_X4 _2048_ (.A1(_1369_),
    .A2(\prev_event_inc[3] ),
    .A3(_1371_),
    .A4(_1372_),
    .ZN(_1373_));
 NAND3_X1 _2049_ (.A1(_1359_),
    .A2(_1358_),
    .A3(_1373_),
    .ZN(_1374_));
 XOR2_X1 _2050_ (.A(_1368_),
    .B(_1374_),
    .Z(_1375_));
 NOR2_X1 _2051_ (.A1(_1357_),
    .A2(_1375_),
    .ZN(_0018_));
 CLKBUF_X2 _2052_ (.A(net11),
    .Z(_1376_));
 NAND3_X1 _2053_ (.A1(_1359_),
    .A2(_1358_),
    .A3(_1368_),
    .ZN(_1377_));
 NOR2_X1 _2054_ (.A1(_1365_),
    .A2(_1377_),
    .ZN(_1378_));
 XNOR2_X1 _2055_ (.A(_1376_),
    .B(_1378_),
    .ZN(_1379_));
 NOR2_X1 _2056_ (.A1(_1357_),
    .A2(_1379_),
    .ZN(_0019_));
 CLKBUF_X2 _2057_ (.A(net12),
    .Z(_1380_));
 INV_X1 _2058_ (.A(_1380_),
    .ZN(_1381_));
 AND4_X2 _2059_ (.A1(_1359_),
    .A2(_1358_),
    .A3(_1368_),
    .A4(_1376_),
    .ZN(_1382_));
 NAND2_X1 _2060_ (.A1(_1373_),
    .A2(_1382_),
    .ZN(_1383_));
 XNOR2_X1 _2061_ (.A(_1381_),
    .B(_1383_),
    .ZN(_1384_));
 NOR2_X1 _2062_ (.A1(_1357_),
    .A2(_1384_),
    .ZN(_0020_));
 BUF_X2 _2063_ (.A(net13),
    .Z(_1385_));
 NAND4_X2 _2064_ (.A1(_1359_),
    .A2(_1358_),
    .A3(_1368_),
    .A4(_1376_),
    .ZN(_1386_));
 NOR3_X1 _2065_ (.A1(_1381_),
    .A2(_1365_),
    .A3(_1386_),
    .ZN(_1387_));
 XNOR2_X1 _2066_ (.A(_1385_),
    .B(_1387_),
    .ZN(_1388_));
 NOR2_X1 _2067_ (.A1(_1357_),
    .A2(_1388_),
    .ZN(_0021_));
 BUF_X2 _2068_ (.A(net14),
    .Z(_1389_));
 NAND4_X1 _2069_ (.A1(_1380_),
    .A2(_1385_),
    .A3(_1373_),
    .A4(_1382_),
    .ZN(_1390_));
 XOR2_X1 _2070_ (.A(_1389_),
    .B(_1390_),
    .Z(_1391_));
 NOR2_X1 _2071_ (.A1(_1357_),
    .A2(_1391_),
    .ZN(_0022_));
 NAND3_X1 _2072_ (.A1(_1380_),
    .A2(_1385_),
    .A3(_1389_),
    .ZN(_1392_));
 NOR3_X1 _2073_ (.A1(_1365_),
    .A2(_1386_),
    .A3(_1392_),
    .ZN(_1393_));
 XNOR2_X1 _2074_ (.A(net15),
    .B(_1393_),
    .ZN(_1394_));
 NOR2_X1 _2075_ (.A1(_1357_),
    .A2(_1394_),
    .ZN(_0023_));
 BUF_X2 _2076_ (.A(net16),
    .Z(_1395_));
 AND4_X2 _2077_ (.A1(_1380_),
    .A2(_1385_),
    .A3(_1389_),
    .A4(net15),
    .ZN(_1396_));
 NAND3_X1 _2078_ (.A1(_1373_),
    .A2(_1382_),
    .A3(_1396_),
    .ZN(_1397_));
 XOR2_X1 _2079_ (.A(_1395_),
    .B(_1397_),
    .Z(_1398_));
 NOR2_X1 _2080_ (.A1(_1357_),
    .A2(_1398_),
    .ZN(_0024_));
 BUF_X2 _2081_ (.A(net17),
    .Z(_1399_));
 NAND2_X1 _2082_ (.A1(_1395_),
    .A2(_1396_),
    .ZN(_1400_));
 NOR3_X1 _2083_ (.A1(_1365_),
    .A2(_1386_),
    .A3(_1400_),
    .ZN(_1401_));
 XNOR2_X1 _2084_ (.A(_1399_),
    .B(_1401_),
    .ZN(_1402_));
 NOR2_X1 _2085_ (.A1(_1357_),
    .A2(_1402_),
    .ZN(_0025_));
 CLKBUF_X2 _2086_ (.A(net18),
    .Z(_1403_));
 INV_X1 _2087_ (.A(_1403_),
    .ZN(_1404_));
 NAND3_X1 _2088_ (.A1(_1350_),
    .A2(_1361_),
    .A3(_1362_),
    .ZN(_1405_));
 NAND2_X1 _2089_ (.A1(net259),
    .A2(_1370_),
    .ZN(_1406_));
 NAND4_X1 _2090_ (.A1(_1363_),
    .A2(_1395_),
    .A3(_1399_),
    .A4(_1396_),
    .ZN(_1407_));
 OR4_X1 _2091_ (.A1(_1405_),
    .A2(_1406_),
    .A3(_1386_),
    .A4(_1407_),
    .ZN(_1408_));
 BUF_X4 _2092_ (.A(_1408_),
    .Z(_1409_));
 XNOR2_X1 _2093_ (.A(_1404_),
    .B(_1409_),
    .ZN(_1410_));
 NOR2_X1 _2094_ (.A1(_1357_),
    .A2(_1410_),
    .ZN(_0026_));
 CLKBUF_X3 _2095_ (.A(_1356_),
    .Z(_1411_));
 INV_X1 _2096_ (.A(_1931_),
    .ZN(_1412_));
 NAND2_X2 _2097_ (.A1(net3),
    .A2(_1350_),
    .ZN(_1413_));
 BUF_X2 _2098_ (.A(net197),
    .Z(_1414_));
 BUF_X2 _2099_ (.A(net208),
    .Z(_1415_));
 NAND4_X4 _2100_ (.A1(net186),
    .A2(_1414_),
    .A3(_1415_),
    .A4(net219),
    .ZN(_1416_));
 NOR4_X4 _2101_ (.A1(\prev_event_inc[0] ),
    .A2(_1412_),
    .A3(_1413_),
    .A4(_1416_),
    .ZN(_1417_));
 BUF_X4 _2102_ (.A(_1417_),
    .Z(_1418_));
 BUF_X2 _2103_ (.A(net230),
    .Z(_1419_));
 CLKBUF_X2 _2104_ (.A(net241),
    .Z(_1420_));
 AND4_X1 _2105_ (.A1(_1419_),
    .A2(_1420_),
    .A3(net252),
    .A4(net263),
    .ZN(_1421_));
 NAND2_X1 _2106_ (.A1(_1418_),
    .A2(_1421_),
    .ZN(_1422_));
 XOR2_X1 _2107_ (.A(net19),
    .B(_1422_),
    .Z(_1423_));
 NOR2_X1 _2108_ (.A1(_1411_),
    .A2(_1423_),
    .ZN(_0027_));
 CLKBUF_X2 _2109_ (.A(net20),
    .Z(_1424_));
 NAND2_X4 _2110_ (.A1(_1382_),
    .A2(_1396_),
    .ZN(_1425_));
 AND4_X1 _2111_ (.A1(_1363_),
    .A2(_1395_),
    .A3(_1399_),
    .A4(_1926_),
    .ZN(_1426_));
 NAND4_X4 _2112_ (.A1(_1351_),
    .A2(_1361_),
    .A3(_1362_),
    .A4(_1426_),
    .ZN(_1427_));
 NOR3_X1 _2113_ (.A1(_1404_),
    .A2(_1425_),
    .A3(_1427_),
    .ZN(_1428_));
 XNOR2_X1 _2114_ (.A(_1424_),
    .B(_1428_),
    .ZN(_1429_));
 NOR2_X1 _2115_ (.A1(_1411_),
    .A2(_1429_),
    .ZN(_0028_));
 NAND4_X2 _2116_ (.A1(_1370_),
    .A2(_1363_),
    .A3(_1395_),
    .A4(_1399_),
    .ZN(_1430_));
 NOR4_X4 _2117_ (.A1(_1369_),
    .A2(\prev_event_inc[3] ),
    .A3(_1372_),
    .A4(_1430_),
    .ZN(_1431_));
 AND2_X1 _2118_ (.A1(_1382_),
    .A2(_1396_),
    .ZN(_1432_));
 NAND4_X1 _2119_ (.A1(_1403_),
    .A2(_1424_),
    .A3(_1431_),
    .A4(_1432_),
    .ZN(_1433_));
 XOR2_X1 _2120_ (.A(net21),
    .B(_1433_),
    .Z(_1434_));
 NOR2_X1 _2121_ (.A1(_1411_),
    .A2(_1434_),
    .ZN(_0029_));
 NAND3_X1 _2122_ (.A1(_1403_),
    .A2(_1424_),
    .A3(net21),
    .ZN(_1435_));
 NOR3_X1 _2123_ (.A1(_1425_),
    .A2(_1427_),
    .A3(_1435_),
    .ZN(_1436_));
 XNOR2_X1 _2124_ (.A(net22),
    .B(_1436_),
    .ZN(_1437_));
 NOR2_X1 _2125_ (.A1(_1411_),
    .A2(_1437_),
    .ZN(_0030_));
 CLKBUF_X2 _2126_ (.A(net23),
    .Z(_1438_));
 AND4_X1 _2127_ (.A1(_1403_),
    .A2(_1424_),
    .A3(net21),
    .A4(net22),
    .ZN(_1439_));
 BUF_X2 _2128_ (.A(_1439_),
    .Z(_1440_));
 NAND3_X1 _2129_ (.A1(_1431_),
    .A2(_1432_),
    .A3(_1440_),
    .ZN(_1441_));
 XOR2_X1 _2130_ (.A(_1438_),
    .B(_1441_),
    .Z(_1442_));
 NOR2_X1 _2131_ (.A1(_1411_),
    .A2(_1442_),
    .ZN(_0031_));
 CLKBUF_X2 _2132_ (.A(net24),
    .Z(_1443_));
 NAND2_X1 _2133_ (.A1(_1438_),
    .A2(_1440_),
    .ZN(_1444_));
 NOR3_X1 _2134_ (.A1(_1425_),
    .A2(_1427_),
    .A3(_1444_),
    .ZN(_1445_));
 XNOR2_X1 _2135_ (.A(_1443_),
    .B(_1445_),
    .ZN(_1446_));
 NOR2_X1 _2136_ (.A1(_1411_),
    .A2(_1446_),
    .ZN(_0032_));
 BUF_X4 _2137_ (.A(_1355_),
    .Z(_1447_));
 BUF_X4 _2138_ (.A(_1447_),
    .Z(_1448_));
 BUF_X1 _2139_ (.A(net25),
    .Z(_1449_));
 NAND3_X1 _2140_ (.A1(_1438_),
    .A2(_1443_),
    .A3(_1440_),
    .ZN(_1450_));
 OAI21_X1 _2141_ (.A(_1449_),
    .B1(_1409_),
    .B2(_1450_),
    .ZN(_1451_));
 OR3_X1 _2142_ (.A1(_1449_),
    .A2(_1409_),
    .A3(_1450_),
    .ZN(_1452_));
 AOI21_X1 _2143_ (.A(_1448_),
    .B1(_1451_),
    .B2(_1452_),
    .ZN(_0033_));
 NAND4_X1 _2144_ (.A1(_1438_),
    .A2(_1443_),
    .A3(_1449_),
    .A4(_1440_),
    .ZN(_1453_));
 NOR3_X1 _2145_ (.A1(_1425_),
    .A2(_1427_),
    .A3(_1453_),
    .ZN(_1454_));
 XNOR2_X1 _2146_ (.A(net26),
    .B(_1454_),
    .ZN(_1455_));
 NOR2_X1 _2147_ (.A1(_1411_),
    .A2(_1455_),
    .ZN(_0034_));
 BUF_X2 _2148_ (.A(net27),
    .Z(_1456_));
 AND4_X1 _2149_ (.A1(_1438_),
    .A2(_1443_),
    .A3(_1449_),
    .A4(net26),
    .ZN(_1457_));
 AND2_X1 _2150_ (.A1(_1440_),
    .A2(_1457_),
    .ZN(_1458_));
 NAND3_X1 _2151_ (.A1(_1431_),
    .A2(_1432_),
    .A3(_1458_),
    .ZN(_1459_));
 XOR2_X1 _2152_ (.A(_1456_),
    .B(_1459_),
    .Z(_1460_));
 NOR2_X1 _2153_ (.A1(_1411_),
    .A2(_1460_),
    .ZN(_0035_));
 NAND3_X1 _2154_ (.A1(_1456_),
    .A2(_1440_),
    .A3(_1457_),
    .ZN(_1461_));
 NOR3_X1 _2155_ (.A1(_1425_),
    .A2(_1427_),
    .A3(_1461_),
    .ZN(_1462_));
 XNOR2_X1 _2156_ (.A(net28),
    .B(_1462_),
    .ZN(_1463_));
 NOR2_X1 _2157_ (.A1(_1411_),
    .A2(_1463_),
    .ZN(_0036_));
 BUF_X2 _2158_ (.A(net29),
    .Z(_1464_));
 NAND4_X4 _2159_ (.A1(_1456_),
    .A2(net28),
    .A3(_1440_),
    .A4(_1457_),
    .ZN(_1465_));
 OAI21_X1 _2160_ (.A(_1464_),
    .B1(_1409_),
    .B2(_1465_),
    .ZN(_1466_));
 OR3_X1 _2161_ (.A1(_1464_),
    .A2(_1409_),
    .A3(_1465_),
    .ZN(_1467_));
 AOI21_X1 _2162_ (.A(_1448_),
    .B1(_1466_),
    .B2(_1467_),
    .ZN(_0037_));
 NAND2_X2 _2163_ (.A1(net8),
    .A2(net119),
    .ZN(_1468_));
 NOR4_X4 _2164_ (.A1(\prev_event_inc[0] ),
    .A2(_1413_),
    .A3(_1416_),
    .A4(_1468_),
    .ZN(_1469_));
 BUF_X4 _2165_ (.A(_1469_),
    .Z(_1470_));
 NAND3_X1 _2166_ (.A1(net19),
    .A2(_1421_),
    .A3(_1470_),
    .ZN(_1471_));
 XOR2_X1 _2167_ (.A(net30),
    .B(_1471_),
    .Z(_1472_));
 NOR2_X1 _2168_ (.A1(_1411_),
    .A2(_1472_),
    .ZN(_0038_));
 BUF_X2 _2169_ (.A(net31),
    .Z(_1473_));
 CLKBUF_X3 _2170_ (.A(_1355_),
    .Z(_1474_));
 NOR2_X1 _2171_ (.A1(_1473_),
    .A2(_1474_),
    .ZN(_1475_));
 AND2_X1 _2172_ (.A1(_1473_),
    .A2(_1347_),
    .ZN(_1476_));
 NOR3_X2 _2173_ (.A1(_1425_),
    .A2(_1427_),
    .A3(_1465_),
    .ZN(_1477_));
 NAND2_X1 _2174_ (.A1(_1464_),
    .A2(_1477_),
    .ZN(_1478_));
 MUX2_X1 _2175_ (.A(_1475_),
    .B(_1476_),
    .S(_1478_),
    .Z(_0039_));
 CLKBUF_X2 _2176_ (.A(net32),
    .Z(_1479_));
 AND2_X1 _2177_ (.A1(_1479_),
    .A2(_1347_),
    .ZN(_1480_));
 NOR2_X1 _2178_ (.A1(_1479_),
    .A2(_1447_),
    .ZN(_1481_));
 NAND2_X1 _2179_ (.A1(_1464_),
    .A2(_1473_),
    .ZN(_1482_));
 NOR3_X1 _2180_ (.A1(_1409_),
    .A2(_1465_),
    .A3(_1482_),
    .ZN(_1483_));
 MUX2_X1 _2181_ (.A(_1480_),
    .B(_1481_),
    .S(_1483_),
    .Z(_0040_));
 CLKBUF_X3 _2182_ (.A(_1356_),
    .Z(_1484_));
 NAND3_X1 _2183_ (.A1(_1464_),
    .A2(_1473_),
    .A3(_1479_),
    .ZN(_1485_));
 NOR4_X1 _2184_ (.A1(_1425_),
    .A2(_1427_),
    .A3(_1465_),
    .A4(_1485_),
    .ZN(_1486_));
 XNOR2_X1 _2185_ (.A(net33),
    .B(_1486_),
    .ZN(_1487_));
 NOR2_X1 _2186_ (.A1(_1484_),
    .A2(_1487_),
    .ZN(_0041_));
 INV_X1 _2187_ (.A(net34),
    .ZN(_1488_));
 NOR2_X1 _2188_ (.A1(_1488_),
    .A2(_1474_),
    .ZN(_1489_));
 CLKBUF_X3 _2189_ (.A(_1355_),
    .Z(_1490_));
 NOR2_X1 _2190_ (.A1(net34),
    .A2(_1490_),
    .ZN(_1491_));
 NAND4_X2 _2191_ (.A1(_1464_),
    .A2(_1473_),
    .A3(_1479_),
    .A4(net33),
    .ZN(_1492_));
 NOR3_X1 _2192_ (.A1(_1409_),
    .A2(_1465_),
    .A3(_1492_),
    .ZN(_1493_));
 MUX2_X1 _2193_ (.A(_1489_),
    .B(_1491_),
    .S(_1493_),
    .Z(_0042_));
 CLKBUF_X2 _2194_ (.A(net35),
    .Z(_1494_));
 NOR2_X1 _2195_ (.A1(_1494_),
    .A2(_1474_),
    .ZN(_1495_));
 AND2_X1 _2196_ (.A1(_1494_),
    .A2(_1347_),
    .ZN(_1496_));
 NOR2_X2 _2197_ (.A1(_1488_),
    .A2(_1492_),
    .ZN(_1497_));
 NAND2_X1 _2198_ (.A1(_1477_),
    .A2(_1497_),
    .ZN(_1498_));
 MUX2_X1 _2199_ (.A(_1495_),
    .B(_1496_),
    .S(_1498_),
    .Z(_0043_));
 CLKBUF_X2 _2200_ (.A(net36),
    .Z(_1499_));
 AND2_X1 _2201_ (.A1(_1499_),
    .A2(_1346_),
    .ZN(_1500_));
 NOR2_X1 _2202_ (.A1(_1499_),
    .A2(_1490_),
    .ZN(_1501_));
 NAND2_X1 _2203_ (.A1(_1494_),
    .A2(_1497_),
    .ZN(_1502_));
 NOR3_X1 _2204_ (.A1(_1409_),
    .A2(_1465_),
    .A3(_1502_),
    .ZN(_1503_));
 MUX2_X1 _2205_ (.A(_1500_),
    .B(_1501_),
    .S(_1503_),
    .Z(_0044_));
 NOR2_X1 _2206_ (.A1(net37),
    .A2(_1474_),
    .ZN(_1504_));
 AND2_X1 _2207_ (.A1(net37),
    .A2(_1347_),
    .ZN(_1505_));
 NAND4_X1 _2208_ (.A1(_1494_),
    .A2(_1499_),
    .A3(_1477_),
    .A4(_1497_),
    .ZN(_1506_));
 MUX2_X1 _2209_ (.A(_1504_),
    .B(_1505_),
    .S(_1506_),
    .Z(_0045_));
 AND2_X1 _2210_ (.A1(net38),
    .A2(_1346_),
    .ZN(_1507_));
 NOR2_X1 _2211_ (.A1(net38),
    .A2(_1490_),
    .ZN(_1508_));
 NAND4_X1 _2212_ (.A1(_1494_),
    .A2(_1499_),
    .A3(net37),
    .A4(_1497_),
    .ZN(_1509_));
 NOR3_X1 _2213_ (.A1(_1409_),
    .A2(_1465_),
    .A3(_1509_),
    .ZN(_1510_));
 MUX2_X1 _2214_ (.A(_1507_),
    .B(_1508_),
    .S(_1510_),
    .Z(_0046_));
 BUF_X4 _2215_ (.A(_1351_),
    .Z(_1511_));
 INV_X1 _2216_ (.A(\prev_event_inc[4] ),
    .ZN(_1512_));
 CLKBUF_X2 _2217_ (.A(event_inc[4]),
    .Z(_1513_));
 NAND3_X1 _2218_ (.A1(_1511_),
    .A2(_1512_),
    .A3(_1513_),
    .ZN(_1514_));
 MUX2_X1 _2219_ (.A(_0006_),
    .B(net39),
    .S(_1514_),
    .Z(_1515_));
 AND2_X1 _2220_ (.A1(_1348_),
    .A2(_1515_),
    .ZN(_0047_));
 MUX2_X1 _2221_ (.A(_0007_),
    .B(net40),
    .S(_1514_),
    .Z(_1516_));
 AND2_X1 _2222_ (.A1(_1348_),
    .A2(_1516_),
    .ZN(_0048_));
 BUF_X2 _2223_ (.A(net41),
    .Z(_1517_));
 AND3_X1 _2224_ (.A1(net19),
    .A2(net30),
    .A3(_1421_),
    .ZN(_1518_));
 CLKBUF_X3 _2225_ (.A(_1518_),
    .Z(_1519_));
 BUF_X4 _2226_ (.A(_1519_),
    .Z(_1520_));
 NAND2_X1 _2227_ (.A1(_1418_),
    .A2(_1520_),
    .ZN(_1521_));
 XOR2_X1 _2228_ (.A(_1517_),
    .B(_1521_),
    .Z(_1522_));
 NOR2_X1 _2229_ (.A1(_1484_),
    .A2(_1522_),
    .ZN(_0049_));
 BUF_X2 _2230_ (.A(net42),
    .Z(_1523_));
 AND2_X1 _2231_ (.A1(_1513_),
    .A2(_1927_),
    .ZN(_1524_));
 AND3_X1 _2232_ (.A1(_1351_),
    .A2(_1512_),
    .A3(_1524_),
    .ZN(_1525_));
 XNOR2_X1 _2233_ (.A(_1523_),
    .B(_1525_),
    .ZN(_1526_));
 NOR2_X1 _2234_ (.A1(_1484_),
    .A2(_1526_),
    .ZN(_0050_));
 AND2_X1 _2235_ (.A1(net39),
    .A2(net40),
    .ZN(_1527_));
 AND4_X2 _2236_ (.A1(_1350_),
    .A2(_1512_),
    .A3(_1513_),
    .A4(_1527_),
    .ZN(_1528_));
 NAND2_X1 _2237_ (.A1(_1523_),
    .A2(_1528_),
    .ZN(_1529_));
 XOR2_X1 _2238_ (.A(net43),
    .B(_1529_),
    .Z(_1530_));
 NOR2_X1 _2239_ (.A1(_1484_),
    .A2(_1530_),
    .ZN(_0051_));
 NAND3_X1 _2240_ (.A1(_1351_),
    .A2(_1512_),
    .A3(_1524_),
    .ZN(_1531_));
 NAND2_X1 _2241_ (.A1(_1523_),
    .A2(net43),
    .ZN(_1532_));
 NOR2_X1 _2242_ (.A1(_1531_),
    .A2(_1532_),
    .ZN(_1533_));
 XNOR2_X1 _2243_ (.A(net44),
    .B(_1533_),
    .ZN(_1534_));
 NOR2_X1 _2244_ (.A1(_1484_),
    .A2(_1534_),
    .ZN(_0052_));
 INV_X1 _2245_ (.A(net44),
    .ZN(_1535_));
 NAND4_X2 _2246_ (.A1(_1350_),
    .A2(_1512_),
    .A3(_1513_),
    .A4(_1527_),
    .ZN(_1536_));
 NOR3_X1 _2247_ (.A1(_1535_),
    .A2(_1536_),
    .A3(_1532_),
    .ZN(_1537_));
 XNOR2_X1 _2248_ (.A(net45),
    .B(_1537_),
    .ZN(_1538_));
 NOR2_X1 _2249_ (.A1(_1484_),
    .A2(_1538_),
    .ZN(_0053_));
 CLKBUF_X3 _2250_ (.A(net46),
    .Z(_1539_));
 AND4_X1 _2251_ (.A1(_1523_),
    .A2(net43),
    .A3(net44),
    .A4(net45),
    .ZN(_1540_));
 AND4_X1 _2252_ (.A1(_1350_),
    .A2(_1512_),
    .A3(_1524_),
    .A4(_1540_),
    .ZN(_1541_));
 BUF_X2 _2253_ (.A(_1541_),
    .Z(_1542_));
 XNOR2_X1 _2254_ (.A(_1539_),
    .B(_1542_),
    .ZN(_1543_));
 NOR2_X1 _2255_ (.A1(_1484_),
    .A2(_1543_),
    .ZN(_0054_));
 CLKBUF_X2 _2256_ (.A(net47),
    .Z(_1544_));
 NAND2_X2 _2257_ (.A1(_1539_),
    .A2(_1540_),
    .ZN(_1545_));
 OR2_X1 _2258_ (.A1(_1536_),
    .A2(_1545_),
    .ZN(_1546_));
 BUF_X2 _2259_ (.A(_1546_),
    .Z(_1547_));
 XOR2_X1 _2260_ (.A(_1544_),
    .B(_1547_),
    .Z(_1548_));
 NOR2_X1 _2261_ (.A1(_1484_),
    .A2(_1548_),
    .ZN(_0055_));
 BUF_X1 _2262_ (.A(net48),
    .Z(_1549_));
 NAND3_X1 _2263_ (.A1(_1539_),
    .A2(_1544_),
    .A3(_1542_),
    .ZN(_1550_));
 XOR2_X1 _2264_ (.A(_1549_),
    .B(_1550_),
    .Z(_1551_));
 NOR2_X1 _2265_ (.A1(_1484_),
    .A2(_1551_),
    .ZN(_0056_));
 BUF_X2 _2266_ (.A(net49),
    .Z(_1552_));
 NAND2_X1 _2267_ (.A1(_1544_),
    .A2(_1549_),
    .ZN(_1553_));
 OAI21_X1 _2268_ (.A(_1552_),
    .B1(_1547_),
    .B2(_1553_),
    .ZN(_1554_));
 OR3_X1 _2269_ (.A1(_1552_),
    .A2(_1547_),
    .A3(_1553_),
    .ZN(_1555_));
 AOI21_X1 _2270_ (.A(_1448_),
    .B1(_1554_),
    .B2(_1555_),
    .ZN(_0057_));
 INV_X1 _2271_ (.A(_1552_),
    .ZN(_1556_));
 NOR4_X1 _2272_ (.A1(_1556_),
    .A2(_1531_),
    .A3(_1545_),
    .A4(_1553_),
    .ZN(_1557_));
 XNOR2_X1 _2273_ (.A(net50),
    .B(_1557_),
    .ZN(_1558_));
 NOR2_X1 _2274_ (.A1(_1484_),
    .A2(_1558_),
    .ZN(_0058_));
 CLKBUF_X3 _2275_ (.A(_1355_),
    .Z(_1559_));
 CLKBUF_X3 _2276_ (.A(_1559_),
    .Z(_1560_));
 BUF_X2 _2277_ (.A(net51),
    .Z(_1561_));
 AND4_X2 _2278_ (.A1(_1544_),
    .A2(_1549_),
    .A3(_1552_),
    .A4(net50),
    .ZN(_1562_));
 AND4_X1 _2279_ (.A1(_1539_),
    .A2(_1528_),
    .A3(_1540_),
    .A4(_1562_),
    .ZN(_1563_));
 XNOR2_X1 _2280_ (.A(_1561_),
    .B(_1563_),
    .ZN(_1564_));
 NOR2_X1 _2281_ (.A1(_1560_),
    .A2(_1564_),
    .ZN(_0059_));
 BUF_X2 _2282_ (.A(net52),
    .Z(_1565_));
 NAND3_X1 _2283_ (.A1(_1517_),
    .A2(_1470_),
    .A3(_1520_),
    .ZN(_1566_));
 XOR2_X1 _2284_ (.A(_1565_),
    .B(_1566_),
    .Z(_1567_));
 NOR2_X1 _2285_ (.A1(_1560_),
    .A2(_1567_),
    .ZN(_0060_));
 CLKBUF_X2 _2286_ (.A(net53),
    .Z(_1568_));
 NAND4_X1 _2287_ (.A1(_1539_),
    .A2(_1561_),
    .A3(_1542_),
    .A4(_1562_),
    .ZN(_1569_));
 XOR2_X1 _2288_ (.A(_1568_),
    .B(_1569_),
    .Z(_1570_));
 NOR2_X1 _2289_ (.A1(_1560_),
    .A2(_1570_),
    .ZN(_0061_));
 BUF_X1 _2290_ (.A(net54),
    .Z(_1571_));
 NAND3_X1 _2291_ (.A1(_1561_),
    .A2(_1568_),
    .A3(_1562_),
    .ZN(_1572_));
 OAI21_X1 _2292_ (.A(_1571_),
    .B1(_1547_),
    .B2(_1572_),
    .ZN(_1573_));
 OR3_X1 _2293_ (.A1(_1571_),
    .A2(_1547_),
    .A3(_1572_),
    .ZN(_1574_));
 AOI21_X1 _2294_ (.A(_1448_),
    .B1(_1573_),
    .B2(_1574_),
    .ZN(_0062_));
 INV_X1 _2295_ (.A(_1571_),
    .ZN(_1575_));
 OR4_X1 _2296_ (.A1(_1575_),
    .A2(_1531_),
    .A3(_1545_),
    .A4(_1572_),
    .ZN(_1576_));
 XOR2_X1 _2297_ (.A(net55),
    .B(_1576_),
    .Z(_1577_));
 NOR2_X1 _2298_ (.A1(_1560_),
    .A2(_1577_),
    .ZN(_0063_));
 CLKBUF_X3 _2299_ (.A(_1447_),
    .Z(_1578_));
 BUF_X2 _2300_ (.A(net56),
    .Z(_1579_));
 AND2_X1 _2301_ (.A1(_1571_),
    .A2(net55),
    .ZN(_1580_));
 NAND4_X2 _2302_ (.A1(_1561_),
    .A2(_1568_),
    .A3(_1562_),
    .A4(_1580_),
    .ZN(_1581_));
 OAI21_X1 _2303_ (.A(_1579_),
    .B1(_1547_),
    .B2(_1581_),
    .ZN(_1582_));
 OR3_X1 _2304_ (.A1(_1579_),
    .A2(_1547_),
    .A3(_1581_),
    .ZN(_1583_));
 AOI21_X1 _2305_ (.A(_1578_),
    .B1(_1582_),
    .B2(_1583_),
    .ZN(_0064_));
 BUF_X1 _2306_ (.A(net57),
    .Z(_1584_));
 AND4_X1 _2307_ (.A1(_1561_),
    .A2(_1568_),
    .A3(_1562_),
    .A4(_1580_),
    .ZN(_1585_));
 BUF_X4 _2308_ (.A(_1585_),
    .Z(_1586_));
 NAND4_X1 _2309_ (.A1(_1539_),
    .A2(_1579_),
    .A3(_1542_),
    .A4(_1586_),
    .ZN(_1587_));
 XOR2_X1 _2310_ (.A(_1584_),
    .B(_1587_),
    .Z(_1588_));
 NOR2_X1 _2311_ (.A1(_1560_),
    .A2(_1588_),
    .ZN(_0065_));
 NAND2_X1 _2312_ (.A1(_1579_),
    .A2(_1584_),
    .ZN(_1589_));
 NOR4_X1 _2313_ (.A1(_1536_),
    .A2(_1545_),
    .A3(_1581_),
    .A4(_1589_),
    .ZN(_1590_));
 XNOR2_X1 _2314_ (.A(net58),
    .B(_1590_),
    .ZN(_1591_));
 NOR2_X1 _2315_ (.A1(_1560_),
    .A2(_1591_),
    .ZN(_0066_));
 AND3_X1 _2316_ (.A1(_1579_),
    .A2(_1584_),
    .A3(net58),
    .ZN(_1592_));
 NAND4_X1 _2317_ (.A1(_1539_),
    .A2(_1542_),
    .A3(_1586_),
    .A4(_1592_),
    .ZN(_1593_));
 XOR2_X1 _2318_ (.A(net59),
    .B(_1593_),
    .Z(_1594_));
 NOR2_X1 _2319_ (.A1(_1560_),
    .A2(_1594_),
    .ZN(_0067_));
 AND4_X1 _2320_ (.A1(_1579_),
    .A2(_1584_),
    .A3(net58),
    .A4(net59),
    .ZN(_1595_));
 INV_X1 _2321_ (.A(_1595_),
    .ZN(_1596_));
 NOR4_X1 _2322_ (.A1(_1536_),
    .A2(_1545_),
    .A3(_1581_),
    .A4(_1596_),
    .ZN(_1597_));
 XNOR2_X1 _2323_ (.A(net60),
    .B(_1597_),
    .ZN(_1598_));
 NOR2_X1 _2324_ (.A1(_1560_),
    .A2(_1598_),
    .ZN(_0068_));
 AND2_X1 _2325_ (.A1(net60),
    .A2(_1595_),
    .ZN(_1599_));
 NAND4_X1 _2326_ (.A1(_1539_),
    .A2(_1542_),
    .A3(_1586_),
    .A4(_1599_),
    .ZN(_1600_));
 XOR2_X1 _2327_ (.A(net61),
    .B(_1600_),
    .Z(_1601_));
 NOR2_X1 _2328_ (.A1(_1560_),
    .A2(_1601_),
    .ZN(_0069_));
 BUF_X1 _2329_ (.A(net62),
    .Z(_1602_));
 AND3_X2 _2330_ (.A1(net60),
    .A2(net61),
    .A3(_1595_),
    .ZN(_1603_));
 NAND2_X1 _2331_ (.A1(_1586_),
    .A2(_1603_),
    .ZN(_1604_));
 OAI21_X1 _2332_ (.A(_1602_),
    .B1(_1547_),
    .B2(_1604_),
    .ZN(_1605_));
 OR3_X1 _2333_ (.A1(_1602_),
    .A2(_1547_),
    .A3(_1604_),
    .ZN(_1606_));
 AOI21_X1 _2334_ (.A(_1578_),
    .B1(_1605_),
    .B2(_1606_),
    .ZN(_0070_));
 BUF_X2 _2335_ (.A(net63),
    .Z(_1607_));
 NAND4_X1 _2336_ (.A1(_1517_),
    .A2(_1565_),
    .A3(_1417_),
    .A4(_1519_),
    .ZN(_1608_));
 XOR2_X1 _2337_ (.A(_1607_),
    .B(_1608_),
    .Z(_1609_));
 NOR2_X1 _2338_ (.A1(_1560_),
    .A2(_1609_),
    .ZN(_0071_));
 NAND4_X1 _2339_ (.A1(_1539_),
    .A2(_1542_),
    .A3(_1586_),
    .A4(_1603_),
    .ZN(_1610_));
 INV_X1 _2340_ (.A(_1602_),
    .ZN(_1611_));
 OAI21_X1 _2341_ (.A(net64),
    .B1(_1610_),
    .B2(_1611_),
    .ZN(_1612_));
 OR3_X1 _2342_ (.A1(_1611_),
    .A2(net64),
    .A3(_1610_),
    .ZN(_1613_));
 AOI21_X1 _2343_ (.A(_1578_),
    .B1(_1612_),
    .B2(_1613_),
    .ZN(_0072_));
 CLKBUF_X3 _2344_ (.A(_1559_),
    .Z(_1614_));
 INV_X1 _2345_ (.A(net65),
    .ZN(_1615_));
 AND4_X2 _2346_ (.A1(net46),
    .A2(_1602_),
    .A3(net64),
    .A4(_1540_),
    .ZN(_1616_));
 NAND4_X4 _2347_ (.A1(_1528_),
    .A2(_1586_),
    .A3(_1603_),
    .A4(_1616_),
    .ZN(_1617_));
 XNOR2_X1 _2348_ (.A(_1615_),
    .B(_1617_),
    .ZN(_1618_));
 NOR2_X1 _2349_ (.A1(_1614_),
    .A2(_1618_),
    .ZN(_0073_));
 BUF_X1 _2350_ (.A(net66),
    .Z(_1619_));
 NAND4_X4 _2351_ (.A1(_1525_),
    .A2(_1586_),
    .A3(_1603_),
    .A4(_1616_),
    .ZN(_1620_));
 OAI21_X1 _2352_ (.A(_1619_),
    .B1(_1620_),
    .B2(_1615_),
    .ZN(_1621_));
 OR3_X1 _2353_ (.A1(_1615_),
    .A2(_1619_),
    .A3(_1620_),
    .ZN(_1622_));
 AOI21_X1 _2354_ (.A(_1578_),
    .B1(_1621_),
    .B2(_1622_),
    .ZN(_0074_));
 NAND2_X1 _2355_ (.A1(net65),
    .A2(_1619_),
    .ZN(_1623_));
 OAI21_X1 _2356_ (.A(net67),
    .B1(_1617_),
    .B2(_1623_),
    .ZN(_1624_));
 OR3_X1 _2357_ (.A1(net67),
    .A2(_1617_),
    .A3(_1623_),
    .ZN(_1625_));
 AOI21_X1 _2358_ (.A(_1578_),
    .B1(_1624_),
    .B2(_1625_),
    .ZN(_0075_));
 NAND3_X1 _2359_ (.A1(net65),
    .A2(_1619_),
    .A3(net67),
    .ZN(_1626_));
 OAI21_X1 _2360_ (.A(net68),
    .B1(_1620_),
    .B2(_1626_),
    .ZN(_1627_));
 OR3_X1 _2361_ (.A1(net68),
    .A2(_1620_),
    .A3(_1626_),
    .ZN(_1628_));
 AOI21_X1 _2362_ (.A(_1578_),
    .B1(_1627_),
    .B2(_1628_),
    .ZN(_0076_));
 CLKBUF_X2 _2363_ (.A(net69),
    .Z(_1629_));
 INV_X1 _2364_ (.A(net68),
    .ZN(_1630_));
 OR2_X1 _2365_ (.A1(_1630_),
    .A2(_1626_),
    .ZN(_1631_));
 OAI21_X1 _2366_ (.A(_1629_),
    .B1(_1617_),
    .B2(_1631_),
    .ZN(_1632_));
 OR3_X1 _2367_ (.A1(_1629_),
    .A2(_1617_),
    .A3(_1631_),
    .ZN(_1633_));
 AOI21_X1 _2368_ (.A(_1578_),
    .B1(_1632_),
    .B2(_1633_),
    .ZN(_0077_));
 NOR2_X1 _2369_ (.A1(_1630_),
    .A2(_1626_),
    .ZN(_1634_));
 NAND2_X1 _2370_ (.A1(_1629_),
    .A2(_1634_),
    .ZN(_1635_));
 OAI21_X1 _2371_ (.A(net70),
    .B1(_1620_),
    .B2(_1635_),
    .ZN(_1636_));
 OR3_X1 _2372_ (.A1(net70),
    .A2(_1620_),
    .A3(_1635_),
    .ZN(_1637_));
 AOI21_X1 _2373_ (.A(_1578_),
    .B1(_1636_),
    .B2(_1637_),
    .ZN(_0078_));
 NAND3_X2 _2374_ (.A1(_1629_),
    .A2(net70),
    .A3(_1634_),
    .ZN(_1638_));
 OAI21_X1 _2375_ (.A(net71),
    .B1(_1617_),
    .B2(_1638_),
    .ZN(_1639_));
 OR3_X1 _2376_ (.A1(net71),
    .A2(_1617_),
    .A3(_1638_),
    .ZN(_1640_));
 AOI21_X1 _2377_ (.A(_1578_),
    .B1(_1639_),
    .B2(_1640_),
    .ZN(_0079_));
 INV_X1 _2378_ (.A(net72),
    .ZN(_1641_));
 NOR2_X1 _2379_ (.A1(_1641_),
    .A2(_1474_),
    .ZN(_1642_));
 NOR2_X1 _2380_ (.A1(net72),
    .A2(_1490_),
    .ZN(_1643_));
 INV_X1 _2381_ (.A(net71),
    .ZN(_1644_));
 NOR3_X1 _2382_ (.A1(_1644_),
    .A2(_1620_),
    .A3(_1638_),
    .ZN(_1645_));
 MUX2_X1 _2383_ (.A(_1642_),
    .B(_1643_),
    .S(_1645_),
    .Z(_0080_));
 AND2_X1 _2384_ (.A1(net73),
    .A2(_1346_),
    .ZN(_1646_));
 NOR2_X1 _2385_ (.A1(net73),
    .A2(_1490_),
    .ZN(_1647_));
 NOR4_X1 _2386_ (.A1(_1644_),
    .A2(_1641_),
    .A3(_1617_),
    .A4(_1638_),
    .ZN(_1648_));
 MUX2_X1 _2387_ (.A(_1646_),
    .B(_1647_),
    .S(_1648_),
    .Z(_0081_));
 AND3_X1 _2388_ (.A1(_1517_),
    .A2(_1565_),
    .A3(_1607_),
    .ZN(_1649_));
 NAND3_X1 _2389_ (.A1(_1470_),
    .A2(_1520_),
    .A3(_1649_),
    .ZN(_1650_));
 XOR2_X1 _2390_ (.A(net74),
    .B(_1650_),
    .Z(_1651_));
 NOR2_X1 _2391_ (.A1(_1614_),
    .A2(_1651_),
    .ZN(_0082_));
 INV_X1 _2392_ (.A(\prev_event_inc[5] ),
    .ZN(_1652_));
 NAND3_X1 _2393_ (.A1(_1511_),
    .A2(_1652_),
    .A3(net5),
    .ZN(_1653_));
 MUX2_X1 _2394_ (.A(_0008_),
    .B(net75),
    .S(_1653_),
    .Z(_1654_));
 AND2_X1 _2395_ (.A1(_1348_),
    .A2(_1654_),
    .ZN(_0083_));
 MUX2_X1 _2396_ (.A(_0009_),
    .B(net76),
    .S(_1653_),
    .Z(_1655_));
 AND2_X1 _2397_ (.A1(_1348_),
    .A2(_1655_),
    .ZN(_0084_));
 CLKBUF_X2 _2398_ (.A(net77),
    .Z(_1656_));
 AND2_X1 _2399_ (.A1(net5),
    .A2(_1928_),
    .ZN(_1657_));
 NAND3_X1 _2400_ (.A1(_1511_),
    .A2(_1652_),
    .A3(_1657_),
    .ZN(_1658_));
 XOR2_X1 _2401_ (.A(_1656_),
    .B(_1658_),
    .Z(_1659_));
 NOR2_X1 _2402_ (.A1(_1614_),
    .A2(_1659_),
    .ZN(_0085_));
 CLKBUF_X2 _2403_ (.A(net78),
    .Z(_1660_));
 INV_X1 _2404_ (.A(net5),
    .ZN(_1661_));
 NAND2_X1 _2405_ (.A1(net75),
    .A2(net76),
    .ZN(_1662_));
 NOR4_X4 _2406_ (.A1(_1369_),
    .A2(\prev_event_inc[5] ),
    .A3(_1661_),
    .A4(_1662_),
    .ZN(_1663_));
 NAND2_X1 _2407_ (.A1(_1656_),
    .A2(_1663_),
    .ZN(_1664_));
 XOR2_X1 _2408_ (.A(_1660_),
    .B(_1664_),
    .Z(_1665_));
 NOR2_X1 _2409_ (.A1(_1614_),
    .A2(_1665_),
    .ZN(_0086_));
 NAND2_X1 _2410_ (.A1(_1656_),
    .A2(_1660_),
    .ZN(_1666_));
 NOR2_X1 _2411_ (.A1(_1658_),
    .A2(_1666_),
    .ZN(_1667_));
 XNOR2_X1 _2412_ (.A(net79),
    .B(_1667_),
    .ZN(_1668_));
 NOR2_X1 _2413_ (.A1(_1614_),
    .A2(_1668_),
    .ZN(_0087_));
 NAND4_X1 _2414_ (.A1(_1656_),
    .A2(_1660_),
    .A3(net79),
    .A4(_1663_),
    .ZN(_0280_));
 XOR2_X1 _2415_ (.A(net80),
    .B(_0280_),
    .Z(_0281_));
 NOR2_X1 _2416_ (.A1(_1614_),
    .A2(_0281_),
    .ZN(_0088_));
 BUF_X2 _2417_ (.A(net81),
    .Z(_0282_));
 AND4_X1 _2418_ (.A1(_1656_),
    .A2(_1660_),
    .A3(net79),
    .A4(net80),
    .ZN(_0283_));
 BUF_X4 _2419_ (.A(_0283_),
    .Z(_0284_));
 AND4_X2 _2420_ (.A1(_1351_),
    .A2(_1652_),
    .A3(_1657_),
    .A4(_0284_),
    .ZN(_0285_));
 BUF_X4 _2421_ (.A(_0285_),
    .Z(_0286_));
 XNOR2_X1 _2422_ (.A(_0282_),
    .B(_0286_),
    .ZN(_0287_));
 NOR2_X1 _2423_ (.A1(_1614_),
    .A2(_0287_),
    .ZN(_0089_));
 CLKBUF_X2 _2424_ (.A(net82),
    .Z(_0288_));
 NAND3_X1 _2425_ (.A1(_0282_),
    .A2(_1663_),
    .A3(_0284_),
    .ZN(_0289_));
 XOR2_X1 _2426_ (.A(_0288_),
    .B(_0289_),
    .Z(_0290_));
 NOR2_X1 _2427_ (.A1(_1614_),
    .A2(_0290_),
    .ZN(_0090_));
 NAND3_X1 _2428_ (.A1(_0282_),
    .A2(_0288_),
    .A3(_0286_),
    .ZN(_0291_));
 XOR2_X1 _2429_ (.A(net83),
    .B(_0291_),
    .Z(_0292_));
 NOR2_X1 _2430_ (.A1(_1614_),
    .A2(_0292_),
    .ZN(_0091_));
 AND3_X1 _2431_ (.A1(_0282_),
    .A2(_0288_),
    .A3(net83),
    .ZN(_0293_));
 NAND3_X1 _2432_ (.A1(_1663_),
    .A2(_0284_),
    .A3(_0293_),
    .ZN(_0294_));
 XOR2_X1 _2433_ (.A(net84),
    .B(_0294_),
    .Z(_0295_));
 NOR2_X1 _2434_ (.A1(_1614_),
    .A2(_0295_),
    .ZN(_0092_));
 CLKBUF_X3 _2435_ (.A(_1559_),
    .Z(_0296_));
 BUF_X2 _2436_ (.A(net85),
    .Z(_0297_));
 AND4_X1 _2437_ (.A1(_1517_),
    .A2(_1565_),
    .A3(_1607_),
    .A4(net74),
    .ZN(_0298_));
 NAND3_X1 _2438_ (.A1(_1418_),
    .A2(_1520_),
    .A3(_0298_),
    .ZN(_0299_));
 XOR2_X1 _2439_ (.A(_0297_),
    .B(_0299_),
    .Z(_0300_));
 NOR2_X1 _2440_ (.A1(_0296_),
    .A2(_0300_),
    .ZN(_0093_));
 BUF_X1 _2441_ (.A(net86),
    .Z(_0301_));
 AND4_X1 _2442_ (.A1(_0282_),
    .A2(_0288_),
    .A3(net83),
    .A4(net84),
    .ZN(_0302_));
 NAND2_X1 _2443_ (.A1(_0286_),
    .A2(_0302_),
    .ZN(_0303_));
 XOR2_X1 _2444_ (.A(_0301_),
    .B(_0303_),
    .Z(_0304_));
 NOR2_X1 _2445_ (.A1(_0296_),
    .A2(_0304_),
    .ZN(_0094_));
 NAND4_X1 _2446_ (.A1(_0301_),
    .A2(_1663_),
    .A3(_0284_),
    .A4(_0302_),
    .ZN(_0305_));
 XOR2_X1 _2447_ (.A(net87),
    .B(_0305_),
    .Z(_0306_));
 NOR2_X1 _2448_ (.A1(_0296_),
    .A2(_0306_),
    .ZN(_0095_));
 BUF_X2 _2449_ (.A(net88),
    .Z(_0307_));
 AND3_X2 _2450_ (.A1(_0301_),
    .A2(net87),
    .A3(_0302_),
    .ZN(_0308_));
 BUF_X4 _2451_ (.A(_0308_),
    .Z(_0309_));
 NAND2_X1 _2452_ (.A1(_0286_),
    .A2(_0309_),
    .ZN(_0310_));
 XOR2_X1 _2453_ (.A(_0307_),
    .B(_0310_),
    .Z(_0311_));
 NOR2_X1 _2454_ (.A1(_0296_),
    .A2(_0311_),
    .ZN(_0096_));
 BUF_X2 _2455_ (.A(net89),
    .Z(_0312_));
 NAND4_X1 _2456_ (.A1(_0307_),
    .A2(_1663_),
    .A3(_0284_),
    .A4(_0308_),
    .ZN(_0313_));
 XOR2_X1 _2457_ (.A(_0312_),
    .B(_0313_),
    .Z(_0314_));
 NOR2_X1 _2458_ (.A1(_0296_),
    .A2(_0314_),
    .ZN(_0097_));
 NAND4_X1 _2459_ (.A1(_0307_),
    .A2(_0312_),
    .A3(_0285_),
    .A4(_0308_),
    .ZN(_0315_));
 XOR2_X1 _2460_ (.A(net90),
    .B(_0315_),
    .Z(_0316_));
 NOR2_X1 _2461_ (.A1(_0296_),
    .A2(_0316_),
    .ZN(_0098_));
 BUF_X2 _2462_ (.A(net91),
    .Z(_0317_));
 AND3_X1 _2463_ (.A1(_0307_),
    .A2(_0312_),
    .A3(net90),
    .ZN(_0318_));
 NAND4_X1 _2464_ (.A1(_1663_),
    .A2(_0284_),
    .A3(_0309_),
    .A4(_0318_),
    .ZN(_0319_));
 XOR2_X1 _2465_ (.A(_0317_),
    .B(_0319_),
    .Z(_0320_));
 NOR2_X1 _2466_ (.A1(_0296_),
    .A2(_0320_),
    .ZN(_0099_));
 INV_X2 _2467_ (.A(net92),
    .ZN(_0321_));
 NAND4_X1 _2468_ (.A1(_0317_),
    .A2(_0286_),
    .A3(_0309_),
    .A4(_0318_),
    .ZN(_0322_));
 XNOR2_X1 _2469_ (.A(_0321_),
    .B(_0322_),
    .ZN(_0323_));
 NOR2_X1 _2470_ (.A1(_0296_),
    .A2(_0323_),
    .ZN(_0100_));
 BUF_X2 _2471_ (.A(net93),
    .Z(_0324_));
 NAND4_X4 _2472_ (.A1(_0307_),
    .A2(_0312_),
    .A3(net90),
    .A4(_0317_),
    .ZN(_0325_));
 NOR2_X2 _2473_ (.A1(_0321_),
    .A2(_0325_),
    .ZN(_0326_));
 NAND4_X2 _2474_ (.A1(_1663_),
    .A2(_0284_),
    .A3(_0308_),
    .A4(_0326_),
    .ZN(_0327_));
 XOR2_X1 _2475_ (.A(_0324_),
    .B(_0327_),
    .Z(_0328_));
 NOR2_X1 _2476_ (.A1(_0296_),
    .A2(_0328_),
    .ZN(_0101_));
 BUF_X2 _2477_ (.A(net94),
    .Z(_0329_));
 NAND4_X1 _2478_ (.A1(_0324_),
    .A2(_0285_),
    .A3(_0309_),
    .A4(_0326_),
    .ZN(_0330_));
 XOR2_X1 _2479_ (.A(_0329_),
    .B(_0330_),
    .Z(_0331_));
 NOR2_X1 _2480_ (.A1(_0296_),
    .A2(_0331_),
    .ZN(_0102_));
 CLKBUF_X2 _2481_ (.A(net95),
    .Z(_0332_));
 NAND2_X1 _2482_ (.A1(_0324_),
    .A2(_0329_),
    .ZN(_0333_));
 OAI21_X1 _2483_ (.A(_0332_),
    .B1(_0327_),
    .B2(_0333_),
    .ZN(_0334_));
 OR3_X1 _2484_ (.A1(_0332_),
    .A2(_0327_),
    .A3(_0333_),
    .ZN(_0335_));
 AOI21_X1 _2485_ (.A(_1578_),
    .B1(_0334_),
    .B2(_0335_),
    .ZN(_0103_));
 BUF_X4 _2486_ (.A(_1559_),
    .Z(_0336_));
 NAND4_X1 _2487_ (.A1(_0297_),
    .A2(_1470_),
    .A3(_1519_),
    .A4(_0298_),
    .ZN(_0337_));
 XOR2_X1 _2488_ (.A(net96),
    .B(_0337_),
    .Z(_0338_));
 NOR2_X1 _2489_ (.A1(_0336_),
    .A2(_0338_),
    .ZN(_0104_));
 AND3_X1 _2490_ (.A1(_0324_),
    .A2(_0329_),
    .A3(_0332_),
    .ZN(_0339_));
 NAND4_X1 _2491_ (.A1(_0286_),
    .A2(_0309_),
    .A3(_0326_),
    .A4(_0339_),
    .ZN(_0340_));
 XOR2_X1 _2492_ (.A(net97),
    .B(_0340_),
    .Z(_0341_));
 NOR2_X1 _2493_ (.A1(_0336_),
    .A2(_0341_),
    .ZN(_0105_));
 BUF_X4 _2494_ (.A(_1447_),
    .Z(_0342_));
 BUF_X1 _2495_ (.A(net98),
    .Z(_0343_));
 NAND4_X4 _2496_ (.A1(_0324_),
    .A2(_0329_),
    .A3(_0332_),
    .A4(net97),
    .ZN(_0344_));
 OAI21_X1 _2497_ (.A(_0343_),
    .B1(_0327_),
    .B2(_0344_),
    .ZN(_0345_));
 OR3_X1 _2498_ (.A1(_0343_),
    .A2(_0327_),
    .A3(_0344_),
    .ZN(_0346_));
 AOI21_X1 _2499_ (.A(_0342_),
    .B1(_0345_),
    .B2(_0346_),
    .ZN(_0106_));
 INV_X1 _2500_ (.A(_0343_),
    .ZN(_0347_));
 NOR2_X1 _2501_ (.A1(_0347_),
    .A2(_0344_),
    .ZN(_0348_));
 NAND4_X1 _2502_ (.A1(_0286_),
    .A2(_0309_),
    .A3(_0326_),
    .A4(_0348_),
    .ZN(_0349_));
 XOR2_X1 _2503_ (.A(net99),
    .B(_0349_),
    .Z(_0350_));
 NOR2_X1 _2504_ (.A1(_0336_),
    .A2(_0350_),
    .ZN(_0107_));
 BUF_X2 _2505_ (.A(net100),
    .Z(_0351_));
 NAND2_X1 _2506_ (.A1(_0343_),
    .A2(net99),
    .ZN(_0352_));
 NOR4_X4 _2507_ (.A1(_0321_),
    .A2(_0325_),
    .A3(_0344_),
    .A4(_0352_),
    .ZN(_0353_));
 NAND4_X4 _2508_ (.A1(_1663_),
    .A2(_0284_),
    .A3(_0308_),
    .A4(_0353_),
    .ZN(_0354_));
 XOR2_X1 _2509_ (.A(_0351_),
    .B(_0354_),
    .Z(_0355_));
 NOR2_X1 _2510_ (.A1(_0336_),
    .A2(_0355_),
    .ZN(_0108_));
 CLKBUF_X2 _2511_ (.A(net101),
    .Z(_0356_));
 NAND4_X1 _2512_ (.A1(_0351_),
    .A2(_0285_),
    .A3(_0309_),
    .A4(_0353_),
    .ZN(_0357_));
 XOR2_X1 _2513_ (.A(_0356_),
    .B(_0357_),
    .Z(_0358_));
 NOR2_X1 _2514_ (.A1(_0336_),
    .A2(_0358_),
    .ZN(_0109_));
 CLKBUF_X2 _2515_ (.A(net102),
    .Z(_0359_));
 NAND2_X1 _2516_ (.A1(_0351_),
    .A2(_0356_),
    .ZN(_0360_));
 OAI21_X1 _2517_ (.A(_0359_),
    .B1(_0354_),
    .B2(_0360_),
    .ZN(_0361_));
 OR3_X1 _2518_ (.A1(_0359_),
    .A2(_0354_),
    .A3(_0360_),
    .ZN(_0362_));
 AOI21_X1 _2519_ (.A(_0342_),
    .B1(_0361_),
    .B2(_0362_),
    .ZN(_0110_));
 AND3_X1 _2520_ (.A1(_0351_),
    .A2(_0356_),
    .A3(_0359_),
    .ZN(_0363_));
 NAND4_X1 _2521_ (.A1(_0286_),
    .A2(_0309_),
    .A3(_0353_),
    .A4(_0363_),
    .ZN(_0364_));
 XOR2_X1 _2522_ (.A(net103),
    .B(_0364_),
    .Z(_0365_));
 NOR2_X1 _2523_ (.A1(_0336_),
    .A2(_0365_),
    .ZN(_0111_));
 BUF_X1 _2524_ (.A(net104),
    .Z(_0366_));
 NAND4_X2 _2525_ (.A1(_0351_),
    .A2(_0356_),
    .A3(_0359_),
    .A4(net103),
    .ZN(_0367_));
 OAI21_X1 _2526_ (.A(_0366_),
    .B1(_0354_),
    .B2(_0367_),
    .ZN(_0368_));
 OR3_X1 _2527_ (.A1(_0366_),
    .A2(_0354_),
    .A3(_0367_),
    .ZN(_0369_));
 AOI21_X1 _2528_ (.A(_0342_),
    .B1(_0368_),
    .B2(_0369_),
    .ZN(_0112_));
 BUF_X1 _2529_ (.A(net105),
    .Z(_0370_));
 INV_X1 _2530_ (.A(_0366_),
    .ZN(_0371_));
 NOR2_X1 _2531_ (.A1(_0371_),
    .A2(_0367_),
    .ZN(_0372_));
 NAND4_X1 _2532_ (.A1(_0286_),
    .A2(_0309_),
    .A3(_0353_),
    .A4(_0372_),
    .ZN(_0373_));
 XOR2_X1 _2533_ (.A(_0370_),
    .B(_0373_),
    .Z(_0374_));
 NOR2_X1 _2534_ (.A1(_0336_),
    .A2(_0374_),
    .ZN(_0113_));
 NAND2_X1 _2535_ (.A1(_0370_),
    .A2(_0372_),
    .ZN(_0375_));
 OAI21_X1 _2536_ (.A(net106),
    .B1(_0354_),
    .B2(_0375_),
    .ZN(_0376_));
 OR3_X1 _2537_ (.A1(net106),
    .A2(_0354_),
    .A3(_0375_),
    .ZN(_0377_));
 AOI21_X1 _2538_ (.A(_0342_),
    .B1(_0376_),
    .B2(_0377_),
    .ZN(_0114_));
 BUF_X2 _2539_ (.A(net107),
    .Z(_0378_));
 AND3_X1 _2540_ (.A1(_0297_),
    .A2(net96),
    .A3(_0298_),
    .ZN(_0379_));
 NAND3_X1 _2541_ (.A1(_1418_),
    .A2(_1520_),
    .A3(_0379_),
    .ZN(_0380_));
 XOR2_X1 _2542_ (.A(_0378_),
    .B(_0380_),
    .Z(_0381_));
 NOR2_X1 _2543_ (.A1(_0336_),
    .A2(_0381_),
    .ZN(_0115_));
 NAND3_X1 _2544_ (.A1(_0366_),
    .A2(_0370_),
    .A3(net106),
    .ZN(_0382_));
 NOR2_X1 _2545_ (.A1(_0367_),
    .A2(_0382_),
    .ZN(_0383_));
 NAND4_X1 _2546_ (.A1(_0286_),
    .A2(_0309_),
    .A3(_0353_),
    .A4(_0383_),
    .ZN(_0384_));
 XOR2_X1 _2547_ (.A(net108),
    .B(_0384_),
    .Z(_0385_));
 NOR2_X1 _2548_ (.A1(_0336_),
    .A2(_0385_),
    .ZN(_0116_));
 NAND2_X1 _2549_ (.A1(net108),
    .A2(_0383_),
    .ZN(_0386_));
 OAI21_X1 _2550_ (.A(net109),
    .B1(_0354_),
    .B2(_0386_),
    .ZN(_0387_));
 OR3_X1 _2551_ (.A1(net109),
    .A2(_0354_),
    .A3(_0386_),
    .ZN(_0388_));
 AOI21_X1 _2552_ (.A(_0342_),
    .B1(_0387_),
    .B2(_0388_),
    .ZN(_0117_));
 INV_X1 _2553_ (.A(net6),
    .ZN(_0389_));
 NOR3_X4 _2554_ (.A1(_1369_),
    .A2(\prev_event_inc[6] ),
    .A3(_0389_),
    .ZN(_0390_));
 MUX2_X1 _2555_ (.A(net110),
    .B(_0010_),
    .S(_0390_),
    .Z(_0391_));
 AND2_X1 _2556_ (.A1(_1348_),
    .A2(_0391_),
    .ZN(_0118_));
 MUX2_X1 _2557_ (.A(net111),
    .B(_0011_),
    .S(_0390_),
    .Z(_0392_));
 AND2_X1 _2558_ (.A1(_1348_),
    .A2(_0392_),
    .ZN(_0119_));
 BUF_X2 _2559_ (.A(net112),
    .Z(_0393_));
 BUF_X1 _2560_ (.A(_1929_),
    .Z(_0394_));
 CLKBUF_X3 _2561_ (.A(_0394_),
    .Z(_0395_));
 NAND2_X1 _2562_ (.A1(_0395_),
    .A2(_0390_),
    .ZN(_0396_));
 XOR2_X1 _2563_ (.A(_0393_),
    .B(_0396_),
    .Z(_0397_));
 NOR2_X1 _2564_ (.A1(_0336_),
    .A2(_0397_),
    .ZN(_0120_));
 CLKBUF_X3 _2565_ (.A(_1559_),
    .Z(_0398_));
 AND2_X1 _2566_ (.A1(net110),
    .A2(net111),
    .ZN(_0399_));
 CLKBUF_X3 _2567_ (.A(_0399_),
    .Z(_0400_));
 NAND3_X1 _2568_ (.A1(_0393_),
    .A2(_0390_),
    .A3(_0400_),
    .ZN(_0401_));
 XOR2_X1 _2569_ (.A(net113),
    .B(_0401_),
    .Z(_0402_));
 NOR2_X1 _2570_ (.A1(_0398_),
    .A2(_0402_),
    .ZN(_0121_));
 BUF_X1 _2571_ (.A(net114),
    .Z(_0403_));
 AND2_X1 _2572_ (.A1(_0393_),
    .A2(net113),
    .ZN(_0404_));
 NAND3_X1 _2573_ (.A1(_0395_),
    .A2(_0390_),
    .A3(_0404_),
    .ZN(_0405_));
 XOR2_X1 _2574_ (.A(_0403_),
    .B(_0405_),
    .Z(_0406_));
 NOR2_X1 _2575_ (.A1(_0398_),
    .A2(_0406_),
    .ZN(_0122_));
 NAND4_X1 _2576_ (.A1(_0403_),
    .A2(_0390_),
    .A3(_0399_),
    .A4(_0404_),
    .ZN(_0407_));
 XOR2_X1 _2577_ (.A(net115),
    .B(_0407_),
    .Z(_0408_));
 NOR2_X1 _2578_ (.A1(_0398_),
    .A2(_0408_),
    .ZN(_0123_));
 AND2_X1 _2579_ (.A1(_0403_),
    .A2(net115),
    .ZN(_0409_));
 NAND4_X1 _2580_ (.A1(_0395_),
    .A2(_0390_),
    .A3(_0404_),
    .A4(_0409_),
    .ZN(_0410_));
 XOR2_X1 _2581_ (.A(net116),
    .B(_0410_),
    .Z(_0411_));
 NOR2_X1 _2582_ (.A1(_0398_),
    .A2(_0411_),
    .ZN(_0124_));
 CLKBUF_X2 _2583_ (.A(net117),
    .Z(_0412_));
 NAND2_X1 _2584_ (.A1(net6),
    .A2(_0403_),
    .ZN(_0413_));
 NAND4_X2 _2585_ (.A1(_0393_),
    .A2(net113),
    .A3(net115),
    .A4(net116),
    .ZN(_0414_));
 NOR4_X4 _2586_ (.A1(_1369_),
    .A2(\prev_event_inc[6] ),
    .A3(_0413_),
    .A4(_0414_),
    .ZN(_0415_));
 CLKBUF_X3 _2587_ (.A(_0415_),
    .Z(_0416_));
 NAND2_X1 _2588_ (.A1(_0400_),
    .A2(_0416_),
    .ZN(_0417_));
 XOR2_X1 _2589_ (.A(_0412_),
    .B(_0417_),
    .Z(_0418_));
 NOR2_X1 _2590_ (.A1(_0398_),
    .A2(_0418_),
    .ZN(_0125_));
 NAND4_X1 _2591_ (.A1(_0378_),
    .A2(_1470_),
    .A3(_1519_),
    .A4(_0379_),
    .ZN(_0419_));
 XOR2_X1 _2592_ (.A(net118),
    .B(_0419_),
    .Z(_0420_));
 NOR2_X1 _2593_ (.A1(_0398_),
    .A2(_0420_),
    .ZN(_0126_));
 MUX2_X1 _2594_ (.A(_0015_),
    .B(net119),
    .S(_1352_),
    .Z(_0421_));
 AND2_X1 _2595_ (.A1(_1348_),
    .A2(_0421_),
    .ZN(_0127_));
 CLKBUF_X2 _2596_ (.A(net120),
    .Z(_0422_));
 NAND3_X1 _2597_ (.A1(_0412_),
    .A2(_0395_),
    .A3(_0416_),
    .ZN(_0423_));
 XOR2_X1 _2598_ (.A(_0422_),
    .B(_0423_),
    .Z(_0424_));
 NOR2_X1 _2599_ (.A1(_0398_),
    .A2(_0424_),
    .ZN(_0128_));
 BUF_X4 _2600_ (.A(_0415_),
    .Z(_0425_));
 NAND4_X1 _2601_ (.A1(_0412_),
    .A2(_0422_),
    .A3(_0399_),
    .A4(_0425_),
    .ZN(_0426_));
 XOR2_X1 _2602_ (.A(net121),
    .B(_0426_),
    .Z(_0427_));
 NOR2_X1 _2603_ (.A1(_0398_),
    .A2(_0427_),
    .ZN(_0129_));
 AND3_X1 _2604_ (.A1(_0412_),
    .A2(_0422_),
    .A3(net121),
    .ZN(_0428_));
 NAND3_X1 _2605_ (.A1(_0395_),
    .A2(_0416_),
    .A3(_0428_),
    .ZN(_0429_));
 XOR2_X1 _2606_ (.A(net122),
    .B(_0429_),
    .Z(_0430_));
 NOR2_X1 _2607_ (.A1(_0398_),
    .A2(_0430_),
    .ZN(_0130_));
 CLKBUF_X2 _2608_ (.A(net123),
    .Z(_0431_));
 AND4_X1 _2609_ (.A1(_0412_),
    .A2(_0422_),
    .A3(net121),
    .A4(net122),
    .ZN(_0432_));
 BUF_X4 _2610_ (.A(_0432_),
    .Z(_0433_));
 NAND3_X1 _2611_ (.A1(_0400_),
    .A2(_0416_),
    .A3(_0433_),
    .ZN(_0434_));
 XOR2_X1 _2612_ (.A(_0431_),
    .B(_0434_),
    .Z(_0435_));
 NOR2_X1 _2613_ (.A1(_0398_),
    .A2(_0435_),
    .ZN(_0131_));
 BUF_X4 _2614_ (.A(_1559_),
    .Z(_0436_));
 NAND4_X1 _2615_ (.A1(_0431_),
    .A2(_0394_),
    .A3(_0425_),
    .A4(_0433_),
    .ZN(_0437_));
 XOR2_X1 _2616_ (.A(net124),
    .B(_0437_),
    .Z(_0438_));
 NOR2_X1 _2617_ (.A1(_0436_),
    .A2(_0438_),
    .ZN(_0132_));
 AND2_X1 _2618_ (.A1(_0431_),
    .A2(net124),
    .ZN(_0439_));
 NAND4_X1 _2619_ (.A1(_0400_),
    .A2(_0416_),
    .A3(_0433_),
    .A4(_0439_),
    .ZN(_0440_));
 XOR2_X1 _2620_ (.A(net125),
    .B(_0440_),
    .Z(_0441_));
 NOR2_X1 _2621_ (.A1(_0436_),
    .A2(_0441_),
    .ZN(_0133_));
 AND2_X1 _2622_ (.A1(net125),
    .A2(_0394_),
    .ZN(_0442_));
 NAND4_X1 _2623_ (.A1(_0416_),
    .A2(_0433_),
    .A3(_0439_),
    .A4(_0442_),
    .ZN(_0443_));
 XOR2_X1 _2624_ (.A(net126),
    .B(_0443_),
    .Z(_0444_));
 NOR2_X1 _2625_ (.A1(_0436_),
    .A2(_0444_),
    .ZN(_0134_));
 AND4_X1 _2626_ (.A1(_0431_),
    .A2(net124),
    .A3(net125),
    .A4(net126),
    .ZN(_0445_));
 NAND4_X1 _2627_ (.A1(_0400_),
    .A2(_0416_),
    .A3(_0433_),
    .A4(_0445_),
    .ZN(_0446_));
 XOR2_X1 _2628_ (.A(net127),
    .B(_0446_),
    .Z(_0447_));
 NOR2_X1 _2629_ (.A1(_0436_),
    .A2(_0447_),
    .ZN(_0135_));
 AND2_X1 _2630_ (.A1(net127),
    .A2(_0445_),
    .ZN(_0448_));
 NAND4_X1 _2631_ (.A1(_0395_),
    .A2(_0416_),
    .A3(_0433_),
    .A4(_0448_),
    .ZN(_0449_));
 XOR2_X1 _2632_ (.A(net128),
    .B(_0449_),
    .Z(_0450_));
 NOR2_X1 _2633_ (.A1(_0436_),
    .A2(_0450_),
    .ZN(_0136_));
 AND2_X1 _2634_ (.A1(net127),
    .A2(net128),
    .ZN(_0451_));
 AND2_X1 _2635_ (.A1(_0445_),
    .A2(_0451_),
    .ZN(_0452_));
 NAND4_X1 _2636_ (.A1(_0400_),
    .A2(_0416_),
    .A3(_0433_),
    .A4(_0452_),
    .ZN(_0453_));
 XOR2_X1 _2637_ (.A(net129),
    .B(_0453_),
    .Z(_0454_));
 NOR2_X1 _2638_ (.A1(_0436_),
    .A2(_0454_),
    .ZN(_0137_));
 INV_X1 _2639_ (.A(net130),
    .ZN(_0455_));
 NAND4_X4 _2640_ (.A1(_1517_),
    .A2(_1565_),
    .A3(_1607_),
    .A4(net74),
    .ZN(_0456_));
 NAND4_X4 _2641_ (.A1(_0297_),
    .A2(net96),
    .A3(_0378_),
    .A4(net118),
    .ZN(_0457_));
 NOR2_X1 _2642_ (.A1(_0456_),
    .A2(_0457_),
    .ZN(_0458_));
 NAND3_X1 _2643_ (.A1(_1418_),
    .A2(_1520_),
    .A3(_0458_),
    .ZN(_0459_));
 XNOR2_X1 _2644_ (.A(_0455_),
    .B(_0459_),
    .ZN(_0460_));
 NOR2_X1 _2645_ (.A1(_0436_),
    .A2(_0460_),
    .ZN(_0138_));
 BUF_X2 _2646_ (.A(net131),
    .Z(_0461_));
 AND4_X1 _2647_ (.A1(net129),
    .A2(_0433_),
    .A3(_0445_),
    .A4(_0451_),
    .ZN(_0462_));
 BUF_X2 _2648_ (.A(_0462_),
    .Z(_0463_));
 NAND3_X2 _2649_ (.A1(_0394_),
    .A2(_0425_),
    .A3(_0463_),
    .ZN(_0464_));
 XOR2_X1 _2650_ (.A(_0461_),
    .B(_0464_),
    .Z(_0465_));
 NOR2_X1 _2651_ (.A1(_0436_),
    .A2(_0465_),
    .ZN(_0139_));
 BUF_X2 _2652_ (.A(net132),
    .Z(_0466_));
 NAND4_X1 _2653_ (.A1(_0461_),
    .A2(_0400_),
    .A3(_0425_),
    .A4(_0463_),
    .ZN(_0467_));
 XOR2_X1 _2654_ (.A(_0466_),
    .B(_0467_),
    .Z(_0468_));
 NOR2_X1 _2655_ (.A1(_0436_),
    .A2(_0468_),
    .ZN(_0140_));
 CLKBUF_X2 _2656_ (.A(net133),
    .Z(_0469_));
 AND2_X1 _2657_ (.A1(_0461_),
    .A2(_0466_),
    .ZN(_0470_));
 NAND4_X1 _2658_ (.A1(_0395_),
    .A2(_0416_),
    .A3(_0463_),
    .A4(_0470_),
    .ZN(_0471_));
 XOR2_X1 _2659_ (.A(_0469_),
    .B(_0471_),
    .Z(_0472_));
 NOR2_X1 _2660_ (.A1(_0436_),
    .A2(_0472_),
    .ZN(_0141_));
 CLKBUF_X3 _2661_ (.A(_1559_),
    .Z(_0473_));
 AND2_X1 _2662_ (.A1(_0469_),
    .A2(_0470_),
    .ZN(_0474_));
 NAND4_X1 _2663_ (.A1(_0400_),
    .A2(_0425_),
    .A3(_0463_),
    .A4(_0474_),
    .ZN(_0475_));
 XOR2_X1 _2664_ (.A(net134),
    .B(_0475_),
    .Z(_0476_));
 NOR2_X1 _2665_ (.A1(_0473_),
    .A2(_0476_),
    .ZN(_0142_));
 CLKBUF_X2 _2666_ (.A(net135),
    .Z(_0477_));
 NAND4_X2 _2667_ (.A1(_0461_),
    .A2(_0466_),
    .A3(_0469_),
    .A4(net134),
    .ZN(_0478_));
 OAI21_X1 _2668_ (.A(_0477_),
    .B1(_0464_),
    .B2(_0478_),
    .ZN(_0479_));
 OR3_X1 _2669_ (.A1(_0477_),
    .A2(_0464_),
    .A3(_0478_),
    .ZN(_0480_));
 AOI21_X1 _2670_ (.A(_0342_),
    .B1(_0479_),
    .B2(_0480_),
    .ZN(_0143_));
 CLKBUF_X2 _2671_ (.A(net136),
    .Z(_0481_));
 AND4_X1 _2672_ (.A1(_0461_),
    .A2(_0466_),
    .A3(_0469_),
    .A4(net134),
    .ZN(_0482_));
 AND2_X1 _2673_ (.A1(_0477_),
    .A2(_0482_),
    .ZN(_0483_));
 NAND4_X1 _2674_ (.A1(_0400_),
    .A2(_0425_),
    .A3(_0463_),
    .A4(_0483_),
    .ZN(_0484_));
 XOR2_X1 _2675_ (.A(_0481_),
    .B(_0484_),
    .Z(_0485_));
 NOR2_X1 _2676_ (.A1(_0473_),
    .A2(_0485_),
    .ZN(_0144_));
 CLKBUF_X2 _2677_ (.A(net137),
    .Z(_0486_));
 NAND2_X1 _2678_ (.A1(_0481_),
    .A2(_0483_),
    .ZN(_0487_));
 OAI21_X1 _2679_ (.A(_0486_),
    .B1(_0464_),
    .B2(_0487_),
    .ZN(_0488_));
 OR3_X1 _2680_ (.A1(_0486_),
    .A2(_0464_),
    .A3(_0487_),
    .ZN(_0489_));
 AOI21_X1 _2681_ (.A(_0342_),
    .B1(_0488_),
    .B2(_0489_),
    .ZN(_0145_));
 AND4_X1 _2682_ (.A1(_0477_),
    .A2(_0481_),
    .A3(_0486_),
    .A4(_0482_),
    .ZN(_0490_));
 NAND4_X1 _2683_ (.A1(_0400_),
    .A2(_0425_),
    .A3(_0463_),
    .A4(_0490_),
    .ZN(_0491_));
 XOR2_X1 _2684_ (.A(net138),
    .B(_0491_),
    .Z(_0492_));
 NOR2_X1 _2685_ (.A1(_0473_),
    .A2(_0492_),
    .ZN(_0146_));
 NAND4_X2 _2686_ (.A1(_0477_),
    .A2(_0481_),
    .A3(_0486_),
    .A4(net138),
    .ZN(_0493_));
 NOR2_X1 _2687_ (.A1(_0478_),
    .A2(_0493_),
    .ZN(_0494_));
 NAND4_X1 _2688_ (.A1(_0395_),
    .A2(_0425_),
    .A3(_0463_),
    .A4(_0494_),
    .ZN(_0495_));
 XOR2_X1 _2689_ (.A(net139),
    .B(_0495_),
    .Z(_0496_));
 NOR2_X1 _2690_ (.A1(_0473_),
    .A2(_0496_),
    .ZN(_0147_));
 CLKBUF_X2 _2691_ (.A(net140),
    .Z(_0497_));
 AND4_X1 _2692_ (.A1(net129),
    .A2(net139),
    .A3(_0399_),
    .A4(_0433_),
    .ZN(_0498_));
 NAND4_X2 _2693_ (.A1(_0415_),
    .A2(_0452_),
    .A3(_0494_),
    .A4(_0498_),
    .ZN(_0499_));
 XOR2_X1 _2694_ (.A(_0497_),
    .B(_0499_),
    .Z(_0500_));
 NOR2_X1 _2695_ (.A1(_0473_),
    .A2(_0500_),
    .ZN(_0148_));
 CLKBUF_X2 _2696_ (.A(net141),
    .Z(_0501_));
 NOR3_X1 _2697_ (.A1(_0455_),
    .A2(_0456_),
    .A3(_0457_),
    .ZN(_0502_));
 NAND3_X1 _2698_ (.A1(_1470_),
    .A2(_1520_),
    .A3(_0502_),
    .ZN(_0503_));
 XOR2_X1 _2699_ (.A(_0501_),
    .B(_0503_),
    .Z(_0504_));
 NOR2_X1 _2700_ (.A1(_0473_),
    .A2(_0504_),
    .ZN(_0149_));
 CLKBUF_X2 _2701_ (.A(net142),
    .Z(_0505_));
 NAND2_X1 _2702_ (.A1(net139),
    .A2(_0497_),
    .ZN(_0506_));
 NOR3_X1 _2703_ (.A1(_0478_),
    .A2(_0493_),
    .A3(_0506_),
    .ZN(_0507_));
 NAND4_X1 _2704_ (.A1(_0395_),
    .A2(_0425_),
    .A3(_0463_),
    .A4(_0507_),
    .ZN(_0508_));
 XOR2_X1 _2705_ (.A(_0505_),
    .B(_0508_),
    .Z(_0509_));
 NOR2_X1 _2706_ (.A1(_0473_),
    .A2(_0509_),
    .ZN(_0150_));
 BUF_X1 _2707_ (.A(net143),
    .Z(_0510_));
 NAND2_X1 _2708_ (.A1(_0497_),
    .A2(_0505_),
    .ZN(_0511_));
 OAI21_X1 _2709_ (.A(_0510_),
    .B1(_0499_),
    .B2(_0511_),
    .ZN(_0512_));
 OR3_X1 _2710_ (.A1(_0510_),
    .A2(_0499_),
    .A3(_0511_),
    .ZN(_0513_));
 AOI21_X1 _2711_ (.A(_0342_),
    .B1(_0512_),
    .B2(_0513_),
    .ZN(_0151_));
 NAND2_X1 _2712_ (.A1(_0505_),
    .A2(_0510_),
    .ZN(_0514_));
 NOR4_X1 _2713_ (.A1(_0478_),
    .A2(_0493_),
    .A3(_0506_),
    .A4(_0514_),
    .ZN(_0515_));
 NAND4_X1 _2714_ (.A1(_0395_),
    .A2(_0425_),
    .A3(_0463_),
    .A4(_0515_),
    .ZN(_0516_));
 XOR2_X1 _2715_ (.A(net144),
    .B(_0516_),
    .Z(_0517_));
 NOR2_X1 _2716_ (.A1(_0473_),
    .A2(_0517_),
    .ZN(_0152_));
 NAND4_X1 _2717_ (.A1(_0497_),
    .A2(_0505_),
    .A3(_0510_),
    .A4(net144),
    .ZN(_0518_));
 OAI21_X1 _2718_ (.A(net145),
    .B1(_0499_),
    .B2(_0518_),
    .ZN(_0519_));
 OR3_X1 _2719_ (.A1(net145),
    .A2(_0499_),
    .A3(_0518_),
    .ZN(_0520_));
 AOI21_X1 _2720_ (.A(_0342_),
    .B1(_0519_),
    .B2(_0520_),
    .ZN(_0153_));
 INV_X1 _2721_ (.A(net146),
    .ZN(_0521_));
 CLKBUF_X2 _2722_ (.A(event_inc[7]),
    .Z(_0522_));
 INV_X1 _2723_ (.A(_0522_),
    .ZN(_0523_));
 NOR3_X4 _2724_ (.A1(_1369_),
    .A2(\prev_event_inc[7] ),
    .A3(_0523_),
    .ZN(_0524_));
 NOR2_X1 _2725_ (.A1(_0521_),
    .A2(_0524_),
    .ZN(_0525_));
 AOI21_X1 _2726_ (.A(_0525_),
    .B1(_0524_),
    .B2(_0012_),
    .ZN(_0526_));
 NOR2_X1 _2727_ (.A1(_0473_),
    .A2(_0526_),
    .ZN(_0154_));
 MUX2_X1 _2728_ (.A(net147),
    .B(_0013_),
    .S(_0524_),
    .Z(_0527_));
 AND2_X1 _2729_ (.A1(_1348_),
    .A2(_0527_),
    .ZN(_0155_));
 INV_X1 _2730_ (.A(net148),
    .ZN(_0528_));
 NAND2_X1 _2731_ (.A1(_1930_),
    .A2(_0524_),
    .ZN(_0529_));
 XNOR2_X1 _2732_ (.A(_0528_),
    .B(_0529_),
    .ZN(_0530_));
 NOR2_X1 _2733_ (.A1(_0473_),
    .A2(_0530_),
    .ZN(_0156_));
 CLKBUF_X3 _2734_ (.A(_1559_),
    .Z(_0531_));
 INV_X1 _2735_ (.A(net149),
    .ZN(_0532_));
 NAND4_X1 _2736_ (.A1(net148),
    .A2(net147),
    .A3(net146),
    .A4(_0524_),
    .ZN(_0533_));
 XNOR2_X1 _2737_ (.A(_0532_),
    .B(_0533_),
    .ZN(_0534_));
 NOR2_X1 _2738_ (.A1(_0531_),
    .A2(_0534_),
    .ZN(_0157_));
 BUF_X2 _2739_ (.A(net150),
    .Z(_0535_));
 INV_X1 _2740_ (.A(\prev_event_inc[7] ),
    .ZN(_0536_));
 AND3_X1 _2741_ (.A1(_1930_),
    .A2(net148),
    .A3(net149),
    .ZN(_0537_));
 AND4_X1 _2742_ (.A1(_1350_),
    .A2(_0536_),
    .A3(_0522_),
    .A4(_0537_),
    .ZN(_0538_));
 BUF_X2 _2743_ (.A(_0538_),
    .Z(_0539_));
 XNOR2_X1 _2744_ (.A(_0535_),
    .B(_0539_),
    .ZN(_0540_));
 NOR2_X1 _2745_ (.A1(_0531_),
    .A2(_0540_),
    .ZN(_0158_));
 BUF_X2 _2746_ (.A(net151),
    .Z(_0541_));
 AND4_X1 _2747_ (.A1(net148),
    .A2(net147),
    .A3(net146),
    .A4(net149),
    .ZN(_0542_));
 NAND4_X1 _2748_ (.A1(_1511_),
    .A2(_0536_),
    .A3(_0522_),
    .A4(_0542_),
    .ZN(_0543_));
 INV_X1 _2749_ (.A(_0535_),
    .ZN(_0544_));
 OAI21_X1 _2750_ (.A(_0541_),
    .B1(_0543_),
    .B2(_0544_),
    .ZN(_0545_));
 INV_X1 _2751_ (.A(_0541_),
    .ZN(_0546_));
 AND4_X1 _2752_ (.A1(_1350_),
    .A2(_0536_),
    .A3(_0522_),
    .A4(_0542_),
    .ZN(_0547_));
 CLKBUF_X3 _2753_ (.A(_0547_),
    .Z(_0548_));
 NAND3_X1 _2754_ (.A1(_0535_),
    .A2(_0546_),
    .A3(_0548_),
    .ZN(_0549_));
 AOI21_X1 _2755_ (.A(_0342_),
    .B1(_0545_),
    .B2(_0549_),
    .ZN(_0159_));
 NAND4_X1 _2756_ (.A1(_0501_),
    .A2(_1417_),
    .A3(_1519_),
    .A4(_0502_),
    .ZN(_0550_));
 XOR2_X1 _2757_ (.A(net152),
    .B(_0550_),
    .Z(_0551_));
 NOR2_X1 _2758_ (.A1(_0531_),
    .A2(_0551_),
    .ZN(_0160_));
 INV_X1 _2759_ (.A(net153),
    .ZN(_0552_));
 NAND3_X1 _2760_ (.A1(_0535_),
    .A2(_0541_),
    .A3(_0539_),
    .ZN(_0553_));
 XNOR2_X1 _2761_ (.A(_0552_),
    .B(_0553_),
    .ZN(_0554_));
 NOR2_X1 _2762_ (.A1(_0531_),
    .A2(_0554_),
    .ZN(_0161_));
 INV_X1 _2763_ (.A(net154),
    .ZN(_0555_));
 NAND4_X1 _2764_ (.A1(_0535_),
    .A2(_0541_),
    .A3(net153),
    .A4(_0548_),
    .ZN(_0556_));
 XNOR2_X1 _2765_ (.A(_0555_),
    .B(_0556_),
    .ZN(_0557_));
 NOR2_X1 _2766_ (.A1(_0531_),
    .A2(_0557_),
    .ZN(_0162_));
 CLKBUF_X2 _2767_ (.A(net155),
    .Z(_0558_));
 NAND4_X4 _2768_ (.A1(_1351_),
    .A2(_0536_),
    .A3(_0522_),
    .A4(_0537_),
    .ZN(_0559_));
 NAND4_X4 _2769_ (.A1(_0535_),
    .A2(_0541_),
    .A3(net153),
    .A4(net154),
    .ZN(_0560_));
 NOR2_X1 _2770_ (.A1(_0559_),
    .A2(_0560_),
    .ZN(_0561_));
 XNOR2_X1 _2771_ (.A(_0558_),
    .B(_0561_),
    .ZN(_0562_));
 NOR2_X1 _2772_ (.A1(_0531_),
    .A2(_0562_),
    .ZN(_0163_));
 INV_X1 _2773_ (.A(net156),
    .ZN(_0563_));
 AND4_X1 _2774_ (.A1(_0535_),
    .A2(_0541_),
    .A3(net153),
    .A4(net154),
    .ZN(_0564_));
 NAND3_X1 _2775_ (.A1(_0558_),
    .A2(_0548_),
    .A3(_0564_),
    .ZN(_0565_));
 XNOR2_X1 _2776_ (.A(_0563_),
    .B(_0565_),
    .ZN(_0566_));
 NOR2_X1 _2777_ (.A1(_0531_),
    .A2(_0566_),
    .ZN(_0164_));
 BUF_X2 _2778_ (.A(net157),
    .Z(_0567_));
 NAND3_X2 _2779_ (.A1(_0558_),
    .A2(net156),
    .A3(_0564_),
    .ZN(_0568_));
 NOR2_X1 _2780_ (.A1(_0559_),
    .A2(_0568_),
    .ZN(_0569_));
 XNOR2_X1 _2781_ (.A(_0567_),
    .B(_0569_),
    .ZN(_0570_));
 NOR2_X1 _2782_ (.A1(_0531_),
    .A2(_0570_),
    .ZN(_0165_));
 BUF_X2 _2783_ (.A(net158),
    .Z(_0571_));
 INV_X1 _2784_ (.A(_0567_),
    .ZN(_0572_));
 NOR3_X1 _2785_ (.A1(_0572_),
    .A2(_0543_),
    .A3(_0568_),
    .ZN(_0573_));
 XNOR2_X1 _2786_ (.A(_0571_),
    .B(_0573_),
    .ZN(_0574_));
 NOR2_X1 _2787_ (.A1(_0531_),
    .A2(_0574_),
    .ZN(_0166_));
 INV_X2 _2788_ (.A(net159),
    .ZN(_0575_));
 NAND4_X2 _2789_ (.A1(_0558_),
    .A2(net156),
    .A3(_0567_),
    .A4(_0571_),
    .ZN(_0576_));
 NOR2_X1 _2790_ (.A1(_0560_),
    .A2(_0576_),
    .ZN(_0577_));
 NAND2_X1 _2791_ (.A1(_0539_),
    .A2(_0577_),
    .ZN(_0578_));
 XNOR2_X1 _2792_ (.A(_0575_),
    .B(_0578_),
    .ZN(_0579_));
 NOR2_X1 _2793_ (.A1(_0531_),
    .A2(_0579_),
    .ZN(_0167_));
 CLKBUF_X3 _2794_ (.A(_1559_),
    .Z(_0580_));
 INV_X2 _2795_ (.A(net160),
    .ZN(_0581_));
 NAND3_X1 _2796_ (.A1(net159),
    .A2(_0548_),
    .A3(_0577_),
    .ZN(_0582_));
 XNOR2_X1 _2797_ (.A(_0581_),
    .B(_0582_),
    .ZN(_0583_));
 NOR2_X1 _2798_ (.A1(_0580_),
    .A2(_0583_),
    .ZN(_0168_));
 INV_X1 _2799_ (.A(net161),
    .ZN(_0584_));
 NOR4_X4 _2800_ (.A1(_0575_),
    .A2(_0581_),
    .A3(_0560_),
    .A4(_0576_),
    .ZN(_0585_));
 NAND2_X1 _2801_ (.A1(_0539_),
    .A2(_0585_),
    .ZN(_0586_));
 XNOR2_X1 _2802_ (.A(_0584_),
    .B(_0586_),
    .ZN(_0587_));
 NOR2_X1 _2803_ (.A1(_0580_),
    .A2(_0587_),
    .ZN(_0169_));
 INV_X1 _2804_ (.A(net162),
    .ZN(_0588_));
 NAND3_X1 _2805_ (.A1(net161),
    .A2(_0548_),
    .A3(_0585_),
    .ZN(_0589_));
 XNOR2_X1 _2806_ (.A(_0588_),
    .B(_0589_),
    .ZN(_0590_));
 NOR2_X1 _2807_ (.A1(_0580_),
    .A2(_0590_),
    .ZN(_0170_));
 BUF_X1 _2808_ (.A(net163),
    .Z(_0591_));
 NAND3_X2 _2809_ (.A1(net130),
    .A2(_0501_),
    .A3(net152),
    .ZN(_0592_));
 NOR3_X4 _2810_ (.A1(_0456_),
    .A2(_0457_),
    .A3(_0592_),
    .ZN(_0593_));
 NAND3_X1 _2811_ (.A1(_1469_),
    .A2(_1519_),
    .A3(_0593_),
    .ZN(_0594_));
 XOR2_X1 _2812_ (.A(_0591_),
    .B(_0594_),
    .Z(_0595_));
 NOR2_X1 _2813_ (.A1(_0580_),
    .A2(_0595_),
    .ZN(_0171_));
 INV_X1 _2814_ (.A(net164),
    .ZN(_0596_));
 AND2_X1 _2815_ (.A1(net161),
    .A2(net162),
    .ZN(_0597_));
 NAND3_X1 _2816_ (.A1(_0539_),
    .A2(_0585_),
    .A3(_0597_),
    .ZN(_0598_));
 XNOR2_X1 _2817_ (.A(_0596_),
    .B(_0598_),
    .ZN(_0599_));
 NOR2_X1 _2818_ (.A1(_0580_),
    .A2(_0599_),
    .ZN(_0172_));
 INV_X1 _2819_ (.A(net165),
    .ZN(_0600_));
 NAND4_X1 _2820_ (.A1(net164),
    .A2(_0548_),
    .A3(_0585_),
    .A4(_0597_),
    .ZN(_0601_));
 XNOR2_X1 _2821_ (.A(_0600_),
    .B(_0601_),
    .ZN(_0602_));
 NOR2_X1 _2822_ (.A1(_0580_),
    .A2(_0602_),
    .ZN(_0173_));
 INV_X1 _2823_ (.A(net166),
    .ZN(_0603_));
 AND3_X1 _2824_ (.A1(net164),
    .A2(net165),
    .A3(_0597_),
    .ZN(_0604_));
 NAND3_X1 _2825_ (.A1(_0539_),
    .A2(_0585_),
    .A3(_0604_),
    .ZN(_0605_));
 XNOR2_X1 _2826_ (.A(_0603_),
    .B(_0605_),
    .ZN(_0606_));
 NOR2_X1 _2827_ (.A1(_0580_),
    .A2(_0606_),
    .ZN(_0174_));
 INV_X1 _2828_ (.A(net167),
    .ZN(_0607_));
 NAND4_X1 _2829_ (.A1(net166),
    .A2(_0548_),
    .A3(_0585_),
    .A4(_0604_),
    .ZN(_0608_));
 XNOR2_X1 _2830_ (.A(_0607_),
    .B(_0608_),
    .ZN(_0609_));
 NOR2_X1 _2831_ (.A1(_0580_),
    .A2(_0609_),
    .ZN(_0175_));
 BUF_X4 _2832_ (.A(net168),
    .Z(_0610_));
 INV_X1 _2833_ (.A(_0610_),
    .ZN(_0611_));
 NAND4_X2 _2834_ (.A1(net161),
    .A2(net162),
    .A3(net164),
    .A4(net165),
    .ZN(_0612_));
 NAND2_X1 _2835_ (.A1(net166),
    .A2(net167),
    .ZN(_0613_));
 NOR2_X1 _2836_ (.A1(_0612_),
    .A2(_0613_),
    .ZN(_0614_));
 NAND3_X1 _2837_ (.A1(_0539_),
    .A2(_0585_),
    .A3(_0614_),
    .ZN(_0615_));
 XNOR2_X1 _2838_ (.A(_0611_),
    .B(_0615_),
    .ZN(_0616_));
 NOR2_X1 _2839_ (.A1(_0580_),
    .A2(_0616_),
    .ZN(_0176_));
 INV_X1 _2840_ (.A(net169),
    .ZN(_0617_));
 NAND4_X1 _2841_ (.A1(_0610_),
    .A2(_0548_),
    .A3(_0585_),
    .A4(_0614_),
    .ZN(_0618_));
 XNOR2_X1 _2842_ (.A(_0617_),
    .B(_0618_),
    .ZN(_0619_));
 NOR2_X1 _2843_ (.A1(_0580_),
    .A2(_0619_),
    .ZN(_0177_));
 NAND2_X1 _2844_ (.A1(_0610_),
    .A2(net169),
    .ZN(_0620_));
 OAI21_X1 _2845_ (.A(net170),
    .B1(_0615_),
    .B2(_0620_),
    .ZN(_0621_));
 OR3_X1 _2846_ (.A1(net170),
    .A2(_0615_),
    .A3(_0620_),
    .ZN(_0622_));
 AOI21_X1 _2847_ (.A(_1356_),
    .B1(_0621_),
    .B2(_0622_),
    .ZN(_0178_));
 BUF_X4 _2848_ (.A(_1559_),
    .Z(_0623_));
 INV_X1 _2849_ (.A(net171),
    .ZN(_0624_));
 NAND3_X1 _2850_ (.A1(_0610_),
    .A2(net169),
    .A3(net170),
    .ZN(_0625_));
 NOR3_X2 _2851_ (.A1(_0612_),
    .A2(_0613_),
    .A3(_0625_),
    .ZN(_0626_));
 NAND3_X2 _2852_ (.A1(_0548_),
    .A2(_0585_),
    .A3(_0626_),
    .ZN(_0627_));
 XNOR2_X1 _2853_ (.A(_0624_),
    .B(_0627_),
    .ZN(_0628_));
 NOR2_X1 _2854_ (.A1(_0623_),
    .A2(_0628_),
    .ZN(_0179_));
 BUF_X1 _2855_ (.A(net172),
    .Z(_0629_));
 INV_X1 _2856_ (.A(net170),
    .ZN(_0630_));
 NAND4_X1 _2857_ (.A1(_0567_),
    .A2(_0571_),
    .A3(net159),
    .A4(net160),
    .ZN(_0631_));
 NAND4_X1 _2858_ (.A1(net166),
    .A2(net167),
    .A3(_0610_),
    .A4(net169),
    .ZN(_0632_));
 OR4_X2 _2859_ (.A1(_0630_),
    .A2(_0631_),
    .A3(_0612_),
    .A4(_0632_),
    .ZN(_0633_));
 NOR4_X1 _2860_ (.A1(_0624_),
    .A2(_0559_),
    .A3(_0568_),
    .A4(_0633_),
    .ZN(_0634_));
 XNOR2_X1 _2861_ (.A(_0629_),
    .B(_0634_),
    .ZN(_0635_));
 NOR2_X1 _2862_ (.A1(_0623_),
    .A2(_0635_),
    .ZN(_0180_));
 BUF_X1 _2863_ (.A(net173),
    .Z(_0636_));
 NAND2_X1 _2864_ (.A1(net171),
    .A2(_0629_),
    .ZN(_0637_));
 OAI21_X1 _2865_ (.A(_0636_),
    .B1(_0627_),
    .B2(_0637_),
    .ZN(_0638_));
 OR3_X1 _2866_ (.A1(_0636_),
    .A2(_0627_),
    .A3(_0637_),
    .ZN(_0639_));
 AOI21_X1 _2867_ (.A(_1356_),
    .B1(_0638_),
    .B2(_0639_),
    .ZN(_0181_));
 BUF_X1 _2868_ (.A(net174),
    .Z(_0640_));
 NAND4_X1 _2869_ (.A1(_0591_),
    .A2(_1417_),
    .A3(_1519_),
    .A4(_0593_),
    .ZN(_0641_));
 XOR2_X1 _2870_ (.A(_0640_),
    .B(_0641_),
    .Z(_0642_));
 NOR2_X1 _2871_ (.A1(_0623_),
    .A2(_0642_),
    .ZN(_0182_));
 NAND3_X1 _2872_ (.A1(net171),
    .A2(_0629_),
    .A3(_0636_),
    .ZN(_0643_));
 NOR4_X1 _2873_ (.A1(_0559_),
    .A2(_0568_),
    .A3(_0633_),
    .A4(_0643_),
    .ZN(_0644_));
 XNOR2_X1 _2874_ (.A(net175),
    .B(_0644_),
    .ZN(_0645_));
 NOR2_X1 _2875_ (.A1(_0623_),
    .A2(_0645_),
    .ZN(_0183_));
 INV_X1 _2876_ (.A(net176),
    .ZN(_0646_));
 AND4_X1 _2877_ (.A1(net171),
    .A2(_0629_),
    .A3(_0636_),
    .A4(net175),
    .ZN(_0647_));
 NAND4_X1 _2878_ (.A1(_0548_),
    .A2(_0585_),
    .A3(_0626_),
    .A4(_0647_),
    .ZN(_0648_));
 XNOR2_X1 _2879_ (.A(_0646_),
    .B(_0648_),
    .ZN(_0649_));
 NOR2_X1 _2880_ (.A1(_0623_),
    .A2(_0649_),
    .ZN(_0184_));
 BUF_X1 _2881_ (.A(net177),
    .Z(_0650_));
 NAND2_X1 _2882_ (.A1(net176),
    .A2(_0647_),
    .ZN(_0651_));
 NOR4_X1 _2883_ (.A1(_0559_),
    .A2(_0568_),
    .A3(_0633_),
    .A4(_0651_),
    .ZN(_0652_));
 XNOR2_X1 _2884_ (.A(_0650_),
    .B(_0652_),
    .ZN(_0653_));
 NOR2_X1 _2885_ (.A1(_0623_),
    .A2(_0653_),
    .ZN(_0185_));
 NAND3_X1 _2886_ (.A1(net176),
    .A2(_0650_),
    .A3(_0647_),
    .ZN(_0654_));
 OAI21_X1 _2887_ (.A(net178),
    .B1(_0627_),
    .B2(_0654_),
    .ZN(_0655_));
 OR3_X1 _2888_ (.A1(net178),
    .A2(_0627_),
    .A3(_0654_),
    .ZN(_0656_));
 AOI21_X1 _2889_ (.A(_1356_),
    .B1(_0655_),
    .B2(_0656_),
    .ZN(_0186_));
 NAND4_X1 _2890_ (.A1(net176),
    .A2(_0650_),
    .A3(net178),
    .A4(_0647_),
    .ZN(_0657_));
 NOR4_X1 _2891_ (.A1(_0559_),
    .A2(_0568_),
    .A3(_0633_),
    .A4(_0657_),
    .ZN(_0658_));
 XNOR2_X1 _2892_ (.A(net179),
    .B(_0658_),
    .ZN(_0659_));
 NOR2_X1 _2893_ (.A1(_0623_),
    .A2(_0659_),
    .ZN(_0187_));
 INV_X1 _2894_ (.A(net179),
    .ZN(_0660_));
 OR2_X1 _2895_ (.A1(_0660_),
    .A2(_0657_),
    .ZN(_0661_));
 OAI21_X1 _2896_ (.A(net180),
    .B1(_0627_),
    .B2(_0661_),
    .ZN(_0662_));
 OR3_X1 _2897_ (.A1(net180),
    .A2(_0627_),
    .A3(_0661_),
    .ZN(_0663_));
 AOI21_X1 _2898_ (.A(_1356_),
    .B1(_0662_),
    .B2(_0663_),
    .ZN(_0188_));
 BUF_X1 _2899_ (.A(net181),
    .Z(_0664_));
 AND2_X1 _2900_ (.A1(_0591_),
    .A2(_0640_),
    .ZN(_0665_));
 NAND4_X1 _2901_ (.A1(_1470_),
    .A2(_1520_),
    .A3(_0593_),
    .A4(_0665_),
    .ZN(_0666_));
 XOR2_X1 _2902_ (.A(_0664_),
    .B(_0666_),
    .Z(_0667_));
 NOR2_X1 _2903_ (.A1(_0623_),
    .A2(_0667_),
    .ZN(_0189_));
 AND2_X1 _2904_ (.A1(_0664_),
    .A2(_0665_),
    .ZN(_0668_));
 NAND4_X1 _2905_ (.A1(_1418_),
    .A2(_1520_),
    .A3(_0593_),
    .A4(_0668_),
    .ZN(_0669_));
 XOR2_X1 _2906_ (.A(net182),
    .B(_0669_),
    .Z(_0670_));
 NOR2_X1 _2907_ (.A1(_0623_),
    .A2(_0670_),
    .ZN(_0190_));
 AND4_X1 _2908_ (.A1(_0591_),
    .A2(_0640_),
    .A3(_0664_),
    .A4(net182),
    .ZN(_0671_));
 NAND4_X1 _2909_ (.A1(_1470_),
    .A2(_1519_),
    .A3(_0593_),
    .A4(_0671_),
    .ZN(_0672_));
 XOR2_X1 _2910_ (.A(net183),
    .B(_0672_),
    .Z(_0673_));
 NOR2_X1 _2911_ (.A1(_0623_),
    .A2(_0673_),
    .ZN(_0191_));
 CLKBUF_X3 _2912_ (.A(_1447_),
    .Z(_0674_));
 BUF_X1 _2913_ (.A(net184),
    .Z(_0675_));
 AND2_X1 _2914_ (.A1(net183),
    .A2(_0671_),
    .ZN(_0676_));
 NAND4_X1 _2915_ (.A1(_1418_),
    .A2(_1519_),
    .A3(_0593_),
    .A4(_0676_),
    .ZN(_0677_));
 XOR2_X1 _2916_ (.A(_0675_),
    .B(_0677_),
    .Z(_0678_));
 NOR2_X1 _2917_ (.A1(_0674_),
    .A2(_0678_),
    .ZN(_0192_));
 NAND2_X1 _2918_ (.A1(_0675_),
    .A2(_0676_),
    .ZN(_0679_));
 OAI21_X1 _2919_ (.A(net185),
    .B1(_0594_),
    .B2(_0679_),
    .ZN(_0680_));
 OR3_X1 _2920_ (.A1(net185),
    .A2(_0594_),
    .A3(_0679_),
    .ZN(_0681_));
 AOI21_X1 _2921_ (.A(_1356_),
    .B1(_0680_),
    .B2(_0681_),
    .ZN(_0193_));
 INV_X1 _2922_ (.A(net186),
    .ZN(_0682_));
 NAND4_X2 _2923_ (.A1(_1349_),
    .A2(net3),
    .A3(_1511_),
    .A4(_1931_),
    .ZN(_0683_));
 XNOR2_X1 _2924_ (.A(_0682_),
    .B(_0683_),
    .ZN(_0684_));
 NOR2_X1 _2925_ (.A1(_0674_),
    .A2(_0684_),
    .ZN(_0194_));
 INV_X1 _2926_ (.A(net187),
    .ZN(_0685_));
 NAND4_X1 _2927_ (.A1(_0591_),
    .A2(_0640_),
    .A3(_0664_),
    .A4(net182),
    .ZN(_0686_));
 NAND3_X1 _2928_ (.A1(net183),
    .A2(_0675_),
    .A3(net185),
    .ZN(_0687_));
 NOR2_X1 _2929_ (.A1(_0686_),
    .A2(_0687_),
    .ZN(_0688_));
 NAND4_X1 _2930_ (.A1(_1418_),
    .A2(_1520_),
    .A3(_0593_),
    .A4(_0688_),
    .ZN(_0689_));
 XNOR2_X1 _2931_ (.A(_0685_),
    .B(_0689_),
    .ZN(_0690_));
 NOR2_X1 _2932_ (.A1(_0674_),
    .A2(_0690_),
    .ZN(_0195_));
 NOR3_X1 _2933_ (.A1(_0685_),
    .A2(_0686_),
    .A3(_0687_),
    .ZN(_0691_));
 NAND4_X1 _2934_ (.A1(_1470_),
    .A2(_1519_),
    .A3(_0593_),
    .A4(_0691_),
    .ZN(_0692_));
 XOR2_X1 _2935_ (.A(net188),
    .B(_0692_),
    .Z(_0693_));
 NOR2_X1 _2936_ (.A1(_0674_),
    .A2(_0693_),
    .ZN(_0196_));
 INV_X2 _2937_ (.A(\prev_event_inc[1] ),
    .ZN(_0694_));
 NAND3_X1 _2938_ (.A1(_1511_),
    .A2(_0694_),
    .A3(net4),
    .ZN(_0695_));
 MUX2_X1 _2939_ (.A(_0000_),
    .B(net189),
    .S(_0695_),
    .Z(_0696_));
 AND2_X1 _2940_ (.A1(_1348_),
    .A2(_0696_),
    .ZN(_0197_));
 MUX2_X1 _2941_ (.A(_0001_),
    .B(net190),
    .S(_0695_),
    .Z(_0697_));
 AND2_X1 _2942_ (.A1(_1347_),
    .A2(_0697_),
    .ZN(_0198_));
 NAND4_X1 _2943_ (.A1(_1511_),
    .A2(_0694_),
    .A3(net4),
    .A4(_1925_),
    .ZN(_0698_));
 XOR2_X1 _2944_ (.A(net191),
    .B(_0698_),
    .Z(_0699_));
 NOR2_X1 _2945_ (.A1(_0674_),
    .A2(_0699_),
    .ZN(_0199_));
 BUF_X2 _2946_ (.A(net192),
    .Z(_0700_));
 INV_X1 _2947_ (.A(_0700_),
    .ZN(_0701_));
 AND2_X2 _2948_ (.A1(net4),
    .A2(net191),
    .ZN(_0702_));
 AND2_X1 _2949_ (.A1(net189),
    .A2(net190),
    .ZN(_0703_));
 NAND4_X4 _2950_ (.A1(_1350_),
    .A2(_0694_),
    .A3(_0702_),
    .A4(_0703_),
    .ZN(_0704_));
 CLKBUF_X3 _2951_ (.A(_0704_),
    .Z(_0705_));
 XNOR2_X1 _2952_ (.A(_0701_),
    .B(_0705_),
    .ZN(_0706_));
 NOR2_X1 _2953_ (.A1(_0674_),
    .A2(_0706_),
    .ZN(_0200_));
 BUF_X4 _2954_ (.A(net193),
    .Z(_0707_));
 NAND4_X4 _2955_ (.A1(_1351_),
    .A2(_0694_),
    .A3(_1925_),
    .A4(_0702_),
    .ZN(_0708_));
 CLKBUF_X3 _2956_ (.A(_0708_),
    .Z(_0709_));
 NOR2_X1 _2957_ (.A1(_0701_),
    .A2(_0709_),
    .ZN(_0710_));
 XNOR2_X1 _2958_ (.A(_0707_),
    .B(_0710_),
    .ZN(_0711_));
 NOR2_X1 _2959_ (.A1(_0674_),
    .A2(_0711_),
    .ZN(_0201_));
 BUF_X4 _2960_ (.A(net194),
    .Z(_0712_));
 NAND2_X1 _2961_ (.A1(_0700_),
    .A2(_0707_),
    .ZN(_0713_));
 NOR2_X1 _2962_ (.A1(_0705_),
    .A2(_0713_),
    .ZN(_0714_));
 XNOR2_X1 _2963_ (.A(_0712_),
    .B(_0714_),
    .ZN(_0715_));
 NOR2_X1 _2964_ (.A1(_0674_),
    .A2(_0715_),
    .ZN(_0202_));
 BUF_X4 _2965_ (.A(net195),
    .Z(_0716_));
 INV_X1 _2966_ (.A(_0712_),
    .ZN(_0717_));
 NOR3_X1 _2967_ (.A1(_0717_),
    .A2(_0709_),
    .A3(_0713_),
    .ZN(_0718_));
 XNOR2_X1 _2968_ (.A(_0716_),
    .B(_0718_),
    .ZN(_0719_));
 NOR2_X1 _2969_ (.A1(_0674_),
    .A2(_0719_),
    .ZN(_0203_));
 BUF_X2 _2970_ (.A(net196),
    .Z(_0720_));
 NAND4_X4 _2971_ (.A1(_0700_),
    .A2(_0707_),
    .A3(_0712_),
    .A4(_0716_),
    .ZN(_0721_));
 NOR2_X1 _2972_ (.A1(_0705_),
    .A2(_0721_),
    .ZN(_0722_));
 XNOR2_X1 _2973_ (.A(_0720_),
    .B(_0722_),
    .ZN(_0723_));
 NOR2_X1 _2974_ (.A1(_0674_),
    .A2(_0723_),
    .ZN(_0204_));
 CLKBUF_X3 _2975_ (.A(_1447_),
    .Z(_0724_));
 NOR3_X1 _2976_ (.A1(_0682_),
    .A2(_1352_),
    .A3(_1468_),
    .ZN(_0725_));
 XNOR2_X1 _2977_ (.A(_1414_),
    .B(_0725_),
    .ZN(_0726_));
 NOR2_X1 _2978_ (.A1(_0724_),
    .A2(_0726_),
    .ZN(_0205_));
 BUF_X2 _2979_ (.A(net198),
    .Z(_0727_));
 INV_X1 _2980_ (.A(_0720_),
    .ZN(_0728_));
 NOR3_X1 _2981_ (.A1(_0728_),
    .A2(_0709_),
    .A3(_0721_),
    .ZN(_0729_));
 XNOR2_X1 _2982_ (.A(_0727_),
    .B(_0729_),
    .ZN(_0730_));
 NOR2_X1 _2983_ (.A1(_0724_),
    .A2(_0730_),
    .ZN(_0206_));
 BUF_X4 _2984_ (.A(net199),
    .Z(_0731_));
 NAND2_X1 _2985_ (.A1(_0720_),
    .A2(_0727_),
    .ZN(_0732_));
 NOR3_X1 _2986_ (.A1(_0705_),
    .A2(_0721_),
    .A3(_0732_),
    .ZN(_0733_));
 XNOR2_X1 _2987_ (.A(_0731_),
    .B(_0733_),
    .ZN(_0734_));
 NOR2_X1 _2988_ (.A1(_0724_),
    .A2(_0734_),
    .ZN(_0207_));
 INV_X1 _2989_ (.A(_0731_),
    .ZN(_0735_));
 NOR4_X1 _2990_ (.A1(_0735_),
    .A2(_0708_),
    .A3(_0721_),
    .A4(_0732_),
    .ZN(_0736_));
 XNOR2_X1 _2991_ (.A(net200),
    .B(_0736_),
    .ZN(_0737_));
 NOR2_X1 _2992_ (.A1(_0724_),
    .A2(_0737_),
    .ZN(_0208_));
 NAND4_X2 _2993_ (.A1(_0720_),
    .A2(_0727_),
    .A3(_0731_),
    .A4(net200),
    .ZN(_0738_));
 NOR3_X1 _2994_ (.A1(_0705_),
    .A2(_0721_),
    .A3(_0738_),
    .ZN(_0739_));
 XNOR2_X1 _2995_ (.A(net201),
    .B(_0739_),
    .ZN(_0740_));
 NOR2_X1 _2996_ (.A1(_0724_),
    .A2(_0740_),
    .ZN(_0209_));
 BUF_X1 _2997_ (.A(net202),
    .Z(_0741_));
 INV_X1 _2998_ (.A(net201),
    .ZN(_0742_));
 OR2_X1 _2999_ (.A1(_0742_),
    .A2(_0738_),
    .ZN(_0743_));
 NOR3_X1 _3000_ (.A1(_0709_),
    .A2(_0721_),
    .A3(_0743_),
    .ZN(_0744_));
 XNOR2_X1 _3001_ (.A(_0741_),
    .B(_0744_),
    .ZN(_0745_));
 NOR2_X1 _3002_ (.A1(_0724_),
    .A2(_0745_),
    .ZN(_0210_));
 INV_X1 _3003_ (.A(_0741_),
    .ZN(_0746_));
 NOR4_X1 _3004_ (.A1(_0746_),
    .A2(_0704_),
    .A3(_0721_),
    .A4(_0743_),
    .ZN(_0747_));
 XNOR2_X1 _3005_ (.A(net203),
    .B(_0747_),
    .ZN(_0748_));
 NOR2_X1 _3006_ (.A1(_0724_),
    .A2(_0748_),
    .ZN(_0211_));
 BUF_X2 _3007_ (.A(net204),
    .Z(_0749_));
 NAND2_X1 _3008_ (.A1(_0741_),
    .A2(net203),
    .ZN(_0750_));
 OR4_X2 _3009_ (.A1(_0742_),
    .A2(_0721_),
    .A3(_0738_),
    .A4(_0750_),
    .ZN(_0751_));
 BUF_X8 _3010_ (.A(_0751_),
    .Z(_0752_));
 BUF_X8 _3011_ (.A(_0752_),
    .Z(_0753_));
 NOR2_X1 _3012_ (.A1(_0709_),
    .A2(_0753_),
    .ZN(_0754_));
 XNOR2_X1 _3013_ (.A(_0749_),
    .B(_0754_),
    .ZN(_0755_));
 NOR2_X1 _3014_ (.A1(_0724_),
    .A2(_0755_),
    .ZN(_0212_));
 INV_X1 _3015_ (.A(_0749_),
    .ZN(_0756_));
 NOR3_X1 _3016_ (.A1(_0756_),
    .A2(_0705_),
    .A3(_0753_),
    .ZN(_0757_));
 XNOR2_X1 _3017_ (.A(net205),
    .B(_0757_),
    .ZN(_0758_));
 NOR2_X1 _3018_ (.A1(_0724_),
    .A2(_0758_),
    .ZN(_0213_));
 NAND2_X1 _3019_ (.A1(_0749_),
    .A2(net205),
    .ZN(_0759_));
 NOR3_X1 _3020_ (.A1(_0709_),
    .A2(_0753_),
    .A3(_0759_),
    .ZN(_0760_));
 XNOR2_X1 _3021_ (.A(net206),
    .B(_0760_),
    .ZN(_0761_));
 NOR2_X1 _3022_ (.A1(_0724_),
    .A2(_0761_),
    .ZN(_0214_));
 CLKBUF_X3 _3023_ (.A(_1447_),
    .Z(_0762_));
 INV_X1 _3024_ (.A(net206),
    .ZN(_0763_));
 NOR4_X1 _3025_ (.A1(_0763_),
    .A2(_0704_),
    .A3(_0752_),
    .A4(_0759_),
    .ZN(_0764_));
 XNOR2_X1 _3026_ (.A(net207),
    .B(_0764_),
    .ZN(_0765_));
 NOR2_X1 _3027_ (.A1(_0762_),
    .A2(_0765_),
    .ZN(_0215_));
 NAND2_X1 _3028_ (.A1(net186),
    .A2(_1414_),
    .ZN(_0766_));
 NOR2_X1 _3029_ (.A1(_0683_),
    .A2(_0766_),
    .ZN(_0767_));
 XNOR2_X1 _3030_ (.A(_1415_),
    .B(_0767_),
    .ZN(_0768_));
 NOR2_X1 _3031_ (.A1(_0762_),
    .A2(_0768_),
    .ZN(_0216_));
 BUF_X2 _3032_ (.A(net209),
    .Z(_0769_));
 AND4_X2 _3033_ (.A1(_0749_),
    .A2(net205),
    .A3(net206),
    .A4(net207),
    .ZN(_0770_));
 INV_X1 _3034_ (.A(_0770_),
    .ZN(_0771_));
 NOR3_X1 _3035_ (.A1(_0709_),
    .A2(_0753_),
    .A3(_0771_),
    .ZN(_0772_));
 XNOR2_X1 _3036_ (.A(_0769_),
    .B(_0772_),
    .ZN(_0773_));
 NOR2_X1 _3037_ (.A1(_0762_),
    .A2(_0773_),
    .ZN(_0217_));
 BUF_X2 _3038_ (.A(net210),
    .Z(_0774_));
 NAND2_X1 _3039_ (.A1(_0769_),
    .A2(_0770_),
    .ZN(_0775_));
 NOR3_X1 _3040_ (.A1(_0705_),
    .A2(_0753_),
    .A3(_0775_),
    .ZN(_0776_));
 XNOR2_X1 _3041_ (.A(_0774_),
    .B(_0776_),
    .ZN(_0777_));
 NOR2_X1 _3042_ (.A1(_0762_),
    .A2(_0777_),
    .ZN(_0218_));
 CLKBUF_X2 _3043_ (.A(net211),
    .Z(_0778_));
 INV_X1 _3044_ (.A(_0774_),
    .ZN(_0779_));
 NOR4_X1 _3045_ (.A1(_0779_),
    .A2(_0708_),
    .A3(_0752_),
    .A4(_0775_),
    .ZN(_0780_));
 XNOR2_X1 _3046_ (.A(_0778_),
    .B(_0780_),
    .ZN(_0781_));
 NOR2_X1 _3047_ (.A1(_0762_),
    .A2(_0781_),
    .ZN(_0219_));
 NAND2_X1 _3048_ (.A1(_0774_),
    .A2(_0778_),
    .ZN(_0782_));
 NOR4_X1 _3049_ (.A1(_0705_),
    .A2(_0753_),
    .A3(_0775_),
    .A4(_0782_),
    .ZN(_0783_));
 XNOR2_X1 _3050_ (.A(net212),
    .B(_0783_),
    .ZN(_0784_));
 NOR2_X1 _3051_ (.A1(_0762_),
    .A2(_0784_),
    .ZN(_0220_));
 NAND3_X1 _3052_ (.A1(_0774_),
    .A2(_0778_),
    .A3(net212),
    .ZN(_0785_));
 NOR4_X1 _3053_ (.A1(_0709_),
    .A2(_0753_),
    .A3(_0775_),
    .A4(_0785_),
    .ZN(_0786_));
 XNOR2_X1 _3054_ (.A(net213),
    .B(_0786_),
    .ZN(_0787_));
 NOR2_X1 _3055_ (.A1(_0762_),
    .A2(_0787_),
    .ZN(_0221_));
 CLKBUF_X2 _3056_ (.A(net214),
    .Z(_0788_));
 AND4_X1 _3057_ (.A1(_0774_),
    .A2(_0778_),
    .A3(net212),
    .A4(net213),
    .ZN(_0789_));
 NAND3_X4 _3058_ (.A1(_0769_),
    .A2(_0770_),
    .A3(_0789_),
    .ZN(_0790_));
 NOR3_X1 _3059_ (.A1(_0705_),
    .A2(_0753_),
    .A3(_0790_),
    .ZN(_0791_));
 XNOR2_X1 _3060_ (.A(_0788_),
    .B(_0791_),
    .ZN(_0792_));
 NOR2_X1 _3061_ (.A1(_0762_),
    .A2(_0792_),
    .ZN(_0222_));
 CLKBUF_X2 _3062_ (.A(net215),
    .Z(_0793_));
 INV_X1 _3063_ (.A(_0788_),
    .ZN(_0794_));
 NOR4_X1 _3064_ (.A1(_0794_),
    .A2(_0708_),
    .A3(_0752_),
    .A4(_0790_),
    .ZN(_0795_));
 XNOR2_X1 _3065_ (.A(_0793_),
    .B(_0795_),
    .ZN(_0796_));
 NOR2_X1 _3066_ (.A1(_0762_),
    .A2(_0796_),
    .ZN(_0223_));
 BUF_X1 _3067_ (.A(net216),
    .Z(_0797_));
 NAND2_X1 _3068_ (.A1(_0788_),
    .A2(_0793_),
    .ZN(_0798_));
 NOR4_X1 _3069_ (.A1(_0705_),
    .A2(_0753_),
    .A3(_0790_),
    .A4(_0798_),
    .ZN(_0799_));
 XNOR2_X1 _3070_ (.A(_0797_),
    .B(_0799_),
    .ZN(_0800_));
 NOR2_X1 _3071_ (.A1(_0762_),
    .A2(_0800_),
    .ZN(_0224_));
 BUF_X4 _3072_ (.A(_1447_),
    .Z(_0801_));
 NAND3_X1 _3073_ (.A1(_0788_),
    .A2(_0793_),
    .A3(_0797_),
    .ZN(_0802_));
 NOR4_X1 _3074_ (.A1(_0709_),
    .A2(_0753_),
    .A3(_0790_),
    .A4(_0802_),
    .ZN(_0803_));
 XNOR2_X1 _3075_ (.A(net217),
    .B(_0803_),
    .ZN(_0804_));
 NOR2_X1 _3076_ (.A1(_0801_),
    .A2(_0804_),
    .ZN(_0225_));
 CLKBUF_X2 _3077_ (.A(net218),
    .Z(_0805_));
 AND4_X1 _3078_ (.A1(_0788_),
    .A2(_0793_),
    .A3(_0797_),
    .A4(net217),
    .ZN(_0806_));
 INV_X1 _3079_ (.A(_0806_),
    .ZN(_0807_));
 NOR4_X1 _3080_ (.A1(_0704_),
    .A2(_0752_),
    .A3(_0790_),
    .A4(_0807_),
    .ZN(_0808_));
 XNOR2_X1 _3081_ (.A(_0805_),
    .B(_0808_),
    .ZN(_0809_));
 NOR2_X1 _3082_ (.A1(_0801_),
    .A2(_0809_),
    .ZN(_0226_));
 INV_X1 _3083_ (.A(_1415_),
    .ZN(_0810_));
 NOR4_X1 _3084_ (.A1(_0810_),
    .A2(_1352_),
    .A3(_0766_),
    .A4(_1468_),
    .ZN(_0811_));
 XNOR2_X1 _3085_ (.A(net219),
    .B(_0811_),
    .ZN(_0812_));
 NOR2_X1 _3086_ (.A1(_0801_),
    .A2(_0812_),
    .ZN(_0227_));
 NAND2_X1 _3087_ (.A1(_0805_),
    .A2(_0806_),
    .ZN(_0813_));
 NOR4_X1 _3088_ (.A1(_0709_),
    .A2(_0752_),
    .A3(_0790_),
    .A4(_0813_),
    .ZN(_0814_));
 XNOR2_X1 _3089_ (.A(net220),
    .B(_0814_),
    .ZN(_0815_));
 NOR2_X1 _3090_ (.A1(_0801_),
    .A2(_0815_),
    .ZN(_0228_));
 NAND3_X1 _3091_ (.A1(_0805_),
    .A2(net220),
    .A3(_0806_),
    .ZN(_0816_));
 NOR4_X1 _3092_ (.A1(_0704_),
    .A2(_0752_),
    .A3(_0790_),
    .A4(_0816_),
    .ZN(_0817_));
 XNOR2_X1 _3093_ (.A(net221),
    .B(_0817_),
    .ZN(_0818_));
 NOR2_X1 _3094_ (.A1(_0801_),
    .A2(_0818_),
    .ZN(_0229_));
 AND3_X1 _3095_ (.A1(_0805_),
    .A2(net220),
    .A3(net221),
    .ZN(_0819_));
 NAND2_X1 _3096_ (.A1(_0806_),
    .A2(_0819_),
    .ZN(_0820_));
 NOR4_X1 _3097_ (.A1(_0708_),
    .A2(_0752_),
    .A3(_0790_),
    .A4(_0820_),
    .ZN(_0821_));
 XNOR2_X1 _3098_ (.A(net222),
    .B(_0821_),
    .ZN(_0822_));
 NOR2_X1 _3099_ (.A1(_0801_),
    .A2(_0822_),
    .ZN(_0230_));
 NAND3_X1 _3100_ (.A1(net222),
    .A2(_0806_),
    .A3(_0819_),
    .ZN(_0823_));
 NOR4_X1 _3101_ (.A1(_0704_),
    .A2(_0752_),
    .A3(_0790_),
    .A4(_0823_),
    .ZN(_0824_));
 XNOR2_X1 _3102_ (.A(net223),
    .B(_0824_),
    .ZN(_0825_));
 NOR2_X1 _3103_ (.A1(_0801_),
    .A2(_0825_),
    .ZN(_0231_));
 INV_X2 _3104_ (.A(\prev_event_inc[2] ),
    .ZN(_0826_));
 BUF_X2 _3105_ (.A(event_inc[2]),
    .Z(_0827_));
 NAND3_X1 _3106_ (.A1(_1511_),
    .A2(_0826_),
    .A3(_0827_),
    .ZN(_0828_));
 MUX2_X1 _3107_ (.A(_0002_),
    .B(net224),
    .S(_0828_),
    .Z(_0829_));
 AND2_X1 _3108_ (.A1(_1347_),
    .A2(_0829_),
    .ZN(_0232_));
 MUX2_X1 _3109_ (.A(_0003_),
    .B(net225),
    .S(_0828_),
    .Z(_0830_));
 AND2_X1 _3110_ (.A1(_1347_),
    .A2(_0830_),
    .ZN(_0233_));
 INV_X1 _3111_ (.A(net226),
    .ZN(_0831_));
 NAND4_X2 _3112_ (.A1(_1511_),
    .A2(_0826_),
    .A3(_0827_),
    .A4(_1932_),
    .ZN(_0832_));
 XNOR2_X1 _3113_ (.A(_0831_),
    .B(_0832_),
    .ZN(_0833_));
 NOR2_X1 _3114_ (.A1(_0801_),
    .A2(_0833_),
    .ZN(_0234_));
 BUF_X4 _3115_ (.A(net227),
    .Z(_0834_));
 AND2_X1 _3116_ (.A1(net224),
    .A2(net225),
    .ZN(_0835_));
 NAND4_X4 _3117_ (.A1(_1351_),
    .A2(_0826_),
    .A3(_0827_),
    .A4(_0835_),
    .ZN(_0836_));
 NOR2_X1 _3118_ (.A1(_0831_),
    .A2(_0836_),
    .ZN(_0837_));
 XNOR2_X1 _3119_ (.A(_0834_),
    .B(_0837_),
    .ZN(_0838_));
 NOR2_X1 _3120_ (.A1(_0801_),
    .A2(_0838_),
    .ZN(_0235_));
 NAND2_X1 _3121_ (.A1(net226),
    .A2(_0834_),
    .ZN(_0839_));
 NOR2_X1 _3122_ (.A1(_0832_),
    .A2(_0839_),
    .ZN(_0840_));
 XNOR2_X1 _3123_ (.A(net228),
    .B(_0840_),
    .ZN(_0841_));
 NOR2_X1 _3124_ (.A1(_0801_),
    .A2(_0841_),
    .ZN(_0236_));
 CLKBUF_X3 _3125_ (.A(_1447_),
    .Z(_0842_));
 INV_X1 _3126_ (.A(net228),
    .ZN(_0843_));
 NOR3_X1 _3127_ (.A1(_0843_),
    .A2(_0836_),
    .A3(_0839_),
    .ZN(_0844_));
 XNOR2_X1 _3128_ (.A(net229),
    .B(_0844_),
    .ZN(_0845_));
 NOR2_X1 _3129_ (.A1(_0842_),
    .A2(_0845_),
    .ZN(_0237_));
 XNOR2_X1 _3130_ (.A(_1419_),
    .B(_1418_),
    .ZN(_0846_));
 NOR2_X1 _3131_ (.A1(_0842_),
    .A2(_0846_),
    .ZN(_0238_));
 BUF_X1 _3132_ (.A(net231),
    .Z(_0847_));
 NAND2_X1 _3133_ (.A1(_0827_),
    .A2(_1932_),
    .ZN(_0848_));
 NAND4_X4 _3134_ (.A1(net226),
    .A2(_0834_),
    .A3(net228),
    .A4(net229),
    .ZN(_0849_));
 NOR4_X4 _3135_ (.A1(_1369_),
    .A2(\prev_event_inc[2] ),
    .A3(_0848_),
    .A4(_0849_),
    .ZN(_0850_));
 XNOR2_X1 _3136_ (.A(_0847_),
    .B(_0850_),
    .ZN(_0851_));
 NOR2_X1 _3137_ (.A1(_0842_),
    .A2(_0851_),
    .ZN(_0239_));
 BUF_X1 _3138_ (.A(net232),
    .Z(_0852_));
 INV_X1 _3139_ (.A(_0847_),
    .ZN(_0853_));
 NOR3_X1 _3140_ (.A1(_0853_),
    .A2(_0836_),
    .A3(_0849_),
    .ZN(_0854_));
 XNOR2_X1 _3141_ (.A(_0852_),
    .B(_0854_),
    .ZN(_0855_));
 NOR2_X1 _3142_ (.A1(_0842_),
    .A2(_0855_),
    .ZN(_0240_));
 INV_X1 _3143_ (.A(net233),
    .ZN(_0856_));
 NAND3_X1 _3144_ (.A1(_0847_),
    .A2(_0852_),
    .A3(_0850_),
    .ZN(_0857_));
 XNOR2_X1 _3145_ (.A(_0856_),
    .B(_0857_),
    .ZN(_0858_));
 NOR2_X1 _3146_ (.A1(_0842_),
    .A2(_0858_),
    .ZN(_0241_));
 NAND3_X1 _3147_ (.A1(_0847_),
    .A2(_0852_),
    .A3(net233),
    .ZN(_0859_));
 NOR3_X1 _3148_ (.A1(_0836_),
    .A2(_0849_),
    .A3(_0859_),
    .ZN(_0860_));
 XNOR2_X1 _3149_ (.A(net234),
    .B(_0860_),
    .ZN(_0861_));
 NOR2_X1 _3150_ (.A1(_0842_),
    .A2(_0861_),
    .ZN(_0242_));
 INV_X1 _3151_ (.A(net235),
    .ZN(_0862_));
 AND4_X1 _3152_ (.A1(_0847_),
    .A2(_0852_),
    .A3(net233),
    .A4(net234),
    .ZN(_0863_));
 NAND2_X1 _3153_ (.A1(_0850_),
    .A2(_0863_),
    .ZN(_0864_));
 XNOR2_X1 _3154_ (.A(_0862_),
    .B(_0864_),
    .ZN(_0865_));
 NOR2_X1 _3155_ (.A1(_0842_),
    .A2(_0865_),
    .ZN(_0243_));
 INV_X1 _3156_ (.A(net236),
    .ZN(_0866_));
 NAND2_X1 _3157_ (.A1(net235),
    .A2(_0863_),
    .ZN(_0867_));
 OR3_X2 _3158_ (.A1(_0836_),
    .A2(_0849_),
    .A3(_0867_),
    .ZN(_0868_));
 XNOR2_X1 _3159_ (.A(_0866_),
    .B(_0868_),
    .ZN(_0869_));
 NOR2_X1 _3160_ (.A1(_0842_),
    .A2(_0869_),
    .ZN(_0244_));
 BUF_X2 _3161_ (.A(net237),
    .Z(_0870_));
 OR4_X2 _3162_ (.A1(_1369_),
    .A2(\prev_event_inc[2] ),
    .A3(_0848_),
    .A4(_0849_),
    .ZN(_0871_));
 BUF_X8 _3163_ (.A(_0871_),
    .Z(_0872_));
 CLKBUF_X3 _3164_ (.A(_0867_),
    .Z(_0873_));
 NOR3_X1 _3165_ (.A1(_0866_),
    .A2(_0872_),
    .A3(_0873_),
    .ZN(_0874_));
 XNOR2_X1 _3166_ (.A(_0870_),
    .B(_0874_),
    .ZN(_0875_));
 NOR2_X1 _3167_ (.A1(_0842_),
    .A2(_0875_),
    .ZN(_0245_));
 INV_X1 _3168_ (.A(_0827_),
    .ZN(_0876_));
 OR4_X2 _3169_ (.A1(_1369_),
    .A2(\prev_event_inc[2] ),
    .A3(_0876_),
    .A4(_0849_),
    .ZN(_0877_));
 NAND3_X1 _3170_ (.A1(net235),
    .A2(_0835_),
    .A3(_0863_),
    .ZN(_0878_));
 NAND2_X1 _3171_ (.A1(net236),
    .A2(_0870_),
    .ZN(_0879_));
 NOR3_X1 _3172_ (.A1(_0877_),
    .A2(_0878_),
    .A3(_0879_),
    .ZN(_0880_));
 XNOR2_X1 _3173_ (.A(net238),
    .B(_0880_),
    .ZN(_0881_));
 NOR2_X1 _3174_ (.A1(_0842_),
    .A2(_0881_),
    .ZN(_0246_));
 CLKBUF_X3 _3175_ (.A(_1447_),
    .Z(_0882_));
 INV_X1 _3176_ (.A(net238),
    .ZN(_0883_));
 NOR4_X1 _3177_ (.A1(_0883_),
    .A2(_0872_),
    .A3(_0873_),
    .A4(_0879_),
    .ZN(_0884_));
 XNOR2_X1 _3178_ (.A(net239),
    .B(_0884_),
    .ZN(_0885_));
 NOR2_X1 _3179_ (.A1(_0882_),
    .A2(_0885_),
    .ZN(_0247_));
 NAND4_X2 _3180_ (.A1(net236),
    .A2(_0870_),
    .A3(net238),
    .A4(net239),
    .ZN(_0886_));
 OAI21_X1 _3181_ (.A(net240),
    .B1(_0868_),
    .B2(_0886_),
    .ZN(_0887_));
 OR3_X1 _3182_ (.A1(net240),
    .A2(_0868_),
    .A3(_0886_),
    .ZN(_0888_));
 AOI21_X1 _3183_ (.A(_1356_),
    .B1(_0887_),
    .B2(_0888_),
    .ZN(_0248_));
 NAND2_X1 _3184_ (.A1(_1419_),
    .A2(_1470_),
    .ZN(_0889_));
 XOR2_X1 _3185_ (.A(_1420_),
    .B(_0889_),
    .Z(_0890_));
 NOR2_X1 _3186_ (.A1(_0882_),
    .A2(_0890_),
    .ZN(_0249_));
 INV_X1 _3187_ (.A(net240),
    .ZN(_0891_));
 NOR4_X1 _3188_ (.A1(_0891_),
    .A2(_0872_),
    .A3(_0873_),
    .A4(_0886_),
    .ZN(_0892_));
 XNOR2_X1 _3189_ (.A(net242),
    .B(_0892_),
    .ZN(_0893_));
 NOR2_X1 _3190_ (.A1(_0882_),
    .A2(_0893_),
    .ZN(_0250_));
 BUF_X2 _3191_ (.A(net243),
    .Z(_0894_));
 NAND2_X1 _3192_ (.A1(net240),
    .A2(net242),
    .ZN(_0895_));
 OR2_X1 _3193_ (.A1(_0886_),
    .A2(_0895_),
    .ZN(_0896_));
 NOR3_X1 _3194_ (.A1(_0877_),
    .A2(_0878_),
    .A3(_0896_),
    .ZN(_0897_));
 XNOR2_X1 _3195_ (.A(_0894_),
    .B(_0897_),
    .ZN(_0898_));
 NOR2_X1 _3196_ (.A1(_0882_),
    .A2(_0898_),
    .ZN(_0251_));
 BUF_X4 _3197_ (.A(net244),
    .Z(_0899_));
 INV_X1 _3198_ (.A(_0894_),
    .ZN(_0900_));
 NOR4_X1 _3199_ (.A1(_0900_),
    .A2(_0872_),
    .A3(_0873_),
    .A4(_0896_),
    .ZN(_0901_));
 XNOR2_X1 _3200_ (.A(_0899_),
    .B(_0901_),
    .ZN(_0902_));
 NOR2_X1 _3201_ (.A1(_0882_),
    .A2(_0902_),
    .ZN(_0252_));
 INV_X1 _3202_ (.A(net245),
    .ZN(_0903_));
 NOR2_X1 _3203_ (.A1(_0903_),
    .A2(_1474_),
    .ZN(_0904_));
 NOR2_X1 _3204_ (.A1(net245),
    .A2(_1490_),
    .ZN(_0905_));
 AND3_X1 _3205_ (.A1(_0894_),
    .A2(_0899_),
    .A3(_0897_),
    .ZN(_0906_));
 MUX2_X1 _3206_ (.A(_0904_),
    .B(_0905_),
    .S(_0906_),
    .Z(_0253_));
 NAND3_X1 _3207_ (.A1(_0894_),
    .A2(_0899_),
    .A3(net245),
    .ZN(_0907_));
 NOR4_X1 _3208_ (.A1(_0872_),
    .A2(_0873_),
    .A3(_0896_),
    .A4(_0907_),
    .ZN(_0908_));
 XNOR2_X1 _3209_ (.A(net246),
    .B(_0908_),
    .ZN(_0909_));
 NOR2_X1 _3210_ (.A1(_0882_),
    .A2(_0909_),
    .ZN(_0254_));
 INV_X1 _3211_ (.A(net247),
    .ZN(_0910_));
 NOR2_X1 _3212_ (.A1(_0910_),
    .A2(_1474_),
    .ZN(_0911_));
 NOR2_X1 _3213_ (.A1(net247),
    .A2(_1490_),
    .ZN(_0912_));
 NAND4_X2 _3214_ (.A1(_0894_),
    .A2(_0899_),
    .A3(net245),
    .A4(net246),
    .ZN(_0913_));
 NOR3_X1 _3215_ (.A1(_0868_),
    .A2(_0896_),
    .A3(_0913_),
    .ZN(_0914_));
 MUX2_X1 _3216_ (.A(_0911_),
    .B(_0912_),
    .S(_0914_),
    .Z(_0255_));
 OR2_X1 _3217_ (.A1(_0910_),
    .A2(_0913_),
    .ZN(_0915_));
 NOR4_X1 _3218_ (.A1(_0872_),
    .A2(_0873_),
    .A3(_0896_),
    .A4(_0915_),
    .ZN(_0916_));
 XNOR2_X1 _3219_ (.A(net248),
    .B(_0916_),
    .ZN(_0917_));
 NOR2_X1 _3220_ (.A1(_0882_),
    .A2(_0917_),
    .ZN(_0256_));
 INV_X1 _3221_ (.A(net249),
    .ZN(_0918_));
 NAND2_X1 _3222_ (.A1(net247),
    .A2(net248),
    .ZN(_0919_));
 OR4_X2 _3223_ (.A1(_0886_),
    .A2(_0895_),
    .A3(_0913_),
    .A4(_0919_),
    .ZN(_0920_));
 OR3_X2 _3224_ (.A1(_0877_),
    .A2(_0878_),
    .A3(_0920_),
    .ZN(_0921_));
 XNOR2_X1 _3225_ (.A(_0918_),
    .B(_0921_),
    .ZN(_0922_));
 NOR2_X1 _3226_ (.A1(_0882_),
    .A2(_0922_),
    .ZN(_0257_));
 NOR4_X1 _3227_ (.A1(_0918_),
    .A2(_0872_),
    .A3(_0873_),
    .A4(_0920_),
    .ZN(_0923_));
 XNOR2_X1 _3228_ (.A(net250),
    .B(_0923_),
    .ZN(_0924_));
 NOR2_X1 _3229_ (.A1(_0882_),
    .A2(_0924_),
    .ZN(_0258_));
 INV_X1 _3230_ (.A(net251),
    .ZN(_0925_));
 NOR2_X1 _3231_ (.A1(_0925_),
    .A2(_1474_),
    .ZN(_0926_));
 NOR2_X1 _3232_ (.A1(net251),
    .A2(_1490_),
    .ZN(_0927_));
 INV_X1 _3233_ (.A(net250),
    .ZN(_0928_));
 NOR3_X1 _3234_ (.A1(_0918_),
    .A2(_0928_),
    .A3(_0921_),
    .ZN(_0929_));
 MUX2_X1 _3235_ (.A(_0926_),
    .B(_0927_),
    .S(_0929_),
    .Z(_0259_));
 NAND3_X1 _3236_ (.A1(_1419_),
    .A2(_1420_),
    .A3(_1418_),
    .ZN(_0930_));
 XOR2_X1 _3237_ (.A(net252),
    .B(_0930_),
    .Z(_0931_));
 NOR2_X1 _3238_ (.A1(_0882_),
    .A2(_0931_),
    .ZN(_0260_));
 NAND3_X1 _3239_ (.A1(net249),
    .A2(net250),
    .A3(net251),
    .ZN(_0932_));
 NOR4_X1 _3240_ (.A1(_0872_),
    .A2(_0873_),
    .A3(_0920_),
    .A4(_0932_),
    .ZN(_0933_));
 XNOR2_X1 _3241_ (.A(net253),
    .B(_0933_),
    .ZN(_0934_));
 NOR2_X1 _3242_ (.A1(_1448_),
    .A2(_0934_),
    .ZN(_0261_));
 BUF_X1 _3243_ (.A(net254),
    .Z(_0935_));
 INV_X1 _3244_ (.A(_0935_),
    .ZN(_0936_));
 NOR2_X1 _3245_ (.A1(_0936_),
    .A2(_1474_),
    .ZN(_0937_));
 NOR2_X1 _3246_ (.A1(_0935_),
    .A2(_1490_),
    .ZN(_0938_));
 INV_X1 _3247_ (.A(net253),
    .ZN(_0939_));
 NOR3_X1 _3248_ (.A1(_0939_),
    .A2(_0921_),
    .A3(_0932_),
    .ZN(_0940_));
 MUX2_X1 _3249_ (.A(_0937_),
    .B(_0938_),
    .S(_0940_),
    .Z(_0262_));
 BUF_X1 _3250_ (.A(net255),
    .Z(_0941_));
 AND4_X1 _3251_ (.A1(net249),
    .A2(net250),
    .A3(net251),
    .A4(net253),
    .ZN(_0942_));
 NAND2_X1 _3252_ (.A1(_0935_),
    .A2(_0942_),
    .ZN(_0943_));
 NOR4_X1 _3253_ (.A1(_0872_),
    .A2(_0873_),
    .A3(_0920_),
    .A4(_0943_),
    .ZN(_0944_));
 XNOR2_X1 _3254_ (.A(_0941_),
    .B(_0944_),
    .ZN(_0945_));
 NOR2_X1 _3255_ (.A1(_1448_),
    .A2(_0945_),
    .ZN(_0263_));
 NAND3_X1 _3256_ (.A1(_0935_),
    .A2(_0941_),
    .A3(_0942_),
    .ZN(_0946_));
 OAI21_X1 _3257_ (.A(net256),
    .B1(_0921_),
    .B2(_0946_),
    .ZN(_0947_));
 OR3_X1 _3258_ (.A1(net256),
    .A2(_0921_),
    .A3(_0946_),
    .ZN(_0948_));
 AOI21_X1 _3259_ (.A(_1356_),
    .B1(_0947_),
    .B2(_0948_),
    .ZN(_0264_));
 NAND4_X1 _3260_ (.A1(_0935_),
    .A2(_0941_),
    .A3(net256),
    .A4(_0942_),
    .ZN(_0949_));
 NOR4_X1 _3261_ (.A1(_0872_),
    .A2(_0873_),
    .A3(_0920_),
    .A4(_0949_),
    .ZN(_0950_));
 XNOR2_X1 _3262_ (.A(net257),
    .B(_0950_),
    .ZN(_0951_));
 NOR2_X1 _3263_ (.A1(_1448_),
    .A2(_0951_),
    .ZN(_0265_));
 INV_X1 _3264_ (.A(net258),
    .ZN(_0952_));
 NOR2_X1 _3265_ (.A1(_0952_),
    .A2(_1474_),
    .ZN(_0953_));
 NOR2_X1 _3266_ (.A1(net258),
    .A2(_1490_),
    .ZN(_0954_));
 INV_X1 _3267_ (.A(net257),
    .ZN(_0955_));
 NOR3_X1 _3268_ (.A1(_0955_),
    .A2(_0921_),
    .A3(_0949_),
    .ZN(_0956_));
 MUX2_X1 _3269_ (.A(_0953_),
    .B(_0954_),
    .S(_0956_),
    .Z(_0266_));
 MUX2_X1 _3270_ (.A(_0004_),
    .B(net259),
    .S(_1405_),
    .Z(_0957_));
 AND2_X1 _3271_ (.A1(_1347_),
    .A2(_0957_),
    .ZN(_0267_));
 MUX2_X1 _3272_ (.A(_0005_),
    .B(_1370_),
    .S(_1405_),
    .Z(_0958_));
 AND2_X1 _3273_ (.A1(_1347_),
    .A2(_0958_),
    .ZN(_0268_));
 NAND4_X1 _3274_ (.A1(_1511_),
    .A2(_1361_),
    .A3(_1362_),
    .A4(_1926_),
    .ZN(_0959_));
 XOR2_X1 _3275_ (.A(_1363_),
    .B(_0959_),
    .Z(_0960_));
 NOR2_X1 _3276_ (.A1(_1448_),
    .A2(_0960_),
    .ZN(_0269_));
 XNOR2_X1 _3277_ (.A(_1359_),
    .B(_1373_),
    .ZN(_0961_));
 NOR2_X1 _3278_ (.A1(_1448_),
    .A2(_0961_),
    .ZN(_0270_));
 NAND4_X1 _3279_ (.A1(_1419_),
    .A2(_1420_),
    .A3(net252),
    .A4(_1469_),
    .ZN(_0962_));
 XOR2_X1 _3280_ (.A(net263),
    .B(_0962_),
    .Z(_0963_));
 NOR2_X1 _3281_ (.A1(_1448_),
    .A2(_0963_),
    .ZN(_0271_));
 NAND2_X1 _3282_ (.A1(\prev_event_inc[0] ),
    .A2(_1344_),
    .ZN(_0964_));
 NAND2_X1 _3283_ (.A1(net3),
    .A2(_1354_),
    .ZN(_0965_));
 AOI21_X1 _3284_ (.A(_1345_),
    .B1(_0964_),
    .B2(_0965_),
    .ZN(_0272_));
 NAND2_X1 _3285_ (.A1(\prev_event_inc[1] ),
    .A2(_1344_),
    .ZN(_0966_));
 NAND2_X1 _3286_ (.A1(net4),
    .A2(_1354_),
    .ZN(_0967_));
 AOI21_X1 _3287_ (.A(_1345_),
    .B1(_0966_),
    .B2(_0967_),
    .ZN(_0273_));
 MUX2_X1 _3288_ (.A(_0826_),
    .B(_0876_),
    .S(_1354_),
    .Z(_0968_));
 NOR2_X1 _3289_ (.A1(_1345_),
    .A2(_0968_),
    .ZN(_0274_));
 NAND2_X1 _3290_ (.A1(\prev_event_inc[3] ),
    .A2(_1344_),
    .ZN(_0969_));
 NAND2_X1 _3291_ (.A1(_1362_),
    .A2(_1354_),
    .ZN(_0970_));
 AOI21_X1 _3292_ (.A(_1345_),
    .B1(_0969_),
    .B2(_0970_),
    .ZN(_0275_));
 NAND2_X1 _3293_ (.A1(\prev_event_inc[4] ),
    .A2(_1344_),
    .ZN(_0971_));
 NAND2_X1 _3294_ (.A1(_1513_),
    .A2(_1354_),
    .ZN(_0972_));
 AOI21_X1 _3295_ (.A(_1345_),
    .B1(_0971_),
    .B2(_0972_),
    .ZN(_0276_));
 MUX2_X1 _3296_ (.A(_1652_),
    .B(_1661_),
    .S(_1354_),
    .Z(_0973_));
 NOR2_X1 _3297_ (.A1(_1345_),
    .A2(_0973_),
    .ZN(_0277_));
 NAND2_X1 _3298_ (.A1(\prev_event_inc[6] ),
    .A2(_1344_),
    .ZN(_0974_));
 NAND2_X1 _3299_ (.A1(net6),
    .A2(_1354_),
    .ZN(_0975_));
 AOI21_X1 _3300_ (.A(_1345_),
    .B1(_0974_),
    .B2(_0975_),
    .ZN(_0278_));
 MUX2_X1 _3301_ (.A(_0536_),
    .B(_0523_),
    .S(_1354_),
    .Z(_0976_));
 NOR2_X1 _3302_ (.A1(_1345_),
    .A2(_0976_),
    .ZN(_0279_));
 INV_X2 _3303_ (.A(net1),
    .ZN(_0977_));
 BUF_X4 _3304_ (.A(net2),
    .Z(_0978_));
 BUF_X4 _3305_ (.A(_0978_),
    .Z(_0979_));
 NOR3_X2 _3306_ (.A1(net110),
    .A2(_0977_),
    .A3(_0979_),
    .ZN(_0980_));
 OR2_X1 _3307_ (.A1(net1),
    .A2(net2),
    .ZN(_0981_));
 BUF_X2 _3308_ (.A(_0981_),
    .Z(_0982_));
 BUF_X2 _3309_ (.A(_0982_),
    .Z(_0983_));
 CLKBUF_X3 _3310_ (.A(counter_sel[5]),
    .Z(_0984_));
 BUF_X2 _3311_ (.A(_0984_),
    .Z(_0985_));
 AOI21_X1 _3312_ (.A(_0983_),
    .B1(_0985_),
    .B2(net75),
    .ZN(_0986_));
 BUF_X2 _3313_ (.A(_0984_),
    .Z(_0987_));
 CLKBUF_X3 _3314_ (.A(counter_sel[4]),
    .Z(_0988_));
 BUF_X4 _3315_ (.A(_0988_),
    .Z(_0989_));
 CLKBUF_X3 _3316_ (.A(counter_sel[2]),
    .Z(_0990_));
 CLKBUF_X3 _3317_ (.A(_0990_),
    .Z(_0991_));
 CLKBUF_X3 _3318_ (.A(counter_sel[1]),
    .Z(_0992_));
 BUF_X2 _3319_ (.A(_0992_),
    .Z(_0993_));
 AOI21_X1 _3320_ (.A(_0991_),
    .B1(_0993_),
    .B2(net189),
    .ZN(_0994_));
 BUF_X1 _3321_ (.A(counter_sel[0]),
    .Z(_0995_));
 BUF_X2 _3322_ (.A(_0995_),
    .Z(_0996_));
 NAND2_X1 _3323_ (.A1(_0996_),
    .A2(net8),
    .ZN(_0997_));
 BUF_X2 _3324_ (.A(_0992_),
    .Z(_0998_));
 OAI21_X1 _3325_ (.A(_0994_),
    .B1(_0997_),
    .B2(_0998_),
    .ZN(_0999_));
 CLKBUF_X3 _3326_ (.A(counter_sel[3]),
    .Z(_1000_));
 BUF_X4 _3327_ (.A(_1000_),
    .Z(_1001_));
 BUF_X2 _3328_ (.A(_0990_),
    .Z(_1002_));
 INV_X1 _3329_ (.A(net224),
    .ZN(_1003_));
 AOI21_X1 _3330_ (.A(_1001_),
    .B1(_1002_),
    .B2(_1003_),
    .ZN(_1004_));
 BUF_X4 _3331_ (.A(_1001_),
    .Z(_1005_));
 AOI221_X2 _3332_ (.A(_0989_),
    .B1(_0999_),
    .B2(_1004_),
    .C1(_1005_),
    .C2(net259),
    .ZN(_1006_));
 INV_X1 _3333_ (.A(_0989_),
    .ZN(_1007_));
 NOR2_X1 _3334_ (.A1(net39),
    .A2(_1007_),
    .ZN(_1008_));
 OR3_X1 _3335_ (.A1(_0987_),
    .A2(_1006_),
    .A3(_1008_),
    .ZN(_1009_));
 BUF_X4 _3336_ (.A(_0979_),
    .Z(_1010_));
 AOI221_X2 _3337_ (.A(_0980_),
    .B1(_0986_),
    .B2(_1009_),
    .C1(_0521_),
    .C2(_1010_),
    .ZN(net264));
 BUF_X4 _3338_ (.A(_0977_),
    .Z(_1011_));
 NOR3_X2 _3339_ (.A1(_1011_),
    .A2(net122),
    .A3(_0979_),
    .ZN(_1012_));
 AOI21_X1 _3340_ (.A(_0983_),
    .B1(_0301_),
    .B2(_0985_),
    .ZN(_1013_));
 AOI21_X1 _3341_ (.A(_0991_),
    .B1(net200),
    .B2(_0993_),
    .ZN(_1014_));
 NAND2_X1 _3342_ (.A1(_0996_),
    .A2(net19),
    .ZN(_1015_));
 OAI21_X1 _3343_ (.A(_1014_),
    .B1(_1015_),
    .B2(_0998_),
    .ZN(_1016_));
 AOI21_X1 _3344_ (.A(_1001_),
    .B1(_0862_),
    .B2(_1002_),
    .ZN(_1017_));
 AOI221_X2 _3345_ (.A(_0989_),
    .B1(_1016_),
    .B2(_1017_),
    .C1(net15),
    .C2(_1005_),
    .ZN(_1018_));
 CLKBUF_X3 _3346_ (.A(_1007_),
    .Z(_1019_));
 NOR2_X1 _3347_ (.A1(_1019_),
    .A2(net50),
    .ZN(_1020_));
 OR3_X1 _3348_ (.A1(_0987_),
    .A2(_1018_),
    .A3(_1020_),
    .ZN(_1021_));
 AOI221_X2 _3349_ (.A(_1012_),
    .B1(_1013_),
    .B2(_1021_),
    .C1(_0572_),
    .C2(_1010_),
    .ZN(net265));
 NOR3_X2 _3350_ (.A1(_1011_),
    .A2(_0431_),
    .A3(_0979_),
    .ZN(_1022_));
 AOI21_X1 _3351_ (.A(_0983_),
    .B1(net87),
    .B2(_0985_),
    .ZN(_1023_));
 AOI21_X1 _3352_ (.A(_0991_),
    .B1(net201),
    .B2(_0993_),
    .ZN(_1024_));
 NAND2_X1 _3353_ (.A1(_0996_),
    .A2(net30),
    .ZN(_1025_));
 OAI21_X1 _3354_ (.A(_1024_),
    .B1(_1025_),
    .B2(_0998_),
    .ZN(_1026_));
 AOI21_X1 _3355_ (.A(_1001_),
    .B1(_0866_),
    .B2(_1002_),
    .ZN(_1027_));
 AOI221_X2 _3356_ (.A(_0989_),
    .B1(_1026_),
    .B2(_1027_),
    .C1(_1395_),
    .C2(_1005_),
    .ZN(_1028_));
 NOR2_X1 _3357_ (.A1(_1019_),
    .A2(_1561_),
    .ZN(_1029_));
 OR3_X1 _3358_ (.A1(_0987_),
    .A2(_1028_),
    .A3(_1029_),
    .ZN(_1030_));
 INV_X1 _3359_ (.A(_0571_),
    .ZN(_1031_));
 AOI221_X2 _3360_ (.A(_1022_),
    .B1(_1023_),
    .B2(_1030_),
    .C1(_1031_),
    .C2(_1010_),
    .ZN(net266));
 NOR3_X2 _3361_ (.A1(_1011_),
    .A2(net124),
    .A3(_0979_),
    .ZN(_1032_));
 AOI21_X1 _3362_ (.A(_0983_),
    .B1(_0307_),
    .B2(_0985_),
    .ZN(_1033_));
 AOI21_X1 _3363_ (.A(_0991_),
    .B1(_0741_),
    .B2(_0993_),
    .ZN(_1034_));
 NAND2_X1 _3364_ (.A1(_0996_),
    .A2(_1517_),
    .ZN(_1035_));
 OAI21_X1 _3365_ (.A(_1034_),
    .B1(_1035_),
    .B2(_0998_),
    .ZN(_1036_));
 INV_X1 _3366_ (.A(_0870_),
    .ZN(_1037_));
 AOI21_X1 _3367_ (.A(_1001_),
    .B1(_1037_),
    .B2(_1002_),
    .ZN(_1038_));
 AOI221_X2 _3368_ (.A(_0989_),
    .B1(_1036_),
    .B2(_1038_),
    .C1(_1399_),
    .C2(_1005_),
    .ZN(_1039_));
 NOR2_X1 _3369_ (.A1(_1019_),
    .A2(_1568_),
    .ZN(_1040_));
 OR3_X1 _3370_ (.A1(_0987_),
    .A2(_1039_),
    .A3(_1040_),
    .ZN(_1041_));
 AOI221_X2 _3371_ (.A(_1032_),
    .B1(_1033_),
    .B2(_1041_),
    .C1(_0575_),
    .C2(_1010_),
    .ZN(net267));
 NOR3_X2 _3372_ (.A1(_1011_),
    .A2(net125),
    .A3(_0979_),
    .ZN(_1042_));
 AOI21_X1 _3373_ (.A(_0983_),
    .B1(_0312_),
    .B2(_0985_),
    .ZN(_1043_));
 AOI21_X1 _3374_ (.A(_0991_),
    .B1(net203),
    .B2(_0993_),
    .ZN(_1044_));
 NAND2_X1 _3375_ (.A1(_0996_),
    .A2(_1565_),
    .ZN(_1045_));
 OAI21_X1 _3376_ (.A(_1044_),
    .B1(_1045_),
    .B2(_0998_),
    .ZN(_1046_));
 AOI21_X1 _3377_ (.A(_1001_),
    .B1(_0883_),
    .B2(_1002_),
    .ZN(_1047_));
 AOI221_X2 _3378_ (.A(_0989_),
    .B1(_1046_),
    .B2(_1047_),
    .C1(_1403_),
    .C2(_1005_),
    .ZN(_1048_));
 NOR2_X1 _3379_ (.A1(_1019_),
    .A2(_1571_),
    .ZN(_1049_));
 OR3_X1 _3380_ (.A1(_0987_),
    .A2(_1048_),
    .A3(_1049_),
    .ZN(_1050_));
 AOI221_X2 _3381_ (.A(_1042_),
    .B1(_1043_),
    .B2(_1050_),
    .C1(_0581_),
    .C2(_1010_),
    .ZN(net268));
 BUF_X4 _3382_ (.A(_0978_),
    .Z(_1051_));
 NOR3_X2 _3383_ (.A1(_1011_),
    .A2(net126),
    .A3(_1051_),
    .ZN(_1052_));
 AOI21_X1 _3384_ (.A(_0983_),
    .B1(net90),
    .B2(_0985_),
    .ZN(_1053_));
 AOI21_X1 _3385_ (.A(_0991_),
    .B1(_0749_),
    .B2(_0993_),
    .ZN(_1054_));
 NAND2_X1 _3386_ (.A1(_0996_),
    .A2(_1607_),
    .ZN(_1055_));
 OAI21_X1 _3387_ (.A(_1054_),
    .B1(_1055_),
    .B2(_0998_),
    .ZN(_1056_));
 CLKBUF_X3 _3388_ (.A(_1000_),
    .Z(_1057_));
 INV_X1 _3389_ (.A(net239),
    .ZN(_1058_));
 AOI21_X1 _3390_ (.A(_1057_),
    .B1(_1058_),
    .B2(_1002_),
    .ZN(_1059_));
 AOI221_X2 _3391_ (.A(_0989_),
    .B1(_1056_),
    .B2(_1059_),
    .C1(_1424_),
    .C2(_1005_),
    .ZN(_1060_));
 NOR2_X1 _3392_ (.A1(_1019_),
    .A2(net55),
    .ZN(_1061_));
 OR3_X1 _3393_ (.A1(_0987_),
    .A2(_1060_),
    .A3(_1061_),
    .ZN(_1062_));
 AOI221_X2 _3394_ (.A(_1052_),
    .B1(_1053_),
    .B2(_1062_),
    .C1(_0584_),
    .C2(_1010_),
    .ZN(net269));
 NOR3_X2 _3395_ (.A1(_1011_),
    .A2(net127),
    .A3(_1051_),
    .ZN(_1063_));
 AOI21_X1 _3396_ (.A(_0983_),
    .B1(_0317_),
    .B2(_0985_),
    .ZN(_1064_));
 AOI21_X1 _3397_ (.A(_0991_),
    .B1(net205),
    .B2(_0993_),
    .ZN(_1065_));
 NAND2_X1 _3398_ (.A1(_0996_),
    .A2(net74),
    .ZN(_1066_));
 OAI21_X1 _3399_ (.A(_1065_),
    .B1(_1066_),
    .B2(_0998_),
    .ZN(_1067_));
 AOI21_X1 _3400_ (.A(_1057_),
    .B1(_0891_),
    .B2(_1002_),
    .ZN(_1068_));
 AOI221_X2 _3401_ (.A(_0989_),
    .B1(_1067_),
    .B2(_1068_),
    .C1(net21),
    .C2(_1005_),
    .ZN(_1069_));
 NOR2_X1 _3402_ (.A1(_1019_),
    .A2(_1579_),
    .ZN(_1070_));
 OR3_X1 _3403_ (.A1(_0987_),
    .A2(_1069_),
    .A3(_1070_),
    .ZN(_1071_));
 AOI221_X2 _3404_ (.A(_1063_),
    .B1(_1064_),
    .B2(_1071_),
    .C1(_0588_),
    .C2(_1010_),
    .ZN(net270));
 NOR3_X2 _3405_ (.A1(_1011_),
    .A2(net128),
    .A3(_1051_),
    .ZN(_1072_));
 AOI21_X1 _3406_ (.A(_0983_),
    .B1(net92),
    .B2(_0985_),
    .ZN(_1073_));
 AOI21_X1 _3407_ (.A(_0991_),
    .B1(net206),
    .B2(_0993_),
    .ZN(_1074_));
 NAND2_X1 _3408_ (.A1(_0996_),
    .A2(_0297_),
    .ZN(_1075_));
 OAI21_X1 _3409_ (.A(_1074_),
    .B1(_1075_),
    .B2(_0998_),
    .ZN(_1076_));
 INV_X1 _3410_ (.A(net242),
    .ZN(_1077_));
 AOI21_X1 _3411_ (.A(_1057_),
    .B1(_1077_),
    .B2(_1002_),
    .ZN(_1078_));
 AOI221_X2 _3412_ (.A(_0989_),
    .B1(_1076_),
    .B2(_1078_),
    .C1(net22),
    .C2(_1005_),
    .ZN(_1079_));
 NOR2_X1 _3413_ (.A1(_1019_),
    .A2(_1584_),
    .ZN(_1080_));
 OR3_X1 _3414_ (.A1(_0987_),
    .A2(_1079_),
    .A3(_1080_),
    .ZN(_1081_));
 AOI221_X2 _3415_ (.A(_1072_),
    .B1(_1073_),
    .B2(_1081_),
    .C1(_0596_),
    .C2(_1010_),
    .ZN(net271));
 NOR3_X2 _3416_ (.A1(_1011_),
    .A2(net129),
    .A3(_1051_),
    .ZN(_1082_));
 AOI21_X1 _3417_ (.A(_0983_),
    .B1(_0324_),
    .B2(_0985_),
    .ZN(_1083_));
 BUF_X2 _3418_ (.A(_0984_),
    .Z(_1084_));
 BUF_X2 _3419_ (.A(_0990_),
    .Z(_1085_));
 CLKBUF_X3 _3420_ (.A(_0992_),
    .Z(_1086_));
 AOI21_X1 _3421_ (.A(_1085_),
    .B1(net207),
    .B2(_1086_),
    .ZN(_1087_));
 NAND2_X1 _3422_ (.A1(_0996_),
    .A2(net96),
    .ZN(_1088_));
 OAI21_X1 _3423_ (.A(_1087_),
    .B1(_1088_),
    .B2(_0998_),
    .ZN(_1089_));
 AOI21_X1 _3424_ (.A(_1057_),
    .B1(_0900_),
    .B2(_1002_),
    .ZN(_1090_));
 AOI221_X2 _3425_ (.A(_0989_),
    .B1(_1089_),
    .B2(_1090_),
    .C1(_1438_),
    .C2(_1005_),
    .ZN(_1091_));
 NOR2_X1 _3426_ (.A1(_1019_),
    .A2(net58),
    .ZN(_1092_));
 OR3_X1 _3427_ (.A1(_1084_),
    .A2(_1091_),
    .A3(_1092_),
    .ZN(_1093_));
 AOI221_X2 _3428_ (.A(_1082_),
    .B1(_1083_),
    .B2(_1093_),
    .C1(_0600_),
    .C2(_1010_),
    .ZN(net272));
 NOR3_X2 _3429_ (.A1(_1011_),
    .A2(_0461_),
    .A3(_1051_),
    .ZN(_1094_));
 AOI21_X1 _3430_ (.A(_0983_),
    .B1(_0329_),
    .B2(_0985_),
    .ZN(_1095_));
 BUF_X4 _3431_ (.A(_0988_),
    .Z(_1096_));
 AOI21_X1 _3432_ (.A(_1085_),
    .B1(_0769_),
    .B2(_1086_),
    .ZN(_1097_));
 NAND2_X1 _3433_ (.A1(_0996_),
    .A2(_0378_),
    .ZN(_1098_));
 OAI21_X1 _3434_ (.A(_1097_),
    .B1(_1098_),
    .B2(_0998_),
    .ZN(_1099_));
 INV_X1 _3435_ (.A(_0899_),
    .ZN(_1100_));
 AOI21_X1 _3436_ (.A(_1057_),
    .B1(_1100_),
    .B2(_1002_),
    .ZN(_1101_));
 AOI221_X2 _3437_ (.A(_1096_),
    .B1(_1099_),
    .B2(_1101_),
    .C1(_1443_),
    .C2(_1005_),
    .ZN(_1102_));
 NOR2_X1 _3438_ (.A1(_1019_),
    .A2(net59),
    .ZN(_1103_));
 OR3_X1 _3439_ (.A1(_1084_),
    .A2(_1102_),
    .A3(_1103_),
    .ZN(_1104_));
 AOI221_X2 _3440_ (.A(_1094_),
    .B1(_1095_),
    .B2(_1104_),
    .C1(_0603_),
    .C2(_1010_),
    .ZN(net273));
 NOR3_X2 _3441_ (.A1(_1011_),
    .A2(_0466_),
    .A3(_1051_),
    .ZN(_1105_));
 CLKBUF_X3 _3442_ (.A(_0982_),
    .Z(_1106_));
 CLKBUF_X3 _3443_ (.A(_0984_),
    .Z(_1107_));
 AOI21_X1 _3444_ (.A(_1106_),
    .B1(_0332_),
    .B2(_1107_),
    .ZN(_1108_));
 AOI21_X1 _3445_ (.A(_1085_),
    .B1(_0774_),
    .B2(_1086_),
    .ZN(_1109_));
 BUF_X2 _3446_ (.A(_0995_),
    .Z(_1110_));
 NAND2_X1 _3447_ (.A1(_1110_),
    .A2(net118),
    .ZN(_1111_));
 BUF_X2 _3448_ (.A(_0992_),
    .Z(_1112_));
 OAI21_X1 _3449_ (.A(_1109_),
    .B1(_1111_),
    .B2(_1112_),
    .ZN(_1113_));
 CLKBUF_X3 _3450_ (.A(_0990_),
    .Z(_1114_));
 AOI21_X1 _3451_ (.A(_1057_),
    .B1(_0903_),
    .B2(_1114_),
    .ZN(_1115_));
 BUF_X4 _3452_ (.A(_1001_),
    .Z(_1116_));
 AOI221_X2 _3453_ (.A(_1096_),
    .B1(_1113_),
    .B2(_1115_),
    .C1(_1449_),
    .C2(_1116_),
    .ZN(_1117_));
 NOR2_X1 _3454_ (.A1(_1019_),
    .A2(net60),
    .ZN(_1118_));
 OR3_X1 _3455_ (.A1(_1084_),
    .A2(_1117_),
    .A3(_1118_),
    .ZN(_1119_));
 BUF_X4 _3456_ (.A(_0979_),
    .Z(_1120_));
 AOI221_X2 _3457_ (.A(_1105_),
    .B1(_1108_),
    .B2(_1119_),
    .C1(_0607_),
    .C2(_1120_),
    .ZN(net274));
 BUF_X2 _3458_ (.A(_0977_),
    .Z(_1121_));
 NOR3_X1 _3459_ (.A1(_1121_),
    .A2(net111),
    .A3(_1051_),
    .ZN(_1122_));
 AOI21_X2 _3460_ (.A(_1106_),
    .B1(net76),
    .B2(_1107_),
    .ZN(_1123_));
 AOI21_X1 _3461_ (.A(_1085_),
    .B1(net190),
    .B2(_1086_),
    .ZN(_1124_));
 NAND2_X1 _3462_ (.A1(_1110_),
    .A2(net119),
    .ZN(_1125_));
 OAI21_X1 _3463_ (.A(_1124_),
    .B1(_1125_),
    .B2(_1112_),
    .ZN(_1126_));
 INV_X1 _3464_ (.A(net225),
    .ZN(_1127_));
 AOI21_X1 _3465_ (.A(_1057_),
    .B1(_1127_),
    .B2(_1114_),
    .ZN(_1128_));
 AOI221_X2 _3466_ (.A(_1096_),
    .B1(_1126_),
    .B2(_1128_),
    .C1(_1370_),
    .C2(_1116_),
    .ZN(_1129_));
 CLKBUF_X3 _3467_ (.A(_1007_),
    .Z(_1130_));
 NOR2_X1 _3468_ (.A1(_1130_),
    .A2(net40),
    .ZN(_1131_));
 OR3_X1 _3469_ (.A1(_1084_),
    .A2(_1129_),
    .A3(_1131_),
    .ZN(_1132_));
 INV_X1 _3470_ (.A(net147),
    .ZN(_1133_));
 AOI221_X2 _3471_ (.A(_1122_),
    .B1(_1123_),
    .B2(_1132_),
    .C1(_1133_),
    .C2(_1120_),
    .ZN(net275));
 NOR3_X1 _3472_ (.A1(_1121_),
    .A2(_0469_),
    .A3(_1051_),
    .ZN(_1134_));
 AOI21_X1 _3473_ (.A(_1106_),
    .B1(net97),
    .B2(_1107_),
    .ZN(_1135_));
 AOI21_X1 _3474_ (.A(_1085_),
    .B1(_0778_),
    .B2(_1086_),
    .ZN(_1136_));
 NAND2_X1 _3475_ (.A1(_1110_),
    .A2(net130),
    .ZN(_1137_));
 OAI21_X1 _3476_ (.A(_1136_),
    .B1(_1137_),
    .B2(_1112_),
    .ZN(_1138_));
 INV_X1 _3477_ (.A(net246),
    .ZN(_1139_));
 AOI21_X1 _3478_ (.A(_1057_),
    .B1(_1139_),
    .B2(_1114_),
    .ZN(_1140_));
 AOI221_X2 _3479_ (.A(_1096_),
    .B1(_1138_),
    .B2(_1140_),
    .C1(net26),
    .C2(_1116_),
    .ZN(_1141_));
 NOR2_X1 _3480_ (.A1(_1130_),
    .A2(net61),
    .ZN(_1142_));
 OR3_X1 _3481_ (.A1(_1084_),
    .A2(_1141_),
    .A3(_1142_),
    .ZN(_1143_));
 AOI221_X1 _3482_ (.A(_1134_),
    .B1(_1135_),
    .B2(_1143_),
    .C1(_0611_),
    .C2(_1120_),
    .ZN(net276));
 NOR3_X1 _3483_ (.A1(_1121_),
    .A2(net134),
    .A3(_1051_),
    .ZN(_1144_));
 AOI21_X1 _3484_ (.A(_1106_),
    .B1(_0343_),
    .B2(_1107_),
    .ZN(_1145_));
 AOI21_X1 _3485_ (.A(_1085_),
    .B1(net212),
    .B2(_1086_),
    .ZN(_1146_));
 NAND2_X1 _3486_ (.A1(_1110_),
    .A2(_0501_),
    .ZN(_1147_));
 OAI21_X1 _3487_ (.A(_1146_),
    .B1(_1147_),
    .B2(_1112_),
    .ZN(_1148_));
 AOI21_X1 _3488_ (.A(_1057_),
    .B1(_0910_),
    .B2(_1114_),
    .ZN(_1149_));
 AOI221_X2 _3489_ (.A(_1096_),
    .B1(_1148_),
    .B2(_1149_),
    .C1(_1456_),
    .C2(_1116_),
    .ZN(_1150_));
 NOR2_X1 _3490_ (.A1(_1130_),
    .A2(_1602_),
    .ZN(_1151_));
 OR3_X1 _3491_ (.A1(_1084_),
    .A2(_1150_),
    .A3(_1151_),
    .ZN(_1152_));
 AOI221_X1 _3492_ (.A(_1144_),
    .B1(_1145_),
    .B2(_1152_),
    .C1(_0617_),
    .C2(_1120_),
    .ZN(net277));
 NOR3_X1 _3493_ (.A1(_1121_),
    .A2(_0477_),
    .A3(_1051_),
    .ZN(_1153_));
 AOI21_X1 _3494_ (.A(_1106_),
    .B1(net99),
    .B2(_1107_),
    .ZN(_1154_));
 AOI21_X1 _3495_ (.A(_1085_),
    .B1(net213),
    .B2(_1086_),
    .ZN(_1155_));
 NAND2_X1 _3496_ (.A1(_1110_),
    .A2(net152),
    .ZN(_1156_));
 OAI21_X1 _3497_ (.A(_1155_),
    .B1(_1156_),
    .B2(_1112_),
    .ZN(_1157_));
 INV_X1 _3498_ (.A(net248),
    .ZN(_1158_));
 AOI21_X1 _3499_ (.A(_1057_),
    .B1(_1158_),
    .B2(_1114_),
    .ZN(_1159_));
 AOI221_X2 _3500_ (.A(_1096_),
    .B1(_1157_),
    .B2(_1159_),
    .C1(net28),
    .C2(_1116_),
    .ZN(_1160_));
 NOR2_X1 _3501_ (.A1(_1130_),
    .A2(net64),
    .ZN(_1161_));
 OR3_X1 _3502_ (.A1(_1084_),
    .A2(_1160_),
    .A3(_1161_),
    .ZN(_1162_));
 AOI221_X1 _3503_ (.A(_1153_),
    .B1(_1154_),
    .B2(_1162_),
    .C1(_0630_),
    .C2(_1120_),
    .ZN(net278));
 BUF_X2 _3504_ (.A(_0978_),
    .Z(_1163_));
 NOR3_X1 _3505_ (.A1(_1121_),
    .A2(_0481_),
    .A3(_1163_),
    .ZN(_1164_));
 AOI21_X1 _3506_ (.A(_1106_),
    .B1(_0351_),
    .B2(_1107_),
    .ZN(_1165_));
 AOI21_X1 _3507_ (.A(_1085_),
    .B1(_0788_),
    .B2(_1086_),
    .ZN(_1166_));
 NAND2_X1 _3508_ (.A1(_1110_),
    .A2(_0591_),
    .ZN(_1167_));
 OAI21_X1 _3509_ (.A(_1166_),
    .B1(_1167_),
    .B2(_1112_),
    .ZN(_1168_));
 CLKBUF_X3 _3510_ (.A(_1000_),
    .Z(_1169_));
 AOI21_X1 _3511_ (.A(_1169_),
    .B1(_0918_),
    .B2(_1114_),
    .ZN(_1170_));
 AOI221_X2 _3512_ (.A(_1096_),
    .B1(_1168_),
    .B2(_1170_),
    .C1(_1464_),
    .C2(_1116_),
    .ZN(_1171_));
 NOR2_X1 _3513_ (.A1(_1130_),
    .A2(net65),
    .ZN(_1172_));
 OR3_X1 _3514_ (.A1(_1084_),
    .A2(_1171_),
    .A3(_1172_),
    .ZN(_1173_));
 AOI221_X1 _3515_ (.A(_1164_),
    .B1(_1165_),
    .B2(_1173_),
    .C1(_0624_),
    .C2(_1120_),
    .ZN(net279));
 NOR3_X1 _3516_ (.A1(_1121_),
    .A2(_0486_),
    .A3(_1163_),
    .ZN(_1174_));
 AOI21_X1 _3517_ (.A(_1106_),
    .B1(_0356_),
    .B2(_1107_),
    .ZN(_1175_));
 AOI21_X1 _3518_ (.A(_1085_),
    .B1(_0793_),
    .B2(_1086_),
    .ZN(_1176_));
 NAND2_X1 _3519_ (.A1(_1110_),
    .A2(_0640_),
    .ZN(_1177_));
 OAI21_X1 _3520_ (.A(_1176_),
    .B1(_1177_),
    .B2(_1112_),
    .ZN(_1178_));
 AOI21_X1 _3521_ (.A(_1169_),
    .B1(_0928_),
    .B2(_1114_),
    .ZN(_1179_));
 AOI221_X2 _3522_ (.A(_1096_),
    .B1(_1178_),
    .B2(_1179_),
    .C1(_1473_),
    .C2(_1116_),
    .ZN(_1180_));
 NOR2_X1 _3523_ (.A1(_1130_),
    .A2(_1619_),
    .ZN(_1181_));
 OR3_X1 _3524_ (.A1(_1084_),
    .A2(_1180_),
    .A3(_1181_),
    .ZN(_1182_));
 INV_X1 _3525_ (.A(_0629_),
    .ZN(_1183_));
 AOI221_X1 _3526_ (.A(_1174_),
    .B1(_1175_),
    .B2(_1182_),
    .C1(_1183_),
    .C2(_1120_),
    .ZN(net280));
 NOR3_X1 _3527_ (.A1(_1121_),
    .A2(net138),
    .A3(_1163_),
    .ZN(_1184_));
 AOI21_X1 _3528_ (.A(_1106_),
    .B1(_0359_),
    .B2(_1107_),
    .ZN(_1185_));
 AOI21_X1 _3529_ (.A(_1085_),
    .B1(_0797_),
    .B2(_1086_),
    .ZN(_1186_));
 NAND2_X1 _3530_ (.A1(_1110_),
    .A2(_0664_),
    .ZN(_1187_));
 OAI21_X1 _3531_ (.A(_1186_),
    .B1(_1187_),
    .B2(_1112_),
    .ZN(_1188_));
 AOI21_X1 _3532_ (.A(_1169_),
    .B1(_0925_),
    .B2(_1114_),
    .ZN(_1189_));
 AOI221_X2 _3533_ (.A(_1096_),
    .B1(_1188_),
    .B2(_1189_),
    .C1(_1479_),
    .C2(_1116_),
    .ZN(_1190_));
 NOR2_X1 _3534_ (.A1(_1130_),
    .A2(net67),
    .ZN(_1191_));
 OR3_X1 _3535_ (.A1(_1084_),
    .A2(_1190_),
    .A3(_1191_),
    .ZN(_1192_));
 INV_X1 _3536_ (.A(_0636_),
    .ZN(_1193_));
 AOI221_X1 _3537_ (.A(_1184_),
    .B1(_1185_),
    .B2(_1192_),
    .C1(_1193_),
    .C2(_1120_),
    .ZN(net281));
 NOR3_X1 _3538_ (.A1(_1121_),
    .A2(net139),
    .A3(_1163_),
    .ZN(_1194_));
 AOI21_X2 _3539_ (.A(_1106_),
    .B1(net103),
    .B2(_1107_),
    .ZN(_1195_));
 BUF_X2 _3540_ (.A(_0984_),
    .Z(_1196_));
 CLKBUF_X3 _3541_ (.A(_0990_),
    .Z(_1197_));
 CLKBUF_X3 _3542_ (.A(_0992_),
    .Z(_1198_));
 AOI21_X1 _3543_ (.A(_1197_),
    .B1(net217),
    .B2(_1198_),
    .ZN(_1199_));
 NAND2_X1 _3544_ (.A1(_1110_),
    .A2(net182),
    .ZN(_1200_));
 OAI21_X1 _3545_ (.A(_1199_),
    .B1(_1200_),
    .B2(_1112_),
    .ZN(_1201_));
 AOI21_X1 _3546_ (.A(_1169_),
    .B1(_0939_),
    .B2(_1114_),
    .ZN(_1202_));
 AOI221_X2 _3547_ (.A(_1096_),
    .B1(_1201_),
    .B2(_1202_),
    .C1(net33),
    .C2(_1116_),
    .ZN(_1203_));
 NOR2_X1 _3548_ (.A1(_1130_),
    .A2(net68),
    .ZN(_1204_));
 OR3_X1 _3549_ (.A1(_1196_),
    .A2(_1203_),
    .A3(_1204_),
    .ZN(_1205_));
 INV_X1 _3550_ (.A(net175),
    .ZN(_1206_));
 AOI221_X2 _3551_ (.A(_1194_),
    .B1(_1195_),
    .B2(_1205_),
    .C1(_1206_),
    .C2(_1120_),
    .ZN(net282));
 NOR3_X1 _3552_ (.A1(_1121_),
    .A2(_0497_),
    .A3(_1163_),
    .ZN(_1207_));
 AOI21_X2 _3553_ (.A(_1106_),
    .B1(_0366_),
    .B2(_1107_),
    .ZN(_1208_));
 BUF_X4 _3554_ (.A(_0988_),
    .Z(_1209_));
 AOI21_X1 _3555_ (.A(_1197_),
    .B1(_0805_),
    .B2(_1198_),
    .ZN(_1210_));
 NAND2_X1 _3556_ (.A1(_1110_),
    .A2(net183),
    .ZN(_1211_));
 OAI21_X1 _3557_ (.A(_1210_),
    .B1(_1211_),
    .B2(_1112_),
    .ZN(_1212_));
 AOI21_X1 _3558_ (.A(_1169_),
    .B1(_0936_),
    .B2(_1114_),
    .ZN(_1213_));
 AOI221_X2 _3559_ (.A(_1209_),
    .B1(_1212_),
    .B2(_1213_),
    .C1(net34),
    .C2(_1116_),
    .ZN(_1214_));
 NOR2_X1 _3560_ (.A1(_1130_),
    .A2(_1629_),
    .ZN(_1215_));
 OR3_X1 _3561_ (.A1(_1196_),
    .A2(_1214_),
    .A3(_1215_),
    .ZN(_1216_));
 AOI221_X2 _3562_ (.A(_1207_),
    .B1(_1208_),
    .B2(_1216_),
    .C1(_0646_),
    .C2(_1120_),
    .ZN(net283));
 NOR3_X1 _3563_ (.A1(_1121_),
    .A2(_0505_),
    .A3(_1163_),
    .ZN(_1217_));
 BUF_X4 _3564_ (.A(_0982_),
    .Z(_1218_));
 BUF_X4 _3565_ (.A(_0984_),
    .Z(_1219_));
 AOI21_X2 _3566_ (.A(_1218_),
    .B1(_0370_),
    .B2(_1219_),
    .ZN(_1220_));
 AOI21_X1 _3567_ (.A(_1197_),
    .B1(net220),
    .B2(_1198_),
    .ZN(_1221_));
 BUF_X2 _3568_ (.A(_0995_),
    .Z(_1222_));
 NAND2_X1 _3569_ (.A1(_1222_),
    .A2(_0675_),
    .ZN(_1223_));
 CLKBUF_X3 _3570_ (.A(_0992_),
    .Z(_1224_));
 OAI21_X1 _3571_ (.A(_1221_),
    .B1(_1223_),
    .B2(_1224_),
    .ZN(_1225_));
 INV_X1 _3572_ (.A(_0941_),
    .ZN(_1226_));
 CLKBUF_X3 _3573_ (.A(_0990_),
    .Z(_1227_));
 AOI21_X1 _3574_ (.A(_1169_),
    .B1(_1226_),
    .B2(_1227_),
    .ZN(_1228_));
 BUF_X4 _3575_ (.A(_1001_),
    .Z(_1229_));
 AOI221_X2 _3576_ (.A(_1209_),
    .B1(_1225_),
    .B2(_1228_),
    .C1(_1494_),
    .C2(_1229_),
    .ZN(_1230_));
 NOR2_X1 _3577_ (.A1(_1130_),
    .A2(net70),
    .ZN(_1231_));
 OR3_X1 _3578_ (.A1(_1196_),
    .A2(_1230_),
    .A3(_1231_),
    .ZN(_1232_));
 INV_X1 _3579_ (.A(_0650_),
    .ZN(_1233_));
 BUF_X4 _3580_ (.A(_0979_),
    .Z(_1234_));
 AOI221_X2 _3581_ (.A(_1217_),
    .B1(_1220_),
    .B2(_1232_),
    .C1(_1233_),
    .C2(_1234_),
    .ZN(net284));
 CLKBUF_X3 _3582_ (.A(_0977_),
    .Z(_1235_));
 NOR3_X1 _3583_ (.A1(_1235_),
    .A2(_0510_),
    .A3(_1163_),
    .ZN(_1236_));
 AOI21_X1 _3584_ (.A(_1218_),
    .B1(net106),
    .B2(_1219_),
    .ZN(_1237_));
 AOI21_X1 _3585_ (.A(_1197_),
    .B1(net221),
    .B2(_1198_),
    .ZN(_1238_));
 NAND2_X1 _3586_ (.A1(_1222_),
    .A2(net185),
    .ZN(_1239_));
 OAI21_X1 _3587_ (.A(_1238_),
    .B1(_1239_),
    .B2(_1224_),
    .ZN(_1240_));
 INV_X1 _3588_ (.A(net256),
    .ZN(_1241_));
 AOI21_X1 _3589_ (.A(_1169_),
    .B1(_1241_),
    .B2(_1227_),
    .ZN(_1242_));
 AOI221_X2 _3590_ (.A(_1209_),
    .B1(_1240_),
    .B2(_1242_),
    .C1(_1499_),
    .C2(_1229_),
    .ZN(_1243_));
 CLKBUF_X3 _3591_ (.A(_1007_),
    .Z(_1244_));
 NOR2_X1 _3592_ (.A1(_1244_),
    .A2(net71),
    .ZN(_1245_));
 OR3_X1 _3593_ (.A1(_1196_),
    .A2(_1243_),
    .A3(_1245_),
    .ZN(_1246_));
 INV_X1 _3594_ (.A(net178),
    .ZN(_1247_));
 AOI221_X1 _3595_ (.A(_1236_),
    .B1(_1237_),
    .B2(_1246_),
    .C1(_1247_),
    .C2(_1234_),
    .ZN(net285));
 NOR3_X1 _3596_ (.A1(_1235_),
    .A2(_0393_),
    .A3(_1163_),
    .ZN(_1248_));
 AOI21_X2 _3597_ (.A(_1218_),
    .B1(_1656_),
    .B2(_1219_),
    .ZN(_1249_));
 AOI21_X1 _3598_ (.A(_1197_),
    .B1(net191),
    .B2(_1198_),
    .ZN(_1250_));
 NAND2_X1 _3599_ (.A1(_1222_),
    .A2(net186),
    .ZN(_1251_));
 OAI21_X1 _3600_ (.A(_1250_),
    .B1(_1251_),
    .B2(_1224_),
    .ZN(_1252_));
 AOI21_X1 _3601_ (.A(_1169_),
    .B1(_0831_),
    .B2(_1227_),
    .ZN(_1253_));
 AOI221_X2 _3602_ (.A(_1209_),
    .B1(_1252_),
    .B2(_1253_),
    .C1(_1363_),
    .C2(_1229_),
    .ZN(_1254_));
 NOR2_X1 _3603_ (.A1(_1244_),
    .A2(_1523_),
    .ZN(_1255_));
 OR3_X1 _3604_ (.A1(_1196_),
    .A2(_1254_),
    .A3(_1255_),
    .ZN(_1256_));
 AOI221_X2 _3605_ (.A(_1248_),
    .B1(_1249_),
    .B2(_1256_),
    .C1(_0528_),
    .C2(_1234_),
    .ZN(net286));
 NOR3_X1 _3606_ (.A1(_1235_),
    .A2(net144),
    .A3(_1163_),
    .ZN(_1257_));
 AOI21_X1 _3607_ (.A(_1218_),
    .B1(net108),
    .B2(_1219_),
    .ZN(_1258_));
 AOI21_X1 _3608_ (.A(_1197_),
    .B1(net222),
    .B2(_1198_),
    .ZN(_1259_));
 NAND2_X1 _3609_ (.A1(_1222_),
    .A2(net187),
    .ZN(_1260_));
 OAI21_X1 _3610_ (.A(_1259_),
    .B1(_1260_),
    .B2(_1224_),
    .ZN(_1261_));
 AOI21_X1 _3611_ (.A(_1169_),
    .B1(_0955_),
    .B2(_1227_),
    .ZN(_1262_));
 AOI221_X2 _3612_ (.A(_1209_),
    .B1(_1261_),
    .B2(_1262_),
    .C1(net37),
    .C2(_1229_),
    .ZN(_1263_));
 NOR2_X1 _3613_ (.A1(_1244_),
    .A2(net72),
    .ZN(_1264_));
 OR3_X1 _3614_ (.A1(_1196_),
    .A2(_1263_),
    .A3(_1264_),
    .ZN(_1265_));
 AOI221_X1 _3615_ (.A(_1257_),
    .B1(_1258_),
    .B2(_1265_),
    .C1(_0660_),
    .C2(_1234_),
    .ZN(net287));
 NOR3_X1 _3616_ (.A1(_1235_),
    .A2(net145),
    .A3(_1163_),
    .ZN(_1266_));
 AOI21_X1 _3617_ (.A(_1218_),
    .B1(net109),
    .B2(_1219_),
    .ZN(_1267_));
 HA_X1 _3618_ (.A(net189),
    .B(net190),
    .CO(_1925_),
    .S(_0001_));
 HA_X1 _3619_ (.A(net259),
    .B(net260),
    .CO(_1926_),
    .S(_0005_));
 HA_X1 _3620_ (.A(net39),
    .B(net40),
    .CO(_1927_),
    .S(_0007_));
 HA_X1 _3621_ (.A(net75),
    .B(net76),
    .CO(_1928_),
    .S(_0009_));
 HA_X1 _3622_ (.A(net110),
    .B(net111),
    .CO(_1929_),
    .S(_0011_));
 HA_X1 _3623_ (.A(net146),
    .B(net147),
    .CO(_1930_),
    .S(_0013_));
 HA_X1 _3624_ (.A(net8),
    .B(net119),
    .CO(_1931_),
    .S(_0015_));
 HA_X1 _3625_ (.A(net224),
    .B(net225),
    .CO(_1932_),
    .S(_0003_));
 DFF_X2 \counters[0]$_SDFFE_PP0P_  (.D(_0016_),
    .CK(clknet_leaf_1_clk),
    .Q(net8),
    .QN(_0014_));
 DFF_X1 \counters[100]$_SDFFE_PP0P_  (.D(_0017_),
    .CK(clknet_leaf_6_clk),
    .Q(net9),
    .QN(_1924_));
 DFF_X1 \counters[101]$_SDFFE_PP0P_  (.D(_0018_),
    .CK(clknet_leaf_6_clk),
    .Q(net10),
    .QN(_1923_));
 DFF_X1 \counters[102]$_SDFFE_PP0P_  (.D(_0019_),
    .CK(clknet_leaf_6_clk),
    .Q(net11),
    .QN(_1922_));
 DFF_X1 \counters[103]$_SDFFE_PP0P_  (.D(_0020_),
    .CK(clknet_leaf_6_clk),
    .Q(net12),
    .QN(_1921_));
 DFF_X1 \counters[104]$_SDFFE_PP0P_  (.D(_0021_),
    .CK(clknet_leaf_2_clk),
    .Q(net13),
    .QN(_1920_));
 DFF_X1 \counters[105]$_SDFFE_PP0P_  (.D(_0022_),
    .CK(clknet_leaf_1_clk),
    .Q(net14),
    .QN(_1919_));
 DFF_X2 \counters[106]$_SDFFE_PP0P_  (.D(_0023_),
    .CK(clknet_leaf_2_clk),
    .Q(net15),
    .QN(_1918_));
 DFF_X1 \counters[107]$_SDFFE_PP0P_  (.D(_0024_),
    .CK(clknet_leaf_2_clk),
    .Q(net16),
    .QN(_1917_));
 DFF_X1 \counters[108]$_SDFFE_PP0P_  (.D(_0025_),
    .CK(clknet_leaf_2_clk),
    .Q(net17),
    .QN(_1916_));
 DFF_X1 \counters[109]$_SDFFE_PP0P_  (.D(_0026_),
    .CK(clknet_leaf_5_clk),
    .Q(net18),
    .QN(_1915_));
 DFF_X2 \counters[10]$_SDFFE_PP0P_  (.D(_0027_),
    .CK(clknet_leaf_3_clk),
    .Q(net19),
    .QN(_1914_));
 DFF_X1 \counters[110]$_SDFFE_PP0P_  (.D(_0028_),
    .CK(clknet_leaf_2_clk),
    .Q(net20),
    .QN(_1913_));
 DFF_X2 \counters[111]$_SDFFE_PP0P_  (.D(_0029_),
    .CK(clknet_leaf_2_clk),
    .Q(net21),
    .QN(_1912_));
 DFF_X2 \counters[112]$_SDFFE_PP0P_  (.D(_0030_),
    .CK(clknet_leaf_3_clk),
    .Q(net22),
    .QN(_1911_));
 DFF_X1 \counters[113]$_SDFFE_PP0P_  (.D(_0031_),
    .CK(clknet_leaf_4_clk),
    .Q(net23),
    .QN(_1910_));
 DFF_X1 \counters[114]$_SDFFE_PP0P_  (.D(_0032_),
    .CK(clknet_leaf_3_clk),
    .Q(net24),
    .QN(_1909_));
 DFF_X1 \counters[115]$_SDFFE_PP0P_  (.D(_0033_),
    .CK(clknet_leaf_4_clk),
    .Q(net25),
    .QN(_1908_));
 DFF_X2 \counters[116]$_SDFFE_PP0P_  (.D(_0034_),
    .CK(clknet_leaf_4_clk),
    .Q(net26),
    .QN(_1907_));
 DFF_X1 \counters[117]$_SDFFE_PP0P_  (.D(_0035_),
    .CK(clknet_leaf_4_clk),
    .Q(net27),
    .QN(_1906_));
 DFF_X2 \counters[118]$_SDFFE_PP0P_  (.D(_0036_),
    .CK(clknet_leaf_4_clk),
    .Q(net28),
    .QN(_1905_));
 DFF_X1 \counters[119]$_SDFFE_PP0P_  (.D(_0037_),
    .CK(clknet_leaf_5_clk),
    .Q(net29),
    .QN(_1904_));
 DFF_X1 \counters[11]$_SDFFE_PP0P_  (.D(_0038_),
    .CK(clknet_leaf_3_clk),
    .Q(net30),
    .QN(_1903_));
 DFF_X1 \counters[120]$_SDFFE_PP0P_  (.D(_0039_),
    .CK(clknet_leaf_12_clk),
    .Q(net31),
    .QN(_1902_));
 DFF_X1 \counters[121]$_SDFFE_PP0P_  (.D(_0040_),
    .CK(clknet_leaf_4_clk),
    .Q(net32),
    .QN(_1901_));
 DFF_X2 \counters[122]$_SDFFE_PP0P_  (.D(_0041_),
    .CK(clknet_leaf_13_clk),
    .Q(net33),
    .QN(_1900_));
 DFF_X2 \counters[123]$_SDFFE_PP0P_  (.D(_0042_),
    .CK(clknet_leaf_13_clk),
    .Q(net34),
    .QN(_1899_));
 DFF_X1 \counters[124]$_SDFFE_PP0P_  (.D(_0043_),
    .CK(clknet_leaf_5_clk),
    .Q(net35),
    .QN(_1898_));
 DFF_X1 \counters[125]$_SDFFE_PP0P_  (.D(_0044_),
    .CK(clknet_leaf_12_clk),
    .Q(net36),
    .QN(_1897_));
 DFF_X2 \counters[126]$_SDFFE_PP0P_  (.D(_0045_),
    .CK(clknet_leaf_12_clk),
    .Q(net37),
    .QN(_1896_));
 DFF_X2 \counters[127]$_SDFFE_PP0P_  (.D(_0046_),
    .CK(clknet_leaf_12_clk),
    .Q(net38),
    .QN(_1895_));
 DFF_X2 \counters[128]$_SDFFE_PP0P_  (.D(_0047_),
    .CK(clknet_leaf_13_clk),
    .Q(net39),
    .QN(_0006_));
 DFF_X2 \counters[129]$_SDFFE_PP0P_  (.D(_0048_),
    .CK(clknet_leaf_13_clk),
    .Q(net40),
    .QN(_1894_));
 DFF_X1 \counters[12]$_SDFFE_PP0P_  (.D(_0049_),
    .CK(clknet_leaf_36_clk),
    .Q(net41),
    .QN(_1893_));
 DFF_X1 \counters[130]$_SDFFE_PP0P_  (.D(_0050_),
    .CK(clknet_leaf_13_clk),
    .Q(net42),
    .QN(_1892_));
 DFF_X2 \counters[131]$_SDFFE_PP0P_  (.D(_0051_),
    .CK(clknet_leaf_14_clk),
    .Q(net43),
    .QN(_1891_));
 DFF_X2 \counters[132]$_SDFFE_PP0P_  (.D(_0052_),
    .CK(clknet_leaf_13_clk),
    .Q(net44),
    .QN(_1890_));
 DFF_X2 \counters[133]$_SDFFE_PP0P_  (.D(_0053_),
    .CK(clknet_leaf_23_clk),
    .Q(net45),
    .QN(_1889_));
 DFF_X1 \counters[134]$_SDFFE_PP0P_  (.D(_0054_),
    .CK(clknet_leaf_23_clk),
    .Q(net46),
    .QN(_1888_));
 DFF_X1 \counters[135]$_SDFFE_PP0P_  (.D(_0055_),
    .CK(clknet_leaf_34_clk),
    .Q(net47),
    .QN(_1887_));
 DFF_X1 \counters[136]$_SDFFE_PP0P_  (.D(_0056_),
    .CK(clknet_leaf_34_clk),
    .Q(net48),
    .QN(_1886_));
 DFF_X1 \counters[137]$_SDFFE_PP0P_  (.D(_0057_),
    .CK(clknet_leaf_4_clk),
    .Q(net49),
    .QN(_1885_));
 DFF_X2 \counters[138]$_SDFFE_PP0P_  (.D(_0058_),
    .CK(clknet_leaf_34_clk),
    .Q(net50),
    .QN(_1884_));
 DFF_X1 \counters[139]$_SDFFE_PP0P_  (.D(_0059_),
    .CK(clknet_leaf_23_clk),
    .Q(net51),
    .QN(_1883_));
 DFF_X1 \counters[13]$_SDFFE_PP0P_  (.D(_0060_),
    .CK(clknet_leaf_32_clk),
    .Q(net52),
    .QN(_1882_));
 DFF_X1 \counters[140]$_SDFFE_PP0P_  (.D(_0061_),
    .CK(clknet_leaf_24_clk),
    .Q(net53),
    .QN(_1881_));
 DFF_X1 \counters[141]$_SDFFE_PP0P_  (.D(_0062_),
    .CK(clknet_leaf_34_clk),
    .Q(net54),
    .QN(_1880_));
 DFF_X2 \counters[142]$_SDFFE_PP0P_  (.D(_0063_),
    .CK(clknet_leaf_33_clk),
    .Q(net55),
    .QN(_1879_));
 DFF_X1 \counters[143]$_SDFFE_PP0P_  (.D(_0064_),
    .CK(clknet_leaf_33_clk),
    .Q(net56),
    .QN(_1878_));
 DFF_X1 \counters[144]$_SDFFE_PP0P_  (.D(_0065_),
    .CK(clknet_leaf_33_clk),
    .Q(net57),
    .QN(_1877_));
 DFF_X2 \counters[145]$_SDFFE_PP0P_  (.D(_0066_),
    .CK(clknet_leaf_24_clk),
    .Q(net58),
    .QN(_1876_));
 DFF_X2 \counters[146]$_SDFFE_PP0P_  (.D(_0067_),
    .CK(clknet_leaf_24_clk),
    .Q(net59),
    .QN(_1875_));
 DFF_X2 \counters[147]$_SDFFE_PP0P_  (.D(_0068_),
    .CK(clknet_leaf_33_clk),
    .Q(net60),
    .QN(_1874_));
 DFF_X2 \counters[148]$_SDFFE_PP0P_  (.D(_0069_),
    .CK(clknet_leaf_33_clk),
    .Q(net61),
    .QN(_1873_));
 DFF_X1 \counters[149]$_SDFFE_PP0P_  (.D(_0070_),
    .CK(clknet_leaf_23_clk),
    .Q(net62),
    .QN(_1872_));
 DFF_X1 \counters[14]$_SDFFE_PP0P_  (.D(_0071_),
    .CK(clknet_leaf_32_clk),
    .Q(net63),
    .QN(_1871_));
 DFF_X2 \counters[150]$_SDFFE_PP0P_  (.D(_0072_),
    .CK(clknet_leaf_23_clk),
    .Q(net64),
    .QN(_1870_));
 DFF_X2 \counters[151]$_SDFFE_PP0P_  (.D(_0073_),
    .CK(clknet_leaf_14_clk),
    .Q(net65),
    .QN(_1869_));
 DFF_X1 \counters[152]$_SDFFE_PP0P_  (.D(_0074_),
    .CK(clknet_leaf_15_clk),
    .Q(net66),
    .QN(_1868_));
 DFF_X2 \counters[153]$_SDFFE_PP0P_  (.D(_0075_),
    .CK(clknet_leaf_15_clk),
    .Q(net67),
    .QN(_1867_));
 DFF_X2 \counters[154]$_SDFFE_PP0P_  (.D(_0076_),
    .CK(clknet_leaf_15_clk),
    .Q(net68),
    .QN(_1866_));
 DFF_X1 \counters[155]$_SDFFE_PP0P_  (.D(_0077_),
    .CK(clknet_leaf_15_clk),
    .Q(net69),
    .QN(_1865_));
 DFF_X2 \counters[156]$_SDFFE_PP0P_  (.D(_0078_),
    .CK(clknet_leaf_15_clk),
    .Q(net70),
    .QN(_1864_));
 DFF_X2 \counters[157]$_SDFFE_PP0P_  (.D(_0079_),
    .CK(clknet_leaf_15_clk),
    .Q(net71),
    .QN(_1863_));
 DFF_X1 \counters[158]$_SDFFE_PP0P_  (.D(_0080_),
    .CK(clknet_leaf_11_clk),
    .Q(net72),
    .QN(_1862_));
 DFF_X1 \counters[159]$_SDFFE_PP0P_  (.D(_0081_),
    .CK(clknet_leaf_11_clk),
    .Q(net73),
    .QN(_1861_));
 DFF_X2 \counters[15]$_SDFFE_PP0P_  (.D(_0082_),
    .CK(clknet_leaf_31_clk),
    .Q(net74),
    .QN(_1860_));
 DFF_X2 \counters[160]$_SDFFE_PP0P_  (.D(_0083_),
    .CK(clknet_leaf_24_clk),
    .Q(net75),
    .QN(_0008_));
 DFF_X2 \counters[161]$_SDFFE_PP0P_  (.D(_0084_),
    .CK(clknet_leaf_27_clk),
    .Q(net76),
    .QN(_1859_));
 DFF_X1 \counters[162]$_SDFFE_PP0P_  (.D(_0085_),
    .CK(clknet_leaf_30_clk),
    .Q(net77),
    .QN(_1858_));
 DFF_X1 \counters[163]$_SDFFE_PP0P_  (.D(_0086_),
    .CK(clknet_leaf_31_clk),
    .Q(net78),
    .QN(_1857_));
 DFF_X2 \counters[164]$_SDFFE_PP0P_  (.D(_0087_),
    .CK(clknet_leaf_32_clk),
    .Q(net79),
    .QN(_1856_));
 DFF_X2 \counters[165]$_SDFFE_PP0P_  (.D(_0088_),
    .CK(clknet_leaf_30_clk),
    .Q(net80),
    .QN(_1855_));
 DFF_X1 \counters[166]$_SDFFE_PP0P_  (.D(_0089_),
    .CK(clknet_leaf_30_clk),
    .Q(net81),
    .QN(_1854_));
 DFF_X1 \counters[167]$_SDFFE_PP0P_  (.D(_0090_),
    .CK(clknet_leaf_30_clk),
    .Q(net82),
    .QN(_1853_));
 DFF_X2 \counters[168]$_SDFFE_PP0P_  (.D(_0091_),
    .CK(clknet_leaf_30_clk),
    .Q(net83),
    .QN(_1852_));
 DFF_X2 \counters[169]$_SDFFE_PP0P_  (.D(_0092_),
    .CK(clknet_leaf_30_clk),
    .Q(net84),
    .QN(_1851_));
 DFF_X1 \counters[16]$_SDFFE_PP0P_  (.D(_0093_),
    .CK(clknet_leaf_31_clk),
    .Q(net85),
    .QN(_1850_));
 DFF_X1 \counters[170]$_SDFFE_PP0P_  (.D(_0094_),
    .CK(clknet_leaf_29_clk),
    .Q(net86),
    .QN(_1849_));
 DFF_X2 \counters[171]$_SDFFE_PP0P_  (.D(_0095_),
    .CK(clknet_leaf_29_clk),
    .Q(net87),
    .QN(_1848_));
 DFF_X1 \counters[172]$_SDFFE_PP0P_  (.D(_0096_),
    .CK(clknet_leaf_29_clk),
    .Q(net88),
    .QN(_1847_));
 DFF_X1 \counters[173]$_SDFFE_PP0P_  (.D(_0097_),
    .CK(clknet_leaf_29_clk),
    .Q(net89),
    .QN(_1846_));
 DFF_X2 \counters[174]$_SDFFE_PP0P_  (.D(_0098_),
    .CK(clknet_leaf_29_clk),
    .Q(net90),
    .QN(_1845_));
 DFF_X1 \counters[175]$_SDFFE_PP0P_  (.D(_0099_),
    .CK(clknet_leaf_29_clk),
    .Q(net91),
    .QN(_1844_));
 DFF_X1 \counters[176]$_SDFFE_PP0P_  (.D(_0100_),
    .CK(clknet_leaf_30_clk),
    .Q(net92),
    .QN(_1843_));
 DFF_X1 \counters[177]$_SDFFE_PP0P_  (.D(_0101_),
    .CK(clknet_leaf_28_clk),
    .Q(net93),
    .QN(_1842_));
 DFF_X1 \counters[178]$_SDFFE_PP0P_  (.D(_0102_),
    .CK(clknet_leaf_28_clk),
    .Q(net94),
    .QN(_1841_));
 DFF_X1 \counters[179]$_SDFFE_PP0P_  (.D(_0103_),
    .CK(clknet_leaf_27_clk),
    .Q(net95),
    .QN(_1840_));
 DFF_X2 \counters[17]$_SDFFE_PP0P_  (.D(_0104_),
    .CK(clknet_leaf_32_clk),
    .Q(net96),
    .QN(_1839_));
 DFF_X2 \counters[180]$_SDFFE_PP0P_  (.D(_0105_),
    .CK(clknet_leaf_27_clk),
    .Q(net97),
    .QN(_1838_));
 DFF_X1 \counters[181]$_SDFFE_PP0P_  (.D(_0106_),
    .CK(clknet_leaf_26_clk),
    .Q(net98),
    .QN(_1837_));
 DFF_X1 \counters[182]$_SDFFE_PP0P_  (.D(_0107_),
    .CK(clknet_leaf_27_clk),
    .Q(net99),
    .QN(_1836_));
 DFF_X1 \counters[183]$_SDFFE_PP0P_  (.D(_0108_),
    .CK(clknet_leaf_28_clk),
    .Q(net100),
    .QN(_1835_));
 DFF_X1 \counters[184]$_SDFFE_PP0P_  (.D(_0109_),
    .CK(clknet_leaf_28_clk),
    .Q(net101),
    .QN(_1834_));
 DFF_X1 \counters[185]$_SDFFE_PP0P_  (.D(_0110_),
    .CK(clknet_leaf_28_clk),
    .Q(net102),
    .QN(_1833_));
 DFF_X2 \counters[186]$_SDFFE_PP0P_  (.D(_0111_),
    .CK(clknet_leaf_28_clk),
    .Q(net103),
    .QN(_1832_));
 DFF_X1 \counters[187]$_SDFFE_PP0P_  (.D(_0112_),
    .CK(clknet_leaf_26_clk),
    .Q(net104),
    .QN(_1831_));
 DFF_X1 \counters[188]$_SDFFE_PP0P_  (.D(_0113_),
    .CK(clknet_leaf_28_clk),
    .Q(net105),
    .QN(_1830_));
 DFF_X1 \counters[189]$_SDFFE_PP0P_  (.D(_0114_),
    .CK(clknet_leaf_26_clk),
    .Q(net106),
    .QN(_1829_));
 DFF_X1 \counters[18]$_SDFFE_PP0P_  (.D(_0115_),
    .CK(clknet_leaf_32_clk),
    .Q(net107),
    .QN(_1828_));
 DFF_X1 \counters[190]$_SDFFE_PP0P_  (.D(_0116_),
    .CK(clknet_leaf_27_clk),
    .Q(net108),
    .QN(_1827_));
 DFF_X1 \counters[191]$_SDFFE_PP0P_  (.D(_0117_),
    .CK(clknet_leaf_26_clk),
    .Q(net109),
    .QN(_1826_));
 DFF_X2 \counters[192]$_SDFFE_PP0P_  (.D(_0118_),
    .CK(clknet_leaf_14_clk),
    .Q(net110),
    .QN(_0010_));
 DFF_X2 \counters[193]$_SDFFE_PP0P_  (.D(_0119_),
    .CK(clknet_leaf_20_clk),
    .Q(net111),
    .QN(_1825_));
 DFF_X1 \counters[194]$_SDFFE_PP0P_  (.D(_0120_),
    .CK(clknet_leaf_14_clk),
    .Q(net112),
    .QN(_1824_));
 DFF_X2 \counters[195]$_SDFFE_PP0P_  (.D(_0121_),
    .CK(clknet_leaf_14_clk),
    .Q(net113),
    .QN(_1823_));
 DFF_X1 \counters[196]$_SDFFE_PP0P_  (.D(_0122_),
    .CK(clknet_leaf_16_clk),
    .Q(net114),
    .QN(_1822_));
 DFF_X2 \counters[197]$_SDFFE_PP0P_  (.D(_0123_),
    .CK(clknet_leaf_16_clk),
    .Q(net115),
    .QN(_1821_));
 DFF_X2 \counters[198]$_SDFFE_PP0P_  (.D(_0124_),
    .CK(clknet_leaf_16_clk),
    .Q(net116),
    .QN(_1820_));
 DFF_X1 \counters[199]$_SDFFE_PP0P_  (.D(_0125_),
    .CK(clknet_leaf_16_clk),
    .Q(net117),
    .QN(_1819_));
 DFF_X2 \counters[19]$_SDFFE_PP0P_  (.D(_0126_),
    .CK(clknet_leaf_33_clk),
    .Q(net118),
    .QN(_1818_));
 DFF_X2 \counters[1]$_SDFFE_PP0P_  (.D(_0127_),
    .CK(clknet_leaf_1_clk),
    .Q(net119),
    .QN(_1817_));
 DFF_X1 \counters[200]$_SDFFE_PP0P_  (.D(_0128_),
    .CK(clknet_leaf_16_clk),
    .Q(net120),
    .QN(_1816_));
 DFF_X2 \counters[201]$_SDFFE_PP0P_  (.D(_0129_),
    .CK(clknet_leaf_16_clk),
    .Q(net121),
    .QN(_1815_));
 DFF_X2 \counters[202]$_SDFFE_PP0P_  (.D(_0130_),
    .CK(clknet_leaf_16_clk),
    .Q(net122),
    .QN(_1814_));
 DFF_X1 \counters[203]$_SDFFE_PP0P_  (.D(_0131_),
    .CK(clknet_leaf_16_clk),
    .Q(net123),
    .QN(_1813_));
 DFF_X2 \counters[204]$_SDFFE_PP0P_  (.D(_0132_),
    .CK(clknet_leaf_17_clk),
    .Q(net124),
    .QN(_1812_));
 DFF_X2 \counters[205]$_SDFFE_PP0P_  (.D(_0133_),
    .CK(clknet_leaf_17_clk),
    .Q(net125),
    .QN(_1811_));
 DFF_X2 \counters[206]$_SDFFE_PP0P_  (.D(_0134_),
    .CK(clknet_leaf_17_clk),
    .Q(net126),
    .QN(_1810_));
 DFF_X2 \counters[207]$_SDFFE_PP0P_  (.D(_0135_),
    .CK(clknet_leaf_19_clk),
    .Q(net127),
    .QN(_1809_));
 DFF_X2 \counters[208]$_SDFFE_PP0P_  (.D(_0136_),
    .CK(clknet_leaf_19_clk),
    .Q(net128),
    .QN(_1808_));
 DFF_X2 \counters[209]$_SDFFE_PP0P_  (.D(_0137_),
    .CK(clknet_leaf_17_clk),
    .Q(net129),
    .QN(_1807_));
 DFF_X2 \counters[20]$_SDFFE_PP0P_  (.D(_0138_),
    .CK(clknet_leaf_33_clk),
    .Q(net130),
    .QN(_1806_));
 DFF_X1 \counters[210]$_SDFFE_PP0P_  (.D(_0139_),
    .CK(clknet_leaf_17_clk),
    .Q(net131),
    .QN(_1805_));
 DFF_X1 \counters[211]$_SDFFE_PP0P_  (.D(_0140_),
    .CK(clknet_leaf_17_clk),
    .Q(net132),
    .QN(_1804_));
 DFF_X1 \counters[212]$_SDFFE_PP0P_  (.D(_0141_),
    .CK(clknet_leaf_17_clk),
    .Q(net133),
    .QN(_1803_));
 DFF_X2 \counters[213]$_SDFFE_PP0P_  (.D(_0142_),
    .CK(clknet_leaf_18_clk),
    .Q(net134),
    .QN(_1802_));
 DFF_X1 \counters[214]$_SDFFE_PP0P_  (.D(_0143_),
    .CK(clknet_leaf_18_clk),
    .Q(net135),
    .QN(_1801_));
 DFF_X1 \counters[215]$_SDFFE_PP0P_  (.D(_0144_),
    .CK(clknet_leaf_18_clk),
    .Q(net136),
    .QN(_1800_));
 DFF_X1 \counters[216]$_SDFFE_PP0P_  (.D(_0145_),
    .CK(clknet_leaf_18_clk),
    .Q(net137),
    .QN(_1799_));
 DFF_X2 \counters[217]$_SDFFE_PP0P_  (.D(_0146_),
    .CK(clknet_leaf_18_clk),
    .Q(net138),
    .QN(_1798_));
 DFF_X2 \counters[218]$_SDFFE_PP0P_  (.D(_0147_),
    .CK(clknet_leaf_19_clk),
    .Q(net139),
    .QN(_1797_));
 DFF_X1 \counters[219]$_SDFFE_PP0P_  (.D(_0148_),
    .CK(clknet_leaf_18_clk),
    .Q(net140),
    .QN(_1796_));
 DFF_X1 \counters[21]$_SDFFE_PP0P_  (.D(_0149_),
    .CK(clknet_leaf_32_clk),
    .Q(net141),
    .QN(_1795_));
 DFF_X1 \counters[220]$_SDFFE_PP0P_  (.D(_0150_),
    .CK(clknet_leaf_18_clk),
    .Q(net142),
    .QN(_1794_));
 DFF_X1 \counters[221]$_SDFFE_PP0P_  (.D(_0151_),
    .CK(clknet_leaf_19_clk),
    .Q(net143),
    .QN(_1793_));
 DFF_X1 \counters[222]$_SDFFE_PP0P_  (.D(_0152_),
    .CK(clknet_leaf_19_clk),
    .Q(net144),
    .QN(_1792_));
 DFF_X1 \counters[223]$_SDFFE_PP0P_  (.D(_0153_),
    .CK(clknet_leaf_19_clk),
    .Q(net145),
    .QN(_1791_));
 DFF_X2 \counters[224]$_SDFFE_PP0P_  (.D(_0154_),
    .CK(clknet_leaf_22_clk),
    .Q(net146),
    .QN(_0012_));
 DFF_X2 \counters[225]$_SDFFE_PP0P_  (.D(_0155_),
    .CK(clknet_leaf_22_clk),
    .Q(net147),
    .QN(_1790_));
 DFF_X2 \counters[226]$_SDFFE_PP0P_  (.D(_0156_),
    .CK(clknet_leaf_22_clk),
    .Q(net148),
    .QN(_1789_));
 DFF_X1 \counters[227]$_SDFFE_PP0P_  (.D(_0157_),
    .CK(clknet_leaf_14_clk),
    .Q(net149),
    .QN(_1788_));
 DFF_X1 \counters[228]$_SDFFE_PP0P_  (.D(_0158_),
    .CK(clknet_leaf_21_clk),
    .Q(net150),
    .QN(_1787_));
 DFF_X1 \counters[229]$_SDFFE_PP0P_  (.D(_0159_),
    .CK(clknet_leaf_22_clk),
    .Q(net151),
    .QN(_1786_));
 DFF_X2 \counters[22]$_SDFFE_PP0P_  (.D(_0160_),
    .CK(clknet_leaf_33_clk),
    .Q(net152),
    .QN(_1785_));
 DFF_X2 \counters[230]$_SDFFE_PP0P_  (.D(_0161_),
    .CK(clknet_leaf_22_clk),
    .Q(net153),
    .QN(_1784_));
 DFF_X2 \counters[231]$_SDFFE_PP0P_  (.D(_0162_),
    .CK(clknet_leaf_23_clk),
    .Q(net154),
    .QN(_1783_));
 DFF_X1 \counters[232]$_SDFFE_PP0P_  (.D(_0163_),
    .CK(clknet_leaf_21_clk),
    .Q(net155),
    .QN(_1782_));
 DFF_X2 \counters[233]$_SDFFE_PP0P_  (.D(_0164_),
    .CK(clknet_leaf_23_clk),
    .Q(net156),
    .QN(_1781_));
 DFF_X1 \counters[234]$_SDFFE_PP0P_  (.D(_0165_),
    .CK(clknet_leaf_21_clk),
    .Q(net157),
    .QN(_1780_));
 DFF_X1 \counters[235]$_SDFFE_PP0P_  (.D(_0166_),
    .CK(clknet_leaf_25_clk),
    .Q(net158),
    .QN(_1779_));
 DFF_X2 \counters[236]$_SDFFE_PP0P_  (.D(_0167_),
    .CK(clknet_leaf_24_clk),
    .Q(net159),
    .QN(_1778_));
 DFF_X1 \counters[237]$_SDFFE_PP0P_  (.D(_0168_),
    .CK(clknet_leaf_25_clk),
    .Q(net160),
    .QN(_1777_));
 DFF_X2 \counters[238]$_SDFFE_PP0P_  (.D(_0169_),
    .CK(clknet_leaf_24_clk),
    .Q(net161),
    .QN(_1776_));
 DFF_X2 \counters[239]$_SDFFE_PP0P_  (.D(_0170_),
    .CK(clknet_leaf_27_clk),
    .Q(net162),
    .QN(_1775_));
 DFF_X1 \counters[23]$_SDFFE_PP0P_  (.D(_0171_),
    .CK(clknet_leaf_34_clk),
    .Q(net163),
    .QN(_1774_));
 DFF_X2 \counters[240]$_SDFFE_PP0P_  (.D(_0172_),
    .CK(clknet_leaf_26_clk),
    .Q(net164),
    .QN(_1773_));
 DFF_X1 \counters[241]$_SDFFE_PP0P_  (.D(_0173_),
    .CK(clknet_leaf_26_clk),
    .Q(net165),
    .QN(_1772_));
 DFF_X2 \counters[242]$_SDFFE_PP0P_  (.D(_0174_),
    .CK(clknet_leaf_26_clk),
    .Q(net166),
    .QN(_1771_));
 DFF_X1 \counters[243]$_SDFFE_PP0P_  (.D(_0175_),
    .CK(clknet_leaf_25_clk),
    .Q(net167),
    .QN(_1770_));
 DFF_X1 \counters[244]$_SDFFE_PP0P_  (.D(_0176_),
    .CK(clknet_leaf_25_clk),
    .Q(net168),
    .QN(_1769_));
 DFF_X2 \counters[245]$_SDFFE_PP0P_  (.D(_0177_),
    .CK(clknet_leaf_25_clk),
    .Q(net169),
    .QN(_1768_));
 DFF_X1 \counters[246]$_SDFFE_PP0P_  (.D(_0178_),
    .CK(clknet_leaf_25_clk),
    .Q(net170),
    .QN(_1767_));
 DFF_X1 \counters[247]$_SDFFE_PP0P_  (.D(_0179_),
    .CK(clknet_leaf_21_clk),
    .Q(net171),
    .QN(_1766_));
 DFF_X1 \counters[248]$_SDFFE_PP0P_  (.D(_0180_),
    .CK(clknet_leaf_21_clk),
    .Q(net172),
    .QN(_1765_));
 DFF_X1 \counters[249]$_SDFFE_PP0P_  (.D(_0181_),
    .CK(clknet_leaf_21_clk),
    .Q(net173),
    .QN(_1764_));
 DFF_X1 \counters[24]$_SDFFE_PP0P_  (.D(_0182_),
    .CK(clknet_leaf_35_clk),
    .Q(net174),
    .QN(_1763_));
 DFF_X1 \counters[250]$_SDFFE_PP0P_  (.D(_0183_),
    .CK(clknet_leaf_21_clk),
    .Q(net175),
    .QN(_1762_));
 DFF_X2 \counters[251]$_SDFFE_PP0P_  (.D(_0184_),
    .CK(clknet_leaf_20_clk),
    .Q(net176),
    .QN(_1761_));
 DFF_X1 \counters[252]$_SDFFE_PP0P_  (.D(_0185_),
    .CK(clknet_leaf_20_clk),
    .Q(net177),
    .QN(_1760_));
 DFF_X1 \counters[253]$_SDFFE_PP0P_  (.D(_0186_),
    .CK(clknet_leaf_20_clk),
    .Q(net178),
    .QN(_1759_));
 DFF_X1 \counters[254]$_SDFFE_PP0P_  (.D(_0187_),
    .CK(clknet_leaf_20_clk),
    .Q(net179),
    .QN(_1758_));
 DFF_X1 \counters[255]$_SDFFE_PP0P_  (.D(_0188_),
    .CK(clknet_leaf_20_clk),
    .Q(net180),
    .QN(_1757_));
 DFF_X1 \counters[25]$_SDFFE_PP0P_  (.D(_0189_),
    .CK(clknet_leaf_35_clk),
    .Q(net181),
    .QN(_1756_));
 DFF_X2 \counters[26]$_SDFFE_PP0P_  (.D(_0190_),
    .CK(clknet_leaf_35_clk),
    .Q(net182),
    .QN(_1755_));
 DFF_X2 \counters[27]$_SDFFE_PP0P_  (.D(_0191_),
    .CK(clknet_leaf_35_clk),
    .Q(net183),
    .QN(_1754_));
 DFF_X1 \counters[28]$_SDFFE_PP0P_  (.D(_0192_),
    .CK(clknet_leaf_35_clk),
    .Q(net184),
    .QN(_1753_));
 DFF_X2 \counters[29]$_SDFFE_PP0P_  (.D(_0193_),
    .CK(clknet_leaf_3_clk),
    .Q(net185),
    .QN(_1752_));
 DFF_X2 \counters[2]$_SDFFE_PP0P_  (.D(_0194_),
    .CK(clknet_leaf_0_clk),
    .Q(net186),
    .QN(_1751_));
 DFF_X1 \counters[30]$_SDFFE_PP0P_  (.D(_0195_),
    .CK(clknet_leaf_35_clk),
    .Q(net187),
    .QN(_1750_));
 DFF_X1 \counters[31]$_SDFFE_PP0P_  (.D(_0196_),
    .CK(clknet_leaf_37_clk),
    .Q(net188),
    .QN(_1749_));
 DFF_X2 \counters[32]$_SDFFE_PP0P_  (.D(_0197_),
    .CK(clknet_leaf_0_clk),
    .Q(net189),
    .QN(_0000_));
 DFF_X2 \counters[33]$_SDFFE_PP0P_  (.D(_0198_),
    .CK(clknet_leaf_3_clk),
    .Q(net190),
    .QN(_1748_));
 DFF_X2 \counters[34]$_SDFFE_PP0P_  (.D(_0199_),
    .CK(clknet_leaf_0_clk),
    .Q(net191),
    .QN(_1747_));
 DFF_X1 \counters[35]$_SDFFE_PP0P_  (.D(_0200_),
    .CK(clknet_leaf_39_clk),
    .Q(net192),
    .QN(_1746_));
 DFF_X1 \counters[36]$_SDFFE_PP0P_  (.D(_0201_),
    .CK(clknet_leaf_39_clk),
    .Q(net193),
    .QN(_1745_));
 DFF_X1 \counters[37]$_SDFFE_PP0P_  (.D(_0202_),
    .CK(clknet_leaf_39_clk),
    .Q(net194),
    .QN(_1744_));
 DFF_X1 \counters[38]$_SDFFE_PP0P_  (.D(_0203_),
    .CK(clknet_leaf_39_clk),
    .Q(net195),
    .QN(_1743_));
 DFF_X1 \counters[39]$_SDFFE_PP0P_  (.D(_0204_),
    .CK(clknet_leaf_38_clk),
    .Q(net196),
    .QN(_1742_));
 DFF_X1 \counters[3]$_SDFFE_PP0P_  (.D(_0205_),
    .CK(clknet_leaf_39_clk),
    .Q(net197),
    .QN(_1741_));
 DFF_X1 \counters[40]$_SDFFE_PP0P_  (.D(_0206_),
    .CK(clknet_leaf_39_clk),
    .Q(net198),
    .QN(_1740_));
 DFF_X1 \counters[41]$_SDFFE_PP0P_  (.D(_0207_),
    .CK(clknet_leaf_38_clk),
    .Q(net199),
    .QN(_1739_));
 DFF_X2 \counters[42]$_SDFFE_PP0P_  (.D(_0208_),
    .CK(clknet_leaf_38_clk),
    .Q(net200),
    .QN(_1738_));
 DFF_X2 \counters[43]$_SDFFE_PP0P_  (.D(_0209_),
    .CK(clknet_leaf_0_clk),
    .Q(net201),
    .QN(_1737_));
 DFF_X1 \counters[44]$_SDFFE_PP0P_  (.D(_0210_),
    .CK(clknet_leaf_38_clk),
    .Q(net202),
    .QN(_1736_));
 DFF_X1 \counters[45]$_SDFFE_PP0P_  (.D(_0211_),
    .CK(clknet_leaf_38_clk),
    .Q(net203),
    .QN(_1735_));
 DFF_X1 \counters[46]$_SDFFE_PP0P_  (.D(_0212_),
    .CK(clknet_leaf_37_clk),
    .Q(net204),
    .QN(_1734_));
 DFF_X2 \counters[47]$_SDFFE_PP0P_  (.D(_0213_),
    .CK(clknet_leaf_38_clk),
    .Q(net205),
    .QN(_1733_));
 DFF_X2 \counters[48]$_SDFFE_PP0P_  (.D(_0214_),
    .CK(clknet_leaf_38_clk),
    .Q(net206),
    .QN(_1732_));
 DFF_X2 \counters[49]$_SDFFE_PP0P_  (.D(_0215_),
    .CK(clknet_leaf_37_clk),
    .Q(net207),
    .QN(_1731_));
 DFF_X1 \counters[4]$_SDFFE_PP0P_  (.D(_0216_),
    .CK(clknet_leaf_39_clk),
    .Q(net208),
    .QN(_1730_));
 DFF_X1 \counters[50]$_SDFFE_PP0P_  (.D(_0217_),
    .CK(clknet_leaf_36_clk),
    .Q(net209),
    .QN(_1729_));
 DFF_X1 \counters[51]$_SDFFE_PP0P_  (.D(_0218_),
    .CK(clknet_leaf_31_clk),
    .Q(net210),
    .QN(_1728_));
 DFF_X1 \counters[52]$_SDFFE_PP0P_  (.D(_0219_),
    .CK(clknet_leaf_31_clk),
    .Q(net211),
    .QN(_1727_));
 DFF_X2 \counters[53]$_SDFFE_PP0P_  (.D(_0220_),
    .CK(clknet_leaf_31_clk),
    .Q(net212),
    .QN(_1726_));
 DFF_X1 \counters[54]$_SDFFE_PP0P_  (.D(_0221_),
    .CK(clknet_leaf_31_clk),
    .Q(net213),
    .QN(_1725_));
 DFF_X1 \counters[55]$_SDFFE_PP0P_  (.D(_0222_),
    .CK(clknet_leaf_36_clk),
    .Q(net214),
    .QN(_1724_));
 DFF_X1 \counters[56]$_SDFFE_PP0P_  (.D(_0223_),
    .CK(clknet_leaf_36_clk),
    .Q(net215),
    .QN(_1723_));
 DFF_X1 \counters[57]$_SDFFE_PP0P_  (.D(_0224_),
    .CK(clknet_leaf_37_clk),
    .Q(net216),
    .QN(_1722_));
 DFF_X2 \counters[58]$_SDFFE_PP0P_  (.D(_0225_),
    .CK(clknet_leaf_36_clk),
    .Q(net217),
    .QN(_1721_));
 DFF_X1 \counters[59]$_SDFFE_PP0P_  (.D(_0226_),
    .CK(clknet_leaf_36_clk),
    .Q(net218),
    .QN(_1720_));
 DFF_X2 \counters[5]$_SDFFE_PP0P_  (.D(_0227_),
    .CK(clknet_leaf_1_clk),
    .Q(net219),
    .QN(_1719_));
 DFF_X2 \counters[60]$_SDFFE_PP0P_  (.D(_0228_),
    .CK(clknet_leaf_37_clk),
    .Q(net220),
    .QN(_1718_));
 DFF_X2 \counters[61]$_SDFFE_PP0P_  (.D(_0229_),
    .CK(clknet_leaf_37_clk),
    .Q(net221),
    .QN(_1717_));
 DFF_X2 \counters[62]$_SDFFE_PP0P_  (.D(_0230_),
    .CK(clknet_leaf_35_clk),
    .Q(net222),
    .QN(_1716_));
 DFF_X1 \counters[63]$_SDFFE_PP0P_  (.D(_0231_),
    .CK(clknet_leaf_37_clk),
    .Q(net223),
    .QN(_1715_));
 DFF_X2 \counters[64]$_SDFFE_PP0P_  (.D(_0232_),
    .CK(clknet_leaf_7_clk),
    .Q(net224),
    .QN(_0002_));
 DFF_X2 \counters[65]$_SDFFE_PP0P_  (.D(_0233_),
    .CK(clknet_leaf_7_clk),
    .Q(net225),
    .QN(_1714_));
 DFF_X2 \counters[66]$_SDFFE_PP0P_  (.D(_0234_),
    .CK(clknet_leaf_7_clk),
    .Q(net226),
    .QN(_1713_));
 DFF_X1 \counters[67]$_SDFFE_PP0P_  (.D(_0235_),
    .CK(clknet_leaf_6_clk),
    .Q(net227),
    .QN(_1712_));
 DFF_X2 \counters[68]$_SDFFE_PP0P_  (.D(_0236_),
    .CK(clknet_leaf_8_clk),
    .Q(net228),
    .QN(_1711_));
 DFF_X2 \counters[69]$_SDFFE_PP0P_  (.D(_0237_),
    .CK(clknet_leaf_7_clk),
    .Q(net229),
    .QN(_1710_));
 DFF_X1 \counters[6]$_SDFFE_PP0P_  (.D(_0238_),
    .CK(clknet_leaf_1_clk),
    .Q(net230),
    .QN(_1709_));
 DFF_X1 \counters[70]$_SDFFE_PP0P_  (.D(_0239_),
    .CK(clknet_leaf_8_clk),
    .Q(net231),
    .QN(_1708_));
 DFF_X1 \counters[71]$_SDFFE_PP0P_  (.D(_0240_),
    .CK(clknet_leaf_8_clk),
    .Q(net232),
    .QN(_1707_));
 DFF_X1 \counters[72]$_SDFFE_PP0P_  (.D(_0241_),
    .CK(clknet_leaf_8_clk),
    .Q(net233),
    .QN(_1706_));
 DFF_X1 \counters[73]$_SDFFE_PP0P_  (.D(_0242_),
    .CK(clknet_leaf_8_clk),
    .Q(net234),
    .QN(_1705_));
 DFF_X1 \counters[74]$_SDFFE_PP0P_  (.D(_0243_),
    .CK(clknet_leaf_7_clk),
    .Q(net235),
    .QN(_1704_));
 DFF_X1 \counters[75]$_SDFFE_PP0P_  (.D(_0244_),
    .CK(clknet_leaf_9_clk),
    .Q(net236),
    .QN(_1703_));
 DFF_X1 \counters[76]$_SDFFE_PP0P_  (.D(_0245_),
    .CK(clknet_leaf_8_clk),
    .Q(net237),
    .QN(_1702_));
 DFF_X2 \counters[77]$_SDFFE_PP0P_  (.D(_0246_),
    .CK(clknet_leaf_9_clk),
    .Q(net238),
    .QN(_1701_));
 DFF_X2 \counters[78]$_SDFFE_PP0P_  (.D(_0247_),
    .CK(clknet_leaf_9_clk),
    .Q(net239),
    .QN(_1700_));
 DFF_X1 \counters[79]$_SDFFE_PP0P_  (.D(_0248_),
    .CK(clknet_leaf_9_clk),
    .Q(net240),
    .QN(_1699_));
 DFF_X1 \counters[7]$_SDFFE_PP0P_  (.D(_0249_),
    .CK(clknet_leaf_1_clk),
    .Q(net241),
    .QN(_1698_));
 DFF_X1 \counters[80]$_SDFFE_PP0P_  (.D(_0250_),
    .CK(clknet_leaf_10_clk),
    .Q(net242),
    .QN(_1697_));
 DFF_X1 \counters[81]$_SDFFE_PP0P_  (.D(_0251_),
    .CK(clknet_leaf_9_clk),
    .Q(net243),
    .QN(_1696_));
 DFF_X1 \counters[82]$_SDFFE_PP0P_  (.D(_0252_),
    .CK(clknet_leaf_9_clk),
    .Q(net244),
    .QN(_1695_));
 DFF_X2 \counters[83]$_SDFFE_PP0P_  (.D(_0253_),
    .CK(clknet_leaf_12_clk),
    .Q(net245),
    .QN(_1694_));
 DFF_X2 \counters[84]$_SDFFE_PP0P_  (.D(_0254_),
    .CK(clknet_leaf_10_clk),
    .Q(net246),
    .QN(_1693_));
 DFF_X1 \counters[85]$_SDFFE_PP0P_  (.D(_0255_),
    .CK(clknet_leaf_10_clk),
    .Q(net247),
    .QN(_1692_));
 DFF_X1 \counters[86]$_SDFFE_PP0P_  (.D(_0256_),
    .CK(clknet_leaf_10_clk),
    .Q(net248),
    .QN(_1691_));
 DFF_X1 \counters[87]$_SDFFE_PP0P_  (.D(_0257_),
    .CK(clknet_leaf_10_clk),
    .Q(net249),
    .QN(_1690_));
 DFF_X2 \counters[88]$_SDFFE_PP0P_  (.D(_0258_),
    .CK(clknet_leaf_10_clk),
    .Q(net250),
    .QN(_1689_));
 DFF_X2 \counters[89]$_SDFFE_PP0P_  (.D(_0259_),
    .CK(clknet_leaf_12_clk),
    .Q(net251),
    .QN(_1688_));
 DFF_X2 \counters[8]$_SDFFE_PP0P_  (.D(_0260_),
    .CK(clknet_leaf_2_clk),
    .Q(net252),
    .QN(_1687_));
 DFF_X1 \counters[90]$_SDFFE_PP0P_  (.D(_0261_),
    .CK(clknet_leaf_11_clk),
    .Q(net253),
    .QN(_1686_));
 DFF_X1 \counters[91]$_SDFFE_PP0P_  (.D(_0262_),
    .CK(clknet_leaf_11_clk),
    .Q(net254),
    .QN(_1685_));
 DFF_X1 \counters[92]$_SDFFE_PP0P_  (.D(_0263_),
    .CK(clknet_leaf_11_clk),
    .Q(net255),
    .QN(_1684_));
 DFF_X2 \counters[93]$_SDFFE_PP0P_  (.D(_0264_),
    .CK(clknet_leaf_11_clk),
    .Q(net256),
    .QN(_1683_));
 DFF_X1 \counters[94]$_SDFFE_PP0P_  (.D(_0265_),
    .CK(clknet_leaf_10_clk),
    .Q(net257),
    .QN(_1682_));
 DFF_X1 \counters[95]$_SDFFE_PP0P_  (.D(_0266_),
    .CK(clknet_leaf_12_clk),
    .Q(net258),
    .QN(_1681_));
 DFF_X2 \counters[96]$_SDFFE_PP0P_  (.D(_0267_),
    .CK(clknet_leaf_5_clk),
    .Q(net259),
    .QN(_0004_));
 DFF_X1 \counters[97]$_SDFFE_PP0P_  (.D(_0268_),
    .CK(clknet_leaf_5_clk),
    .Q(net260),
    .QN(_1680_));
 DFF_X1 \counters[98]$_SDFFE_PP0P_  (.D(_0269_),
    .CK(clknet_leaf_6_clk),
    .Q(net261),
    .QN(_1679_));
 DFF_X1 \counters[99]$_SDFFE_PP0P_  (.D(_0270_),
    .CK(clknet_leaf_6_clk),
    .Q(net262),
    .QN(_1678_));
 DFF_X1 \counters[9]$_SDFFE_PP0P_  (.D(_0271_),
    .CK(clknet_leaf_1_clk),
    .Q(net263),
    .QN(_1677_));
 DFF_X2 \prev_event_inc[0]$_SDFFE_PN0N_  (.D(_0272_),
    .CK(clknet_leaf_0_clk),
    .Q(\prev_event_inc[0] ),
    .QN(_1676_));
 DFF_X1 \prev_event_inc[1]$_SDFFE_PN0N_  (.D(_0273_),
    .CK(clknet_leaf_0_clk),
    .Q(\prev_event_inc[1] ),
    .QN(_1675_));
 DFF_X2 \prev_event_inc[2]$_SDFFE_PN0N_  (.D(_0274_),
    .CK(clknet_leaf_7_clk),
    .Q(\prev_event_inc[2] ),
    .QN(_1674_));
 DFF_X2 \prev_event_inc[3]$_SDFFE_PN0N_  (.D(_0275_),
    .CK(clknet_leaf_5_clk),
    .Q(\prev_event_inc[3] ),
    .QN(_1673_));
 DFF_X1 \prev_event_inc[4]$_SDFFE_PN0N_  (.D(_0276_),
    .CK(clknet_leaf_13_clk),
    .Q(\prev_event_inc[4] ),
    .QN(_1672_));
 DFF_X1 \prev_event_inc[5]$_SDFFE_PN0N_  (.D(_0277_),
    .CK(clknet_leaf_32_clk),
    .Q(\prev_event_inc[5] ),
    .QN(_1671_));
 DFF_X2 \prev_event_inc[6]$_SDFFE_PN0N_  (.D(_0278_),
    .CK(clknet_leaf_14_clk),
    .Q(\prev_event_inc[6] ),
    .QN(_1670_));
 DFF_X1 \prev_event_inc[7]$_SDFFE_PN0N_  (.D(_0279_),
    .CK(clknet_leaf_22_clk),
    .Q(\prev_event_inc[7] ),
    .QN(_1669_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_111 ();
 BUF_X1 input1 (.A(counter_sel[6]),
    .Z(net1));
 BUF_X1 input2 (.A(counter_sel[7]),
    .Z(net2));
 BUF_X2 input3 (.A(event_inc[0]),
    .Z(net3));
 BUF_X1 input4 (.A(event_inc[1]),
    .Z(net4));
 BUF_X1 input5 (.A(event_inc[5]),
    .Z(net5));
 BUF_X1 input6 (.A(event_inc[6]),
    .Z(net6));
 CLKBUF_X2 input7 (.A(rst_n),
    .Z(net7));
 BUF_X1 output8 (.A(net8),
    .Z(all_counts[0]));
 BUF_X1 output9 (.A(net9),
    .Z(all_counts[100]));
 BUF_X1 output10 (.A(net10),
    .Z(all_counts[101]));
 BUF_X1 output11 (.A(net11),
    .Z(all_counts[102]));
 BUF_X1 output12 (.A(net12),
    .Z(all_counts[103]));
 BUF_X1 output13 (.A(net13),
    .Z(all_counts[104]));
 BUF_X1 output14 (.A(net14),
    .Z(all_counts[105]));
 BUF_X1 output15 (.A(net15),
    .Z(all_counts[106]));
 BUF_X1 output16 (.A(net16),
    .Z(all_counts[107]));
 BUF_X1 output17 (.A(net17),
    .Z(all_counts[108]));
 BUF_X1 output18 (.A(net18),
    .Z(all_counts[109]));
 BUF_X1 output19 (.A(net19),
    .Z(all_counts[10]));
 BUF_X1 output20 (.A(net20),
    .Z(all_counts[110]));
 BUF_X1 output21 (.A(net21),
    .Z(all_counts[111]));
 BUF_X1 output22 (.A(net22),
    .Z(all_counts[112]));
 BUF_X1 output23 (.A(net23),
    .Z(all_counts[113]));
 BUF_X1 output24 (.A(net24),
    .Z(all_counts[114]));
 BUF_X1 output25 (.A(net25),
    .Z(all_counts[115]));
 BUF_X1 output26 (.A(net26),
    .Z(all_counts[116]));
 BUF_X1 output27 (.A(net27),
    .Z(all_counts[117]));
 BUF_X1 output28 (.A(net28),
    .Z(all_counts[118]));
 BUF_X1 output29 (.A(net29),
    .Z(all_counts[119]));
 BUF_X1 output30 (.A(net30),
    .Z(all_counts[11]));
 BUF_X1 output31 (.A(net31),
    .Z(all_counts[120]));
 BUF_X1 output32 (.A(net32),
    .Z(all_counts[121]));
 BUF_X1 output33 (.A(net33),
    .Z(all_counts[122]));
 BUF_X1 output34 (.A(net34),
    .Z(all_counts[123]));
 BUF_X1 output35 (.A(net35),
    .Z(all_counts[124]));
 BUF_X1 output36 (.A(net36),
    .Z(all_counts[125]));
 BUF_X1 output37 (.A(net37),
    .Z(all_counts[126]));
 BUF_X1 output38 (.A(net38),
    .Z(all_counts[127]));
 BUF_X1 output39 (.A(net39),
    .Z(all_counts[128]));
 BUF_X1 output40 (.A(net40),
    .Z(all_counts[129]));
 BUF_X1 output41 (.A(net41),
    .Z(all_counts[12]));
 BUF_X1 output42 (.A(net42),
    .Z(all_counts[130]));
 BUF_X1 output43 (.A(net43),
    .Z(all_counts[131]));
 BUF_X1 output44 (.A(net44),
    .Z(all_counts[132]));
 BUF_X1 output45 (.A(net45),
    .Z(all_counts[133]));
 BUF_X1 output46 (.A(net46),
    .Z(all_counts[134]));
 BUF_X1 output47 (.A(net47),
    .Z(all_counts[135]));
 BUF_X1 output48 (.A(net48),
    .Z(all_counts[136]));
 BUF_X1 output49 (.A(net49),
    .Z(all_counts[137]));
 BUF_X1 output50 (.A(net50),
    .Z(all_counts[138]));
 BUF_X1 output51 (.A(net51),
    .Z(all_counts[139]));
 BUF_X1 output52 (.A(net52),
    .Z(all_counts[13]));
 BUF_X1 output53 (.A(net53),
    .Z(all_counts[140]));
 BUF_X1 output54 (.A(net54),
    .Z(all_counts[141]));
 BUF_X1 output55 (.A(net55),
    .Z(all_counts[142]));
 BUF_X1 output56 (.A(net56),
    .Z(all_counts[143]));
 BUF_X1 output57 (.A(net57),
    .Z(all_counts[144]));
 BUF_X1 output58 (.A(net58),
    .Z(all_counts[145]));
 BUF_X1 output59 (.A(net59),
    .Z(all_counts[146]));
 BUF_X1 output60 (.A(net60),
    .Z(all_counts[147]));
 BUF_X1 output61 (.A(net61),
    .Z(all_counts[148]));
 BUF_X1 output62 (.A(net62),
    .Z(all_counts[149]));
 BUF_X1 output63 (.A(net63),
    .Z(all_counts[14]));
 BUF_X1 output64 (.A(net64),
    .Z(all_counts[150]));
 BUF_X1 output65 (.A(net65),
    .Z(all_counts[151]));
 BUF_X1 output66 (.A(net66),
    .Z(all_counts[152]));
 BUF_X1 output67 (.A(net67),
    .Z(all_counts[153]));
 BUF_X1 output68 (.A(net68),
    .Z(all_counts[154]));
 BUF_X1 output69 (.A(net69),
    .Z(all_counts[155]));
 BUF_X1 output70 (.A(net70),
    .Z(all_counts[156]));
 BUF_X1 output71 (.A(net71),
    .Z(all_counts[157]));
 BUF_X1 output72 (.A(net72),
    .Z(all_counts[158]));
 BUF_X1 output73 (.A(net73),
    .Z(all_counts[159]));
 BUF_X1 output74 (.A(net74),
    .Z(all_counts[15]));
 BUF_X1 output75 (.A(net75),
    .Z(all_counts[160]));
 BUF_X1 output76 (.A(net76),
    .Z(all_counts[161]));
 BUF_X1 output77 (.A(net77),
    .Z(all_counts[162]));
 BUF_X1 output78 (.A(net78),
    .Z(all_counts[163]));
 BUF_X1 output79 (.A(net79),
    .Z(all_counts[164]));
 BUF_X1 output80 (.A(net80),
    .Z(all_counts[165]));
 BUF_X1 output81 (.A(net81),
    .Z(all_counts[166]));
 BUF_X1 output82 (.A(net82),
    .Z(all_counts[167]));
 BUF_X1 output83 (.A(net83),
    .Z(all_counts[168]));
 BUF_X1 output84 (.A(net84),
    .Z(all_counts[169]));
 BUF_X1 output85 (.A(net85),
    .Z(all_counts[16]));
 BUF_X1 output86 (.A(net86),
    .Z(all_counts[170]));
 BUF_X1 output87 (.A(net87),
    .Z(all_counts[171]));
 BUF_X1 output88 (.A(net88),
    .Z(all_counts[172]));
 BUF_X1 output89 (.A(net89),
    .Z(all_counts[173]));
 BUF_X1 output90 (.A(net90),
    .Z(all_counts[174]));
 BUF_X1 output91 (.A(net91),
    .Z(all_counts[175]));
 BUF_X1 output92 (.A(net92),
    .Z(all_counts[176]));
 BUF_X1 output93 (.A(net93),
    .Z(all_counts[177]));
 BUF_X1 output94 (.A(net94),
    .Z(all_counts[178]));
 BUF_X1 output95 (.A(net95),
    .Z(all_counts[179]));
 BUF_X1 output96 (.A(net96),
    .Z(all_counts[17]));
 BUF_X1 output97 (.A(net97),
    .Z(all_counts[180]));
 BUF_X1 output98 (.A(net98),
    .Z(all_counts[181]));
 BUF_X1 output99 (.A(net99),
    .Z(all_counts[182]));
 BUF_X1 output100 (.A(net100),
    .Z(all_counts[183]));
 BUF_X1 output101 (.A(net101),
    .Z(all_counts[184]));
 BUF_X1 output102 (.A(net102),
    .Z(all_counts[185]));
 BUF_X1 output103 (.A(net103),
    .Z(all_counts[186]));
 BUF_X1 output104 (.A(net104),
    .Z(all_counts[187]));
 BUF_X1 output105 (.A(net105),
    .Z(all_counts[188]));
 BUF_X1 output106 (.A(net106),
    .Z(all_counts[189]));
 BUF_X1 output107 (.A(net107),
    .Z(all_counts[18]));
 BUF_X1 output108 (.A(net108),
    .Z(all_counts[190]));
 BUF_X1 output109 (.A(net109),
    .Z(all_counts[191]));
 BUF_X1 output110 (.A(net110),
    .Z(all_counts[192]));
 BUF_X1 output111 (.A(net111),
    .Z(all_counts[193]));
 BUF_X1 output112 (.A(net112),
    .Z(all_counts[194]));
 BUF_X1 output113 (.A(net113),
    .Z(all_counts[195]));
 BUF_X1 output114 (.A(net114),
    .Z(all_counts[196]));
 BUF_X1 output115 (.A(net115),
    .Z(all_counts[197]));
 BUF_X1 output116 (.A(net116),
    .Z(all_counts[198]));
 BUF_X1 output117 (.A(net117),
    .Z(all_counts[199]));
 BUF_X1 output118 (.A(net118),
    .Z(all_counts[19]));
 BUF_X1 output119 (.A(net119),
    .Z(all_counts[1]));
 BUF_X1 output120 (.A(net120),
    .Z(all_counts[200]));
 BUF_X1 output121 (.A(net121),
    .Z(all_counts[201]));
 BUF_X1 output122 (.A(net122),
    .Z(all_counts[202]));
 BUF_X1 output123 (.A(net123),
    .Z(all_counts[203]));
 BUF_X1 output124 (.A(net124),
    .Z(all_counts[204]));
 BUF_X1 output125 (.A(net125),
    .Z(all_counts[205]));
 BUF_X1 output126 (.A(net126),
    .Z(all_counts[206]));
 BUF_X1 output127 (.A(net127),
    .Z(all_counts[207]));
 BUF_X1 output128 (.A(net128),
    .Z(all_counts[208]));
 BUF_X1 output129 (.A(net129),
    .Z(all_counts[209]));
 BUF_X1 output130 (.A(net130),
    .Z(all_counts[20]));
 BUF_X1 output131 (.A(net131),
    .Z(all_counts[210]));
 BUF_X1 output132 (.A(net132),
    .Z(all_counts[211]));
 BUF_X1 output133 (.A(net133),
    .Z(all_counts[212]));
 BUF_X1 output134 (.A(net134),
    .Z(all_counts[213]));
 BUF_X1 output135 (.A(net135),
    .Z(all_counts[214]));
 BUF_X1 output136 (.A(net136),
    .Z(all_counts[215]));
 BUF_X1 output137 (.A(net137),
    .Z(all_counts[216]));
 BUF_X1 output138 (.A(net138),
    .Z(all_counts[217]));
 BUF_X1 output139 (.A(net139),
    .Z(all_counts[218]));
 BUF_X1 output140 (.A(net140),
    .Z(all_counts[219]));
 BUF_X1 output141 (.A(net141),
    .Z(all_counts[21]));
 BUF_X1 output142 (.A(net142),
    .Z(all_counts[220]));
 BUF_X1 output143 (.A(net143),
    .Z(all_counts[221]));
 BUF_X1 output144 (.A(net144),
    .Z(all_counts[222]));
 BUF_X1 output145 (.A(net145),
    .Z(all_counts[223]));
 BUF_X1 output146 (.A(net146),
    .Z(all_counts[224]));
 BUF_X1 output147 (.A(net147),
    .Z(all_counts[225]));
 BUF_X1 output148 (.A(net148),
    .Z(all_counts[226]));
 BUF_X1 output149 (.A(net149),
    .Z(all_counts[227]));
 BUF_X1 output150 (.A(net150),
    .Z(all_counts[228]));
 BUF_X1 output151 (.A(net151),
    .Z(all_counts[229]));
 BUF_X1 output152 (.A(net152),
    .Z(all_counts[22]));
 BUF_X1 output153 (.A(net153),
    .Z(all_counts[230]));
 BUF_X1 output154 (.A(net154),
    .Z(all_counts[231]));
 BUF_X1 output155 (.A(net155),
    .Z(all_counts[232]));
 BUF_X1 output156 (.A(net156),
    .Z(all_counts[233]));
 BUF_X1 output157 (.A(net157),
    .Z(all_counts[234]));
 BUF_X1 output158 (.A(net158),
    .Z(all_counts[235]));
 BUF_X1 output159 (.A(net159),
    .Z(all_counts[236]));
 BUF_X1 output160 (.A(net160),
    .Z(all_counts[237]));
 BUF_X1 output161 (.A(net161),
    .Z(all_counts[238]));
 BUF_X1 output162 (.A(net162),
    .Z(all_counts[239]));
 BUF_X1 output163 (.A(net163),
    .Z(all_counts[23]));
 BUF_X1 output164 (.A(net164),
    .Z(all_counts[240]));
 BUF_X1 output165 (.A(net165),
    .Z(all_counts[241]));
 BUF_X1 output166 (.A(net166),
    .Z(all_counts[242]));
 BUF_X1 output167 (.A(net167),
    .Z(all_counts[243]));
 BUF_X1 output168 (.A(net168),
    .Z(all_counts[244]));
 BUF_X1 output169 (.A(net169),
    .Z(all_counts[245]));
 BUF_X1 output170 (.A(net170),
    .Z(all_counts[246]));
 BUF_X1 output171 (.A(net171),
    .Z(all_counts[247]));
 BUF_X1 output172 (.A(net172),
    .Z(all_counts[248]));
 BUF_X1 output173 (.A(net173),
    .Z(all_counts[249]));
 BUF_X1 output174 (.A(net174),
    .Z(all_counts[24]));
 BUF_X1 output175 (.A(net175),
    .Z(all_counts[250]));
 BUF_X1 output176 (.A(net176),
    .Z(all_counts[251]));
 BUF_X1 output177 (.A(net177),
    .Z(all_counts[252]));
 BUF_X1 output178 (.A(net178),
    .Z(all_counts[253]));
 BUF_X1 output179 (.A(net179),
    .Z(all_counts[254]));
 BUF_X1 output180 (.A(net180),
    .Z(all_counts[255]));
 BUF_X1 output181 (.A(net181),
    .Z(all_counts[25]));
 BUF_X1 output182 (.A(net182),
    .Z(all_counts[26]));
 BUF_X1 output183 (.A(net183),
    .Z(all_counts[27]));
 BUF_X1 output184 (.A(net184),
    .Z(all_counts[28]));
 BUF_X1 output185 (.A(net185),
    .Z(all_counts[29]));
 BUF_X1 output186 (.A(net186),
    .Z(all_counts[2]));
 BUF_X1 output187 (.A(net187),
    .Z(all_counts[30]));
 BUF_X1 output188 (.A(net188),
    .Z(all_counts[31]));
 BUF_X1 output189 (.A(net189),
    .Z(all_counts[32]));
 BUF_X1 output190 (.A(net190),
    .Z(all_counts[33]));
 BUF_X1 output191 (.A(net191),
    .Z(all_counts[34]));
 BUF_X1 output192 (.A(net192),
    .Z(all_counts[35]));
 BUF_X1 output193 (.A(net193),
    .Z(all_counts[36]));
 BUF_X1 output194 (.A(net194),
    .Z(all_counts[37]));
 BUF_X1 output195 (.A(net195),
    .Z(all_counts[38]));
 BUF_X1 output196 (.A(net196),
    .Z(all_counts[39]));
 BUF_X1 output197 (.A(net197),
    .Z(all_counts[3]));
 BUF_X1 output198 (.A(net198),
    .Z(all_counts[40]));
 BUF_X1 output199 (.A(net199),
    .Z(all_counts[41]));
 BUF_X1 output200 (.A(net200),
    .Z(all_counts[42]));
 BUF_X1 output201 (.A(net201),
    .Z(all_counts[43]));
 BUF_X1 output202 (.A(net202),
    .Z(all_counts[44]));
 BUF_X1 output203 (.A(net203),
    .Z(all_counts[45]));
 BUF_X1 output204 (.A(net204),
    .Z(all_counts[46]));
 BUF_X1 output205 (.A(net205),
    .Z(all_counts[47]));
 BUF_X1 output206 (.A(net206),
    .Z(all_counts[48]));
 BUF_X1 output207 (.A(net207),
    .Z(all_counts[49]));
 BUF_X1 output208 (.A(net208),
    .Z(all_counts[4]));
 BUF_X1 output209 (.A(net209),
    .Z(all_counts[50]));
 BUF_X1 output210 (.A(net210),
    .Z(all_counts[51]));
 BUF_X1 output211 (.A(net211),
    .Z(all_counts[52]));
 BUF_X1 output212 (.A(net212),
    .Z(all_counts[53]));
 BUF_X1 output213 (.A(net213),
    .Z(all_counts[54]));
 BUF_X1 output214 (.A(net214),
    .Z(all_counts[55]));
 BUF_X1 output215 (.A(net215),
    .Z(all_counts[56]));
 BUF_X1 output216 (.A(net216),
    .Z(all_counts[57]));
 BUF_X1 output217 (.A(net217),
    .Z(all_counts[58]));
 BUF_X1 output218 (.A(net218),
    .Z(all_counts[59]));
 BUF_X1 output219 (.A(net219),
    .Z(all_counts[5]));
 BUF_X1 output220 (.A(net220),
    .Z(all_counts[60]));
 BUF_X1 output221 (.A(net221),
    .Z(all_counts[61]));
 BUF_X1 output222 (.A(net222),
    .Z(all_counts[62]));
 BUF_X1 output223 (.A(net223),
    .Z(all_counts[63]));
 BUF_X1 output224 (.A(net224),
    .Z(all_counts[64]));
 BUF_X1 output225 (.A(net225),
    .Z(all_counts[65]));
 BUF_X1 output226 (.A(net226),
    .Z(all_counts[66]));
 BUF_X1 output227 (.A(net227),
    .Z(all_counts[67]));
 BUF_X1 output228 (.A(net228),
    .Z(all_counts[68]));
 BUF_X1 output229 (.A(net229),
    .Z(all_counts[69]));
 BUF_X1 output230 (.A(net230),
    .Z(all_counts[6]));
 BUF_X1 output231 (.A(net231),
    .Z(all_counts[70]));
 BUF_X1 output232 (.A(net232),
    .Z(all_counts[71]));
 BUF_X1 output233 (.A(net233),
    .Z(all_counts[72]));
 BUF_X1 output234 (.A(net234),
    .Z(all_counts[73]));
 BUF_X1 output235 (.A(net235),
    .Z(all_counts[74]));
 BUF_X1 output236 (.A(net236),
    .Z(all_counts[75]));
 BUF_X1 output237 (.A(net237),
    .Z(all_counts[76]));
 BUF_X1 output238 (.A(net238),
    .Z(all_counts[77]));
 BUF_X1 output239 (.A(net239),
    .Z(all_counts[78]));
 BUF_X1 output240 (.A(net240),
    .Z(all_counts[79]));
 BUF_X1 output241 (.A(net241),
    .Z(all_counts[7]));
 BUF_X1 output242 (.A(net242),
    .Z(all_counts[80]));
 BUF_X1 output243 (.A(net243),
    .Z(all_counts[81]));
 BUF_X1 output244 (.A(net244),
    .Z(all_counts[82]));
 BUF_X1 output245 (.A(net245),
    .Z(all_counts[83]));
 BUF_X1 output246 (.A(net246),
    .Z(all_counts[84]));
 BUF_X1 output247 (.A(net247),
    .Z(all_counts[85]));
 BUF_X1 output248 (.A(net248),
    .Z(all_counts[86]));
 BUF_X1 output249 (.A(net249),
    .Z(all_counts[87]));
 BUF_X1 output250 (.A(net250),
    .Z(all_counts[88]));
 BUF_X1 output251 (.A(net251),
    .Z(all_counts[89]));
 BUF_X1 output252 (.A(net252),
    .Z(all_counts[8]));
 BUF_X1 output253 (.A(net253),
    .Z(all_counts[90]));
 BUF_X1 output254 (.A(net254),
    .Z(all_counts[91]));
 BUF_X1 output255 (.A(net255),
    .Z(all_counts[92]));
 BUF_X1 output256 (.A(net256),
    .Z(all_counts[93]));
 BUF_X1 output257 (.A(net257),
    .Z(all_counts[94]));
 BUF_X1 output258 (.A(net258),
    .Z(all_counts[95]));
 BUF_X1 output259 (.A(net259),
    .Z(all_counts[96]));
 BUF_X1 output260 (.A(net260),
    .Z(all_counts[97]));
 BUF_X1 output261 (.A(net261),
    .Z(all_counts[98]));
 BUF_X1 output262 (.A(net262),
    .Z(all_counts[99]));
 BUF_X1 output263 (.A(net263),
    .Z(all_counts[9]));
 BUF_X1 output264 (.A(net264),
    .Z(count_value[0]));
 BUF_X1 output265 (.A(net265),
    .Z(count_value[10]));
 BUF_X1 output266 (.A(net266),
    .Z(count_value[11]));
 BUF_X1 output267 (.A(net267),
    .Z(count_value[12]));
 BUF_X1 output268 (.A(net268),
    .Z(count_value[13]));
 BUF_X1 output269 (.A(net269),
    .Z(count_value[14]));
 BUF_X1 output270 (.A(net270),
    .Z(count_value[15]));
 BUF_X1 output271 (.A(net271),
    .Z(count_value[16]));
 BUF_X1 output272 (.A(net272),
    .Z(count_value[17]));
 BUF_X1 output273 (.A(net273),
    .Z(count_value[18]));
 BUF_X1 output274 (.A(net274),
    .Z(count_value[19]));
 BUF_X1 output275 (.A(net275),
    .Z(count_value[1]));
 BUF_X1 output276 (.A(net276),
    .Z(count_value[20]));
 BUF_X1 output277 (.A(net277),
    .Z(count_value[21]));
 BUF_X1 output278 (.A(net278),
    .Z(count_value[22]));
 BUF_X1 output279 (.A(net279),
    .Z(count_value[23]));
 BUF_X1 output280 (.A(net280),
    .Z(count_value[24]));
 BUF_X1 output281 (.A(net281),
    .Z(count_value[25]));
 BUF_X1 output282 (.A(net282),
    .Z(count_value[26]));
 BUF_X1 output283 (.A(net283),
    .Z(count_value[27]));
 BUF_X1 output284 (.A(net284),
    .Z(count_value[28]));
 BUF_X1 output285 (.A(net285),
    .Z(count_value[29]));
 BUF_X1 output286 (.A(net286),
    .Z(count_value[2]));
 BUF_X1 output287 (.A(net287),
    .Z(count_value[30]));
 BUF_X1 output288 (.A(net288),
    .Z(count_value[31]));
 BUF_X1 output289 (.A(net289),
    .Z(count_value[3]));
 BUF_X1 output290 (.A(net290),
    .Z(count_value[4]));
 BUF_X1 output291 (.A(net291),
    .Z(count_value[5]));
 BUF_X1 output292 (.A(net292),
    .Z(count_value[6]));
 BUF_X1 output293 (.A(net293),
    .Z(count_value[7]));
 BUF_X1 output294 (.A(net294),
    .Z(count_value[8]));
 BUF_X1 output295 (.A(net295),
    .Z(count_value[9]));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_leaf_0_clk));
 CLKBUF_X1 clkload1 (.A(clknet_leaf_1_clk));
 CLKBUF_X1 clkload2 (.A(clknet_leaf_2_clk));
 CLKBUF_X1 clkload3 (.A(clknet_leaf_3_clk));
 INV_X1 clkload4 (.A(clknet_leaf_34_clk));
 CLKBUF_X1 clkload5 (.A(clknet_leaf_35_clk));
 CLKBUF_X1 clkload6 (.A(clknet_leaf_36_clk));
 CLKBUF_X1 clkload7 (.A(clknet_leaf_37_clk));
 CLKBUF_X1 clkload8 (.A(clknet_leaf_38_clk));
 CLKBUF_X1 clkload9 (.A(clknet_leaf_4_clk));
 CLKBUF_X1 clkload10 (.A(clknet_leaf_5_clk));
 CLKBUF_X1 clkload11 (.A(clknet_leaf_7_clk));
 CLKBUF_X1 clkload12 (.A(clknet_leaf_8_clk));
 CLKBUF_X1 clkload13 (.A(clknet_leaf_9_clk));
 CLKBUF_X1 clkload14 (.A(clknet_leaf_10_clk));
 CLKBUF_X1 clkload15 (.A(clknet_leaf_11_clk));
 CLKBUF_X1 clkload16 (.A(clknet_leaf_12_clk));
 CLKBUF_X1 clkload17 (.A(clknet_leaf_13_clk));
 INV_X1 clkload18 (.A(clknet_leaf_24_clk));
 INV_X1 clkload19 (.A(clknet_leaf_25_clk));
 CLKBUF_X1 clkload20 (.A(clknet_leaf_26_clk));
 INV_X1 clkload21 (.A(clknet_leaf_27_clk));
 CLKBUF_X1 clkload22 (.A(clknet_leaf_28_clk));
 INV_X1 clkload23 (.A(clknet_leaf_29_clk));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_30_clk));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_31_clk));
 CLKBUF_X1 clkload26 (.A(clknet_leaf_32_clk));
 CLKBUF_X1 clkload27 (.A(clknet_leaf_14_clk));
 INV_X1 clkload28 (.A(clknet_leaf_15_clk));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_17_clk));
 CLKBUF_X1 clkload30 (.A(clknet_leaf_18_clk));
 INV_X1 clkload31 (.A(clknet_leaf_19_clk));
 INV_X1 clkload32 (.A(clknet_leaf_20_clk));
 CLKBUF_X1 clkload33 (.A(clknet_leaf_21_clk));
 INV_X1 clkload34 (.A(clknet_leaf_22_clk));
 CLKBUF_X1 clkload35 (.A(clknet_leaf_23_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X16 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_49 ();
 FILLCELL_X2 FILLER_0_60 ();
 FILLCELL_X4 FILLER_0_65 ();
 FILLCELL_X2 FILLER_0_69 ();
 FILLCELL_X8 FILLER_0_77 ();
 FILLCELL_X4 FILLER_0_85 ();
 FILLCELL_X1 FILLER_0_89 ();
 FILLCELL_X1 FILLER_0_111 ();
 FILLCELL_X1 FILLER_0_115 ();
 FILLCELL_X1 FILLER_0_119 ();
 FILLCELL_X4 FILLER_0_123 ();
 FILLCELL_X1 FILLER_0_127 ();
 FILLCELL_X1 FILLER_0_137 ();
 FILLCELL_X1 FILLER_0_141 ();
 FILLCELL_X1 FILLER_0_145 ();
 FILLCELL_X1 FILLER_0_149 ();
 FILLCELL_X1 FILLER_0_181 ();
 FILLCELL_X2 FILLER_0_252 ();
 FILLCELL_X2 FILLER_0_260 ();
 FILLCELL_X2 FILLER_0_265 ();
 FILLCELL_X4 FILLER_0_270 ();
 FILLCELL_X1 FILLER_0_274 ();
 FILLCELL_X8 FILLER_0_281 ();
 FILLCELL_X4 FILLER_0_292 ();
 FILLCELL_X2 FILLER_0_296 ();
 FILLCELL_X2 FILLER_0_301 ();
 FILLCELL_X8 FILLER_0_306 ();
 FILLCELL_X2 FILLER_0_314 ();
 FILLCELL_X1 FILLER_0_316 ();
 FILLCELL_X16 FILLER_0_320 ();
 FILLCELL_X1 FILLER_0_336 ();
 FILLCELL_X2 FILLER_0_340 ();
 FILLCELL_X1 FILLER_0_342 ();
 FILLCELL_X8 FILLER_0_346 ();
 FILLCELL_X2 FILLER_0_354 ();
 FILLCELL_X1 FILLER_0_356 ();
 FILLCELL_X32 FILLER_0_360 ();
 FILLCELL_X16 FILLER_0_392 ();
 FILLCELL_X8 FILLER_0_408 ();
 FILLCELL_X2 FILLER_0_416 ();
 FILLCELL_X1 FILLER_0_418 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X16 FILLER_1_65 ();
 FILLCELL_X4 FILLER_1_81 ();
 FILLCELL_X2 FILLER_1_85 ();
 FILLCELL_X1 FILLER_1_123 ();
 FILLCELL_X2 FILLER_1_144 ();
 FILLCELL_X1 FILLER_1_152 ();
 FILLCELL_X1 FILLER_1_170 ();
 FILLCELL_X1 FILLER_1_175 ();
 FILLCELL_X1 FILLER_1_193 ();
 FILLCELL_X2 FILLER_1_211 ();
 FILLCELL_X1 FILLER_1_233 ();
 FILLCELL_X16 FILLER_1_258 ();
 FILLCELL_X1 FILLER_1_274 ();
 FILLCELL_X2 FILLER_1_278 ();
 FILLCELL_X1 FILLER_1_280 ();
 FILLCELL_X8 FILLER_1_284 ();
 FILLCELL_X2 FILLER_1_292 ();
 FILLCELL_X32 FILLER_1_297 ();
 FILLCELL_X32 FILLER_1_329 ();
 FILLCELL_X32 FILLER_1_361 ();
 FILLCELL_X16 FILLER_1_393 ();
 FILLCELL_X8 FILLER_1_409 ();
 FILLCELL_X2 FILLER_1_417 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X2 FILLER_2_49 ();
 FILLCELL_X1 FILLER_2_51 ();
 FILLCELL_X16 FILLER_2_79 ();
 FILLCELL_X4 FILLER_2_95 ();
 FILLCELL_X2 FILLER_2_99 ();
 FILLCELL_X1 FILLER_2_101 ();
 FILLCELL_X1 FILLER_2_115 ();
 FILLCELL_X16 FILLER_2_125 ();
 FILLCELL_X8 FILLER_2_141 ();
 FILLCELL_X2 FILLER_2_155 ();
 FILLCELL_X1 FILLER_2_162 ();
 FILLCELL_X2 FILLER_2_166 ();
 FILLCELL_X4 FILLER_2_171 ();
 FILLCELL_X8 FILLER_2_185 ();
 FILLCELL_X1 FILLER_2_193 ();
 FILLCELL_X2 FILLER_2_200 ();
 FILLCELL_X2 FILLER_2_207 ();
 FILLCELL_X2 FILLER_2_215 ();
 FILLCELL_X1 FILLER_2_217 ();
 FILLCELL_X2 FILLER_2_222 ();
 FILLCELL_X1 FILLER_2_224 ();
 FILLCELL_X8 FILLER_2_231 ();
 FILLCELL_X2 FILLER_2_239 ();
 FILLCELL_X1 FILLER_2_241 ();
 FILLCELL_X32 FILLER_2_246 ();
 FILLCELL_X2 FILLER_2_278 ();
 FILLCELL_X32 FILLER_2_297 ();
 FILLCELL_X2 FILLER_2_329 ();
 FILLCELL_X32 FILLER_2_348 ();
 FILLCELL_X32 FILLER_2_380 ();
 FILLCELL_X4 FILLER_2_412 ();
 FILLCELL_X2 FILLER_2_416 ();
 FILLCELL_X1 FILLER_2_418 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X8 FILLER_3_33 ();
 FILLCELL_X1 FILLER_3_41 ();
 FILLCELL_X1 FILLER_3_63 ();
 FILLCELL_X4 FILLER_3_73 ();
 FILLCELL_X1 FILLER_3_77 ();
 FILLCELL_X8 FILLER_3_81 ();
 FILLCELL_X2 FILLER_3_89 ();
 FILLCELL_X4 FILLER_3_110 ();
 FILLCELL_X4 FILLER_3_121 ();
 FILLCELL_X2 FILLER_3_125 ();
 FILLCELL_X16 FILLER_3_146 ();
 FILLCELL_X4 FILLER_3_162 ();
 FILLCELL_X1 FILLER_3_166 ();
 FILLCELL_X2 FILLER_3_173 ();
 FILLCELL_X8 FILLER_3_177 ();
 FILLCELL_X1 FILLER_3_185 ();
 FILLCELL_X4 FILLER_3_195 ();
 FILLCELL_X1 FILLER_3_199 ();
 FILLCELL_X16 FILLER_3_204 ();
 FILLCELL_X8 FILLER_3_220 ();
 FILLCELL_X2 FILLER_3_228 ();
 FILLCELL_X1 FILLER_3_230 ();
 FILLCELL_X16 FILLER_3_248 ();
 FILLCELL_X2 FILLER_3_264 ();
 FILLCELL_X2 FILLER_3_287 ();
 FILLCELL_X16 FILLER_3_312 ();
 FILLCELL_X8 FILLER_3_328 ();
 FILLCELL_X1 FILLER_3_336 ();
 FILLCELL_X2 FILLER_3_340 ();
 FILLCELL_X1 FILLER_3_342 ();
 FILLCELL_X32 FILLER_3_347 ();
 FILLCELL_X32 FILLER_3_379 ();
 FILLCELL_X8 FILLER_3_411 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X16 FILLER_4_33 ();
 FILLCELL_X4 FILLER_4_49 ();
 FILLCELL_X4 FILLER_4_63 ();
 FILLCELL_X2 FILLER_4_67 ();
 FILLCELL_X4 FILLER_4_94 ();
 FILLCELL_X2 FILLER_4_98 ();
 FILLCELL_X2 FILLER_4_103 ();
 FILLCELL_X8 FILLER_4_120 ();
 FILLCELL_X2 FILLER_4_128 ();
 FILLCELL_X1 FILLER_4_130 ();
 FILLCELL_X8 FILLER_4_134 ();
 FILLCELL_X1 FILLER_4_142 ();
 FILLCELL_X4 FILLER_4_149 ();
 FILLCELL_X2 FILLER_4_153 ();
 FILLCELL_X1 FILLER_4_155 ();
 FILLCELL_X1 FILLER_4_178 ();
 FILLCELL_X1 FILLER_4_184 ();
 FILLCELL_X16 FILLER_4_204 ();
 FILLCELL_X4 FILLER_4_220 ();
 FILLCELL_X2 FILLER_4_224 ();
 FILLCELL_X1 FILLER_4_226 ();
 FILLCELL_X32 FILLER_4_230 ();
 FILLCELL_X16 FILLER_4_262 ();
 FILLCELL_X2 FILLER_4_278 ();
 FILLCELL_X1 FILLER_4_280 ();
 FILLCELL_X1 FILLER_4_290 ();
 FILLCELL_X8 FILLER_4_300 ();
 FILLCELL_X1 FILLER_4_308 ();
 FILLCELL_X2 FILLER_4_343 ();
 FILLCELL_X1 FILLER_4_345 ();
 FILLCELL_X32 FILLER_4_367 ();
 FILLCELL_X16 FILLER_4_399 ();
 FILLCELL_X4 FILLER_4_415 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X16 FILLER_5_33 ();
 FILLCELL_X2 FILLER_5_49 ();
 FILLCELL_X1 FILLER_5_54 ();
 FILLCELL_X2 FILLER_5_63 ();
 FILLCELL_X1 FILLER_5_65 ();
 FILLCELL_X4 FILLER_5_80 ();
 FILLCELL_X1 FILLER_5_84 ();
 FILLCELL_X8 FILLER_5_93 ();
 FILLCELL_X4 FILLER_5_101 ();
 FILLCELL_X1 FILLER_5_105 ();
 FILLCELL_X4 FILLER_5_111 ();
 FILLCELL_X1 FILLER_5_115 ();
 FILLCELL_X8 FILLER_5_121 ();
 FILLCELL_X8 FILLER_5_134 ();
 FILLCELL_X4 FILLER_5_163 ();
 FILLCELL_X1 FILLER_5_187 ();
 FILLCELL_X4 FILLER_5_195 ();
 FILLCELL_X8 FILLER_5_205 ();
 FILLCELL_X2 FILLER_5_213 ();
 FILLCELL_X1 FILLER_5_215 ();
 FILLCELL_X2 FILLER_5_224 ();
 FILLCELL_X4 FILLER_5_235 ();
 FILLCELL_X1 FILLER_5_239 ();
 FILLCELL_X16 FILLER_5_248 ();
 FILLCELL_X8 FILLER_5_264 ();
 FILLCELL_X4 FILLER_5_272 ();
 FILLCELL_X1 FILLER_5_276 ();
 FILLCELL_X1 FILLER_5_284 ();
 FILLCELL_X1 FILLER_5_291 ();
 FILLCELL_X16 FILLER_5_296 ();
 FILLCELL_X2 FILLER_5_315 ();
 FILLCELL_X1 FILLER_5_317 ();
 FILLCELL_X2 FILLER_5_321 ();
 FILLCELL_X1 FILLER_5_323 ();
 FILLCELL_X2 FILLER_5_350 ();
 FILLCELL_X32 FILLER_5_364 ();
 FILLCELL_X16 FILLER_5_396 ();
 FILLCELL_X4 FILLER_5_412 ();
 FILLCELL_X2 FILLER_5_416 ();
 FILLCELL_X1 FILLER_5_418 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X2 FILLER_6_9 ();
 FILLCELL_X1 FILLER_6_11 ();
 FILLCELL_X8 FILLER_6_15 ();
 FILLCELL_X2 FILLER_6_23 ();
 FILLCELL_X1 FILLER_6_46 ();
 FILLCELL_X8 FILLER_6_68 ();
 FILLCELL_X4 FILLER_6_76 ();
 FILLCELL_X2 FILLER_6_80 ();
 FILLCELL_X1 FILLER_6_82 ();
 FILLCELL_X16 FILLER_6_100 ();
 FILLCELL_X1 FILLER_6_116 ();
 FILLCELL_X1 FILLER_6_123 ();
 FILLCELL_X4 FILLER_6_157 ();
 FILLCELL_X32 FILLER_6_172 ();
 FILLCELL_X8 FILLER_6_204 ();
 FILLCELL_X32 FILLER_6_231 ();
 FILLCELL_X2 FILLER_6_289 ();
 FILLCELL_X16 FILLER_6_295 ();
 FILLCELL_X4 FILLER_6_317 ();
 FILLCELL_X2 FILLER_6_321 ();
 FILLCELL_X8 FILLER_6_328 ();
 FILLCELL_X2 FILLER_6_336 ();
 FILLCELL_X4 FILLER_6_343 ();
 FILLCELL_X1 FILLER_6_347 ();
 FILLCELL_X1 FILLER_6_355 ();
 FILLCELL_X16 FILLER_6_386 ();
 FILLCELL_X2 FILLER_6_402 ();
 FILLCELL_X1 FILLER_6_404 ();
 FILLCELL_X1 FILLER_6_408 ();
 FILLCELL_X4 FILLER_6_412 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X2 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_46 ();
 FILLCELL_X1 FILLER_7_54 ();
 FILLCELL_X16 FILLER_7_58 ();
 FILLCELL_X8 FILLER_7_74 ();
 FILLCELL_X2 FILLER_7_82 ();
 FILLCELL_X4 FILLER_7_93 ();
 FILLCELL_X1 FILLER_7_97 ();
 FILLCELL_X8 FILLER_7_101 ();
 FILLCELL_X4 FILLER_7_109 ();
 FILLCELL_X2 FILLER_7_113 ();
 FILLCELL_X1 FILLER_7_115 ();
 FILLCELL_X8 FILLER_7_119 ();
 FILLCELL_X2 FILLER_7_127 ();
 FILLCELL_X8 FILLER_7_132 ();
 FILLCELL_X2 FILLER_7_140 ();
 FILLCELL_X1 FILLER_7_147 ();
 FILLCELL_X4 FILLER_7_157 ();
 FILLCELL_X2 FILLER_7_161 ();
 FILLCELL_X1 FILLER_7_163 ();
 FILLCELL_X32 FILLER_7_173 ();
 FILLCELL_X8 FILLER_7_205 ();
 FILLCELL_X4 FILLER_7_235 ();
 FILLCELL_X2 FILLER_7_239 ();
 FILLCELL_X8 FILLER_7_262 ();
 FILLCELL_X4 FILLER_7_270 ();
 FILLCELL_X2 FILLER_7_274 ();
 FILLCELL_X1 FILLER_7_276 ();
 FILLCELL_X1 FILLER_7_292 ();
 FILLCELL_X1 FILLER_7_307 ();
 FILLCELL_X8 FILLER_7_311 ();
 FILLCELL_X4 FILLER_7_325 ();
 FILLCELL_X2 FILLER_7_329 ();
 FILLCELL_X4 FILLER_7_337 ();
 FILLCELL_X16 FILLER_7_363 ();
 FILLCELL_X4 FILLER_7_379 ();
 FILLCELL_X2 FILLER_7_383 ();
 FILLCELL_X1 FILLER_7_385 ();
 FILLCELL_X2 FILLER_7_389 ();
 FILLCELL_X1 FILLER_7_391 ();
 FILLCELL_X2 FILLER_7_395 ();
 FILLCELL_X1 FILLER_7_397 ();
 FILLCELL_X1 FILLER_7_418 ();
 FILLCELL_X4 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_35 ();
 FILLCELL_X16 FILLER_8_48 ();
 FILLCELL_X4 FILLER_8_64 ();
 FILLCELL_X1 FILLER_8_68 ();
 FILLCELL_X8 FILLER_8_78 ();
 FILLCELL_X2 FILLER_8_86 ();
 FILLCELL_X8 FILLER_8_95 ();
 FILLCELL_X4 FILLER_8_103 ();
 FILLCELL_X2 FILLER_8_131 ();
 FILLCELL_X2 FILLER_8_154 ();
 FILLCELL_X4 FILLER_8_161 ();
 FILLCELL_X16 FILLER_8_184 ();
 FILLCELL_X8 FILLER_8_200 ();
 FILLCELL_X8 FILLER_8_225 ();
 FILLCELL_X4 FILLER_8_233 ();
 FILLCELL_X2 FILLER_8_237 ();
 FILLCELL_X1 FILLER_8_239 ();
 FILLCELL_X4 FILLER_8_246 ();
 FILLCELL_X2 FILLER_8_250 ();
 FILLCELL_X8 FILLER_8_255 ();
 FILLCELL_X4 FILLER_8_263 ();
 FILLCELL_X1 FILLER_8_289 ();
 FILLCELL_X8 FILLER_8_301 ();
 FILLCELL_X4 FILLER_8_309 ();
 FILLCELL_X2 FILLER_8_327 ();
 FILLCELL_X1 FILLER_8_375 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X8 FILLER_9_17 ();
 FILLCELL_X2 FILLER_9_25 ();
 FILLCELL_X8 FILLER_9_56 ();
 FILLCELL_X2 FILLER_9_64 ();
 FILLCELL_X1 FILLER_9_75 ();
 FILLCELL_X4 FILLER_9_100 ();
 FILLCELL_X2 FILLER_9_104 ();
 FILLCELL_X4 FILLER_9_119 ();
 FILLCELL_X2 FILLER_9_123 ();
 FILLCELL_X1 FILLER_9_125 ();
 FILLCELL_X8 FILLER_9_145 ();
 FILLCELL_X16 FILLER_9_159 ();
 FILLCELL_X2 FILLER_9_175 ();
 FILLCELL_X4 FILLER_9_198 ();
 FILLCELL_X1 FILLER_9_202 ();
 FILLCELL_X2 FILLER_9_220 ();
 FILLCELL_X1 FILLER_9_222 ();
 FILLCELL_X1 FILLER_9_227 ();
 FILLCELL_X1 FILLER_9_234 ();
 FILLCELL_X16 FILLER_9_254 ();
 FILLCELL_X8 FILLER_9_270 ();
 FILLCELL_X2 FILLER_9_278 ();
 FILLCELL_X8 FILLER_9_302 ();
 FILLCELL_X2 FILLER_9_310 ();
 FILLCELL_X4 FILLER_9_331 ();
 FILLCELL_X4 FILLER_9_366 ();
 FILLCELL_X1 FILLER_9_406 ();
 FILLCELL_X2 FILLER_9_417 ();
 FILLCELL_X2 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_3 ();
 FILLCELL_X4 FILLER_10_7 ();
 FILLCELL_X1 FILLER_10_11 ();
 FILLCELL_X2 FILLER_10_39 ();
 FILLCELL_X4 FILLER_10_59 ();
 FILLCELL_X2 FILLER_10_63 ();
 FILLCELL_X8 FILLER_10_84 ();
 FILLCELL_X16 FILLER_10_101 ();
 FILLCELL_X8 FILLER_10_117 ();
 FILLCELL_X4 FILLER_10_125 ();
 FILLCELL_X8 FILLER_10_132 ();
 FILLCELL_X4 FILLER_10_140 ();
 FILLCELL_X8 FILLER_10_166 ();
 FILLCELL_X4 FILLER_10_174 ();
 FILLCELL_X1 FILLER_10_178 ();
 FILLCELL_X8 FILLER_10_191 ();
 FILLCELL_X1 FILLER_10_199 ();
 FILLCELL_X4 FILLER_10_213 ();
 FILLCELL_X1 FILLER_10_217 ();
 FILLCELL_X1 FILLER_10_222 ();
 FILLCELL_X1 FILLER_10_228 ();
 FILLCELL_X2 FILLER_10_233 ();
 FILLCELL_X2 FILLER_10_248 ();
 FILLCELL_X2 FILLER_10_259 ();
 FILLCELL_X16 FILLER_10_266 ();
 FILLCELL_X8 FILLER_10_282 ();
 FILLCELL_X4 FILLER_10_290 ();
 FILLCELL_X2 FILLER_10_297 ();
 FILLCELL_X1 FILLER_10_299 ();
 FILLCELL_X32 FILLER_10_309 ();
 FILLCELL_X8 FILLER_10_341 ();
 FILLCELL_X2 FILLER_10_349 ();
 FILLCELL_X1 FILLER_10_351 ();
 FILLCELL_X4 FILLER_10_359 ();
 FILLCELL_X4 FILLER_10_388 ();
 FILLCELL_X1 FILLER_10_392 ();
 FILLCELL_X2 FILLER_10_396 ();
 FILLCELL_X1 FILLER_10_398 ();
 FILLCELL_X1 FILLER_10_412 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_9 ();
 FILLCELL_X2 FILLER_11_13 ();
 FILLCELL_X16 FILLER_11_58 ();
 FILLCELL_X8 FILLER_11_77 ();
 FILLCELL_X8 FILLER_11_112 ();
 FILLCELL_X4 FILLER_11_120 ();
 FILLCELL_X1 FILLER_11_124 ();
 FILLCELL_X16 FILLER_11_142 ();
 FILLCELL_X8 FILLER_11_158 ();
 FILLCELL_X4 FILLER_11_166 ();
 FILLCELL_X2 FILLER_11_170 ();
 FILLCELL_X8 FILLER_11_195 ();
 FILLCELL_X2 FILLER_11_203 ();
 FILLCELL_X1 FILLER_11_205 ();
 FILLCELL_X8 FILLER_11_228 ();
 FILLCELL_X1 FILLER_11_236 ();
 FILLCELL_X1 FILLER_11_242 ();
 FILLCELL_X2 FILLER_11_248 ();
 FILLCELL_X2 FILLER_11_270 ();
 FILLCELL_X2 FILLER_11_297 ();
 FILLCELL_X1 FILLER_11_299 ();
 FILLCELL_X4 FILLER_11_319 ();
 FILLCELL_X2 FILLER_11_326 ();
 FILLCELL_X1 FILLER_11_328 ();
 FILLCELL_X4 FILLER_11_353 ();
 FILLCELL_X2 FILLER_11_357 ();
 FILLCELL_X2 FILLER_11_364 ();
 FILLCELL_X1 FILLER_11_366 ();
 FILLCELL_X8 FILLER_11_370 ();
 FILLCELL_X2 FILLER_11_378 ();
 FILLCELL_X1 FILLER_11_380 ();
 FILLCELL_X2 FILLER_11_414 ();
 FILLCELL_X1 FILLER_12_4 ();
 FILLCELL_X1 FILLER_12_8 ();
 FILLCELL_X1 FILLER_12_26 ();
 FILLCELL_X1 FILLER_12_31 ();
 FILLCELL_X4 FILLER_12_36 ();
 FILLCELL_X2 FILLER_12_40 ();
 FILLCELL_X2 FILLER_12_45 ();
 FILLCELL_X1 FILLER_12_47 ();
 FILLCELL_X8 FILLER_12_55 ();
 FILLCELL_X4 FILLER_12_63 ();
 FILLCELL_X2 FILLER_12_67 ();
 FILLCELL_X2 FILLER_12_88 ();
 FILLCELL_X4 FILLER_12_95 ();
 FILLCELL_X4 FILLER_12_103 ();
 FILLCELL_X2 FILLER_12_122 ();
 FILLCELL_X1 FILLER_12_124 ();
 FILLCELL_X4 FILLER_12_137 ();
 FILLCELL_X2 FILLER_12_141 ();
 FILLCELL_X1 FILLER_12_148 ();
 FILLCELL_X1 FILLER_12_153 ();
 FILLCELL_X2 FILLER_12_173 ();
 FILLCELL_X4 FILLER_12_178 ();
 FILLCELL_X2 FILLER_12_185 ();
 FILLCELL_X4 FILLER_12_190 ();
 FILLCELL_X2 FILLER_12_194 ();
 FILLCELL_X2 FILLER_12_239 ();
 FILLCELL_X1 FILLER_12_241 ();
 FILLCELL_X8 FILLER_12_267 ();
 FILLCELL_X2 FILLER_12_275 ();
 FILLCELL_X4 FILLER_12_292 ();
 FILLCELL_X8 FILLER_12_305 ();
 FILLCELL_X4 FILLER_12_313 ();
 FILLCELL_X2 FILLER_12_317 ();
 FILLCELL_X1 FILLER_12_319 ();
 FILLCELL_X8 FILLER_12_371 ();
 FILLCELL_X2 FILLER_12_389 ();
 FILLCELL_X1 FILLER_12_391 ();
 FILLCELL_X1 FILLER_12_415 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_17 ();
 FILLCELL_X2 FILLER_13_21 ();
 FILLCELL_X1 FILLER_13_23 ();
 FILLCELL_X2 FILLER_13_29 ();
 FILLCELL_X2 FILLER_13_45 ();
 FILLCELL_X1 FILLER_13_47 ();
 FILLCELL_X2 FILLER_13_55 ();
 FILLCELL_X8 FILLER_13_60 ();
 FILLCELL_X1 FILLER_13_68 ();
 FILLCELL_X16 FILLER_13_78 ();
 FILLCELL_X2 FILLER_13_94 ();
 FILLCELL_X1 FILLER_13_108 ();
 FILLCELL_X1 FILLER_13_127 ();
 FILLCELL_X1 FILLER_13_131 ();
 FILLCELL_X4 FILLER_13_154 ();
 FILLCELL_X2 FILLER_13_158 ();
 FILLCELL_X2 FILLER_13_188 ();
 FILLCELL_X2 FILLER_13_204 ();
 FILLCELL_X1 FILLER_13_206 ();
 FILLCELL_X4 FILLER_13_212 ();
 FILLCELL_X2 FILLER_13_216 ();
 FILLCELL_X1 FILLER_13_236 ();
 FILLCELL_X1 FILLER_13_242 ();
 FILLCELL_X1 FILLER_13_249 ();
 FILLCELL_X32 FILLER_13_261 ();
 FILLCELL_X2 FILLER_13_293 ();
 FILLCELL_X1 FILLER_13_295 ();
 FILLCELL_X2 FILLER_13_300 ();
 FILLCELL_X1 FILLER_13_302 ();
 FILLCELL_X8 FILLER_13_310 ();
 FILLCELL_X4 FILLER_13_318 ();
 FILLCELL_X2 FILLER_13_322 ();
 FILLCELL_X4 FILLER_13_334 ();
 FILLCELL_X2 FILLER_13_338 ();
 FILLCELL_X1 FILLER_13_343 ();
 FILLCELL_X4 FILLER_13_366 ();
 FILLCELL_X2 FILLER_13_370 ();
 FILLCELL_X4 FILLER_13_375 ();
 FILLCELL_X1 FILLER_13_379 ();
 FILLCELL_X2 FILLER_13_386 ();
 FILLCELL_X8 FILLER_13_397 ();
 FILLCELL_X1 FILLER_13_405 ();
 FILLCELL_X1 FILLER_13_415 ();
 FILLCELL_X16 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_20 ();
 FILLCELL_X2 FILLER_14_39 ();
 FILLCELL_X1 FILLER_14_104 ();
 FILLCELL_X4 FILLER_14_109 ();
 FILLCELL_X2 FILLER_14_113 ();
 FILLCELL_X1 FILLER_14_127 ();
 FILLCELL_X2 FILLER_14_132 ();
 FILLCELL_X1 FILLER_14_134 ();
 FILLCELL_X8 FILLER_14_138 ();
 FILLCELL_X4 FILLER_14_146 ();
 FILLCELL_X2 FILLER_14_156 ();
 FILLCELL_X4 FILLER_14_163 ();
 FILLCELL_X4 FILLER_14_171 ();
 FILLCELL_X2 FILLER_14_175 ();
 FILLCELL_X1 FILLER_14_186 ();
 FILLCELL_X8 FILLER_14_195 ();
 FILLCELL_X2 FILLER_14_203 ();
 FILLCELL_X1 FILLER_14_205 ();
 FILLCELL_X1 FILLER_14_240 ();
 FILLCELL_X2 FILLER_14_247 ();
 FILLCELL_X1 FILLER_14_252 ();
 FILLCELL_X1 FILLER_14_287 ();
 FILLCELL_X2 FILLER_14_299 ();
 FILLCELL_X8 FILLER_14_309 ();
 FILLCELL_X4 FILLER_14_317 ();
 FILLCELL_X2 FILLER_14_321 ();
 FILLCELL_X1 FILLER_14_323 ();
 FILLCELL_X2 FILLER_14_371 ();
 FILLCELL_X1 FILLER_14_373 ();
 FILLCELL_X2 FILLER_14_391 ();
 FILLCELL_X2 FILLER_14_401 ();
 FILLCELL_X1 FILLER_14_403 ();
 FILLCELL_X2 FILLER_14_407 ();
 FILLCELL_X1 FILLER_14_412 ();
 FILLCELL_X4 FILLER_15_39 ();
 FILLCELL_X1 FILLER_15_43 ();
 FILLCELL_X2 FILLER_15_49 ();
 FILLCELL_X1 FILLER_15_73 ();
 FILLCELL_X1 FILLER_15_88 ();
 FILLCELL_X4 FILLER_15_111 ();
 FILLCELL_X16 FILLER_15_123 ();
 FILLCELL_X8 FILLER_15_139 ();
 FILLCELL_X4 FILLER_15_147 ();
 FILLCELL_X2 FILLER_15_151 ();
 FILLCELL_X1 FILLER_15_162 ();
 FILLCELL_X1 FILLER_15_173 ();
 FILLCELL_X4 FILLER_15_178 ();
 FILLCELL_X2 FILLER_15_182 ();
 FILLCELL_X1 FILLER_15_184 ();
 FILLCELL_X16 FILLER_15_197 ();
 FILLCELL_X2 FILLER_15_213 ();
 FILLCELL_X4 FILLER_15_220 ();
 FILLCELL_X4 FILLER_15_237 ();
 FILLCELL_X4 FILLER_15_260 ();
 FILLCELL_X2 FILLER_15_264 ();
 FILLCELL_X1 FILLER_15_266 ();
 FILLCELL_X1 FILLER_15_280 ();
 FILLCELL_X32 FILLER_15_315 ();
 FILLCELL_X8 FILLER_15_347 ();
 FILLCELL_X1 FILLER_15_355 ();
 FILLCELL_X4 FILLER_15_376 ();
 FILLCELL_X1 FILLER_15_380 ();
 FILLCELL_X1 FILLER_15_397 ();
 FILLCELL_X1 FILLER_15_418 ();
 FILLCELL_X4 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_11 ();
 FILLCELL_X1 FILLER_16_13 ();
 FILLCELL_X1 FILLER_16_17 ();
 FILLCELL_X1 FILLER_16_24 ();
 FILLCELL_X1 FILLER_16_77 ();
 FILLCELL_X8 FILLER_16_85 ();
 FILLCELL_X2 FILLER_16_116 ();
 FILLCELL_X2 FILLER_16_126 ();
 FILLCELL_X16 FILLER_16_131 ();
 FILLCELL_X1 FILLER_16_147 ();
 FILLCELL_X1 FILLER_16_167 ();
 FILLCELL_X1 FILLER_16_172 ();
 FILLCELL_X1 FILLER_16_176 ();
 FILLCELL_X2 FILLER_16_180 ();
 FILLCELL_X1 FILLER_16_199 ();
 FILLCELL_X8 FILLER_16_203 ();
 FILLCELL_X4 FILLER_16_211 ();
 FILLCELL_X2 FILLER_16_221 ();
 FILLCELL_X1 FILLER_16_223 ();
 FILLCELL_X4 FILLER_16_243 ();
 FILLCELL_X2 FILLER_16_250 ();
 FILLCELL_X1 FILLER_16_252 ();
 FILLCELL_X16 FILLER_16_263 ();
 FILLCELL_X8 FILLER_16_288 ();
 FILLCELL_X1 FILLER_16_296 ();
 FILLCELL_X2 FILLER_16_311 ();
 FILLCELL_X1 FILLER_16_317 ();
 FILLCELL_X4 FILLER_16_346 ();
 FILLCELL_X1 FILLER_16_350 ();
 FILLCELL_X16 FILLER_16_361 ();
 FILLCELL_X4 FILLER_16_377 ();
 FILLCELL_X2 FILLER_16_381 ();
 FILLCELL_X1 FILLER_16_398 ();
 FILLCELL_X2 FILLER_16_413 ();
 FILLCELL_X1 FILLER_16_418 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_5 ();
 FILLCELL_X2 FILLER_17_30 ();
 FILLCELL_X1 FILLER_17_32 ();
 FILLCELL_X1 FILLER_17_55 ();
 FILLCELL_X4 FILLER_17_60 ();
 FILLCELL_X2 FILLER_17_64 ();
 FILLCELL_X1 FILLER_17_66 ();
 FILLCELL_X8 FILLER_17_71 ();
 FILLCELL_X2 FILLER_17_79 ();
 FILLCELL_X1 FILLER_17_81 ();
 FILLCELL_X4 FILLER_17_89 ();
 FILLCELL_X2 FILLER_17_93 ();
 FILLCELL_X8 FILLER_17_103 ();
 FILLCELL_X4 FILLER_17_111 ();
 FILLCELL_X2 FILLER_17_115 ();
 FILLCELL_X1 FILLER_17_153 ();
 FILLCELL_X8 FILLER_17_159 ();
 FILLCELL_X2 FILLER_17_167 ();
 FILLCELL_X1 FILLER_17_172 ();
 FILLCELL_X2 FILLER_17_177 ();
 FILLCELL_X1 FILLER_17_179 ();
 FILLCELL_X2 FILLER_17_187 ();
 FILLCELL_X1 FILLER_17_189 ();
 FILLCELL_X8 FILLER_17_194 ();
 FILLCELL_X1 FILLER_17_202 ();
 FILLCELL_X8 FILLER_17_230 ();
 FILLCELL_X4 FILLER_17_238 ();
 FILLCELL_X2 FILLER_17_242 ();
 FILLCELL_X1 FILLER_17_244 ();
 FILLCELL_X8 FILLER_17_274 ();
 FILLCELL_X1 FILLER_17_282 ();
 FILLCELL_X16 FILLER_17_313 ();
 FILLCELL_X2 FILLER_17_329 ();
 FILLCELL_X2 FILLER_17_352 ();
 FILLCELL_X2 FILLER_17_358 ();
 FILLCELL_X1 FILLER_17_360 ();
 FILLCELL_X2 FILLER_17_365 ();
 FILLCELL_X2 FILLER_17_371 ();
 FILLCELL_X1 FILLER_17_377 ();
 FILLCELL_X2 FILLER_17_382 ();
 FILLCELL_X2 FILLER_17_394 ();
 FILLCELL_X1 FILLER_17_401 ();
 FILLCELL_X8 FILLER_18_36 ();
 FILLCELL_X2 FILLER_18_44 ();
 FILLCELL_X1 FILLER_18_46 ();
 FILLCELL_X4 FILLER_18_60 ();
 FILLCELL_X4 FILLER_18_68 ();
 FILLCELL_X4 FILLER_18_95 ();
 FILLCELL_X1 FILLER_18_99 ();
 FILLCELL_X1 FILLER_18_104 ();
 FILLCELL_X2 FILLER_18_119 ();
 FILLCELL_X1 FILLER_18_121 ();
 FILLCELL_X8 FILLER_18_127 ();
 FILLCELL_X2 FILLER_18_145 ();
 FILLCELL_X2 FILLER_18_151 ();
 FILLCELL_X1 FILLER_18_153 ();
 FILLCELL_X1 FILLER_18_158 ();
 FILLCELL_X2 FILLER_18_163 ();
 FILLCELL_X1 FILLER_18_165 ();
 FILLCELL_X2 FILLER_18_179 ();
 FILLCELL_X16 FILLER_18_184 ();
 FILLCELL_X8 FILLER_18_200 ();
 FILLCELL_X2 FILLER_18_208 ();
 FILLCELL_X1 FILLER_18_210 ();
 FILLCELL_X2 FILLER_18_216 ();
 FILLCELL_X4 FILLER_18_223 ();
 FILLCELL_X2 FILLER_18_227 ();
 FILLCELL_X2 FILLER_18_265 ();
 FILLCELL_X1 FILLER_18_267 ();
 FILLCELL_X8 FILLER_18_271 ();
 FILLCELL_X16 FILLER_18_300 ();
 FILLCELL_X4 FILLER_18_316 ();
 FILLCELL_X2 FILLER_18_320 ();
 FILLCELL_X1 FILLER_18_322 ();
 FILLCELL_X2 FILLER_18_327 ();
 FILLCELL_X1 FILLER_18_329 ();
 FILLCELL_X8 FILLER_18_334 ();
 FILLCELL_X2 FILLER_18_342 ();
 FILLCELL_X1 FILLER_18_348 ();
 FILLCELL_X2 FILLER_18_368 ();
 FILLCELL_X2 FILLER_18_381 ();
 FILLCELL_X2 FILLER_18_391 ();
 FILLCELL_X1 FILLER_18_393 ();
 FILLCELL_X2 FILLER_18_417 ();
 FILLCELL_X2 FILLER_19_4 ();
 FILLCELL_X1 FILLER_19_9 ();
 FILLCELL_X4 FILLER_19_13 ();
 FILLCELL_X1 FILLER_19_17 ();
 FILLCELL_X4 FILLER_19_58 ();
 FILLCELL_X1 FILLER_19_62 ();
 FILLCELL_X8 FILLER_19_70 ();
 FILLCELL_X1 FILLER_19_78 ();
 FILLCELL_X8 FILLER_19_86 ();
 FILLCELL_X1 FILLER_19_116 ();
 FILLCELL_X8 FILLER_19_121 ();
 FILLCELL_X1 FILLER_19_143 ();
 FILLCELL_X1 FILLER_19_151 ();
 FILLCELL_X1 FILLER_19_156 ();
 FILLCELL_X1 FILLER_19_164 ();
 FILLCELL_X8 FILLER_19_169 ();
 FILLCELL_X2 FILLER_19_177 ();
 FILLCELL_X4 FILLER_19_217 ();
 FILLCELL_X2 FILLER_19_221 ();
 FILLCELL_X1 FILLER_19_223 ();
 FILLCELL_X8 FILLER_19_270 ();
 FILLCELL_X4 FILLER_19_278 ();
 FILLCELL_X1 FILLER_19_282 ();
 FILLCELL_X4 FILLER_19_290 ();
 FILLCELL_X1 FILLER_19_294 ();
 FILLCELL_X4 FILLER_19_302 ();
 FILLCELL_X1 FILLER_19_332 ();
 FILLCELL_X4 FILLER_19_345 ();
 FILLCELL_X1 FILLER_19_349 ();
 FILLCELL_X1 FILLER_19_354 ();
 FILLCELL_X2 FILLER_19_360 ();
 FILLCELL_X1 FILLER_19_362 ();
 FILLCELL_X1 FILLER_19_382 ();
 FILLCELL_X2 FILLER_19_398 ();
 FILLCELL_X2 FILLER_19_417 ();
 FILLCELL_X4 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_5 ();
 FILLCELL_X1 FILLER_20_7 ();
 FILLCELL_X4 FILLER_20_11 ();
 FILLCELL_X2 FILLER_20_30 ();
 FILLCELL_X8 FILLER_20_35 ();
 FILLCELL_X1 FILLER_20_43 ();
 FILLCELL_X1 FILLER_20_55 ();
 FILLCELL_X8 FILLER_20_67 ();
 FILLCELL_X4 FILLER_20_75 ();
 FILLCELL_X1 FILLER_20_79 ();
 FILLCELL_X1 FILLER_20_84 ();
 FILLCELL_X1 FILLER_20_104 ();
 FILLCELL_X16 FILLER_20_108 ();
 FILLCELL_X2 FILLER_20_124 ();
 FILLCELL_X1 FILLER_20_126 ();
 FILLCELL_X1 FILLER_20_146 ();
 FILLCELL_X2 FILLER_20_154 ();
 FILLCELL_X32 FILLER_20_164 ();
 FILLCELL_X4 FILLER_20_196 ();
 FILLCELL_X16 FILLER_20_216 ();
 FILLCELL_X2 FILLER_20_235 ();
 FILLCELL_X4 FILLER_20_248 ();
 FILLCELL_X1 FILLER_20_252 ();
 FILLCELL_X2 FILLER_20_258 ();
 FILLCELL_X4 FILLER_20_270 ();
 FILLCELL_X4 FILLER_20_283 ();
 FILLCELL_X1 FILLER_20_306 ();
 FILLCELL_X4 FILLER_20_312 ();
 FILLCELL_X2 FILLER_20_316 ();
 FILLCELL_X4 FILLER_20_337 ();
 FILLCELL_X1 FILLER_20_341 ();
 FILLCELL_X2 FILLER_20_380 ();
 FILLCELL_X16 FILLER_20_402 ();
 FILLCELL_X1 FILLER_20_418 ();
 FILLCELL_X2 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_6 ();
 FILLCELL_X2 FILLER_21_14 ();
 FILLCELL_X1 FILLER_21_16 ();
 FILLCELL_X1 FILLER_21_26 ();
 FILLCELL_X2 FILLER_21_36 ();
 FILLCELL_X2 FILLER_21_43 ();
 FILLCELL_X1 FILLER_21_45 ();
 FILLCELL_X4 FILLER_21_65 ();
 FILLCELL_X2 FILLER_21_69 ();
 FILLCELL_X8 FILLER_21_80 ();
 FILLCELL_X8 FILLER_21_98 ();
 FILLCELL_X2 FILLER_21_106 ();
 FILLCELL_X1 FILLER_21_108 ();
 FILLCELL_X1 FILLER_21_117 ();
 FILLCELL_X8 FILLER_21_123 ();
 FILLCELL_X2 FILLER_21_131 ();
 FILLCELL_X1 FILLER_21_133 ();
 FILLCELL_X2 FILLER_21_138 ();
 FILLCELL_X1 FILLER_21_140 ();
 FILLCELL_X8 FILLER_21_158 ();
 FILLCELL_X2 FILLER_21_166 ();
 FILLCELL_X32 FILLER_21_173 ();
 FILLCELL_X4 FILLER_21_205 ();
 FILLCELL_X1 FILLER_21_209 ();
 FILLCELL_X8 FILLER_21_229 ();
 FILLCELL_X4 FILLER_21_237 ();
 FILLCELL_X4 FILLER_21_245 ();
 FILLCELL_X1 FILLER_21_249 ();
 FILLCELL_X2 FILLER_21_263 ();
 FILLCELL_X2 FILLER_21_271 ();
 FILLCELL_X4 FILLER_21_282 ();
 FILLCELL_X2 FILLER_21_315 ();
 FILLCELL_X1 FILLER_21_317 ();
 FILLCELL_X1 FILLER_21_327 ();
 FILLCELL_X4 FILLER_21_331 ();
 FILLCELL_X1 FILLER_21_335 ();
 FILLCELL_X1 FILLER_21_338 ();
 FILLCELL_X4 FILLER_21_352 ();
 FILLCELL_X4 FILLER_21_358 ();
 FILLCELL_X2 FILLER_21_362 ();
 FILLCELL_X1 FILLER_21_364 ();
 FILLCELL_X2 FILLER_21_414 ();
 FILLCELL_X2 FILLER_22_1 ();
 FILLCELL_X1 FILLER_22_3 ();
 FILLCELL_X4 FILLER_22_14 ();
 FILLCELL_X1 FILLER_22_48 ();
 FILLCELL_X8 FILLER_22_59 ();
 FILLCELL_X4 FILLER_22_67 ();
 FILLCELL_X2 FILLER_22_71 ();
 FILLCELL_X4 FILLER_22_109 ();
 FILLCELL_X2 FILLER_22_113 ();
 FILLCELL_X8 FILLER_22_120 ();
 FILLCELL_X4 FILLER_22_145 ();
 FILLCELL_X2 FILLER_22_149 ();
 FILLCELL_X1 FILLER_22_151 ();
 FILLCELL_X16 FILLER_22_156 ();
 FILLCELL_X8 FILLER_22_172 ();
 FILLCELL_X2 FILLER_22_180 ();
 FILLCELL_X1 FILLER_22_182 ();
 FILLCELL_X8 FILLER_22_210 ();
 FILLCELL_X2 FILLER_22_218 ();
 FILLCELL_X1 FILLER_22_220 ();
 FILLCELL_X1 FILLER_22_230 ();
 FILLCELL_X4 FILLER_22_234 ();
 FILLCELL_X1 FILLER_22_238 ();
 FILLCELL_X2 FILLER_22_246 ();
 FILLCELL_X1 FILLER_22_248 ();
 FILLCELL_X1 FILLER_22_254 ();
 FILLCELL_X4 FILLER_22_258 ();
 FILLCELL_X2 FILLER_22_262 ();
 FILLCELL_X4 FILLER_22_267 ();
 FILLCELL_X2 FILLER_22_274 ();
 FILLCELL_X16 FILLER_22_287 ();
 FILLCELL_X16 FILLER_22_305 ();
 FILLCELL_X8 FILLER_22_321 ();
 FILLCELL_X8 FILLER_22_340 ();
 FILLCELL_X1 FILLER_22_376 ();
 FILLCELL_X1 FILLER_22_396 ();
 FILLCELL_X2 FILLER_22_403 ();
 FILLCELL_X1 FILLER_22_405 ();
 FILLCELL_X2 FILLER_22_411 ();
 FILLCELL_X2 FILLER_22_416 ();
 FILLCELL_X1 FILLER_22_418 ();
 FILLCELL_X2 FILLER_23_4 ();
 FILLCELL_X1 FILLER_23_33 ();
 FILLCELL_X2 FILLER_23_40 ();
 FILLCELL_X1 FILLER_23_42 ();
 FILLCELL_X16 FILLER_23_55 ();
 FILLCELL_X4 FILLER_23_71 ();
 FILLCELL_X2 FILLER_23_75 ();
 FILLCELL_X1 FILLER_23_77 ();
 FILLCELL_X4 FILLER_23_81 ();
 FILLCELL_X4 FILLER_23_90 ();
 FILLCELL_X1 FILLER_23_94 ();
 FILLCELL_X4 FILLER_23_98 ();
 FILLCELL_X2 FILLER_23_102 ();
 FILLCELL_X1 FILLER_23_104 ();
 FILLCELL_X4 FILLER_23_127 ();
 FILLCELL_X2 FILLER_23_131 ();
 FILLCELL_X8 FILLER_23_136 ();
 FILLCELL_X2 FILLER_23_144 ();
 FILLCELL_X32 FILLER_23_160 ();
 FILLCELL_X4 FILLER_23_192 ();
 FILLCELL_X2 FILLER_23_196 ();
 FILLCELL_X1 FILLER_23_198 ();
 FILLCELL_X2 FILLER_23_212 ();
 FILLCELL_X2 FILLER_23_222 ();
 FILLCELL_X2 FILLER_23_231 ();
 FILLCELL_X2 FILLER_23_238 ();
 FILLCELL_X1 FILLER_23_240 ();
 FILLCELL_X16 FILLER_23_247 ();
 FILLCELL_X1 FILLER_23_263 ();
 FILLCELL_X1 FILLER_23_274 ();
 FILLCELL_X2 FILLER_23_283 ();
 FILLCELL_X1 FILLER_23_290 ();
 FILLCELL_X2 FILLER_23_295 ();
 FILLCELL_X1 FILLER_23_297 ();
 FILLCELL_X8 FILLER_23_302 ();
 FILLCELL_X2 FILLER_23_313 ();
 FILLCELL_X8 FILLER_23_365 ();
 FILLCELL_X4 FILLER_23_373 ();
 FILLCELL_X1 FILLER_23_377 ();
 FILLCELL_X2 FILLER_23_398 ();
 FILLCELL_X1 FILLER_23_400 ();
 FILLCELL_X4 FILLER_23_407 ();
 FILLCELL_X1 FILLER_23_411 ();
 FILLCELL_X1 FILLER_23_415 ();
 FILLCELL_X8 FILLER_24_4 ();
 FILLCELL_X4 FILLER_24_12 ();
 FILLCELL_X2 FILLER_24_16 ();
 FILLCELL_X1 FILLER_24_18 ();
 FILLCELL_X4 FILLER_24_42 ();
 FILLCELL_X1 FILLER_24_84 ();
 FILLCELL_X2 FILLER_24_104 ();
 FILLCELL_X1 FILLER_24_145 ();
 FILLCELL_X16 FILLER_24_176 ();
 FILLCELL_X8 FILLER_24_192 ();
 FILLCELL_X1 FILLER_24_200 ();
 FILLCELL_X2 FILLER_24_221 ();
 FILLCELL_X1 FILLER_24_223 ();
 FILLCELL_X1 FILLER_24_227 ();
 FILLCELL_X4 FILLER_24_233 ();
 FILLCELL_X2 FILLER_24_267 ();
 FILLCELL_X2 FILLER_24_275 ();
 FILLCELL_X1 FILLER_24_277 ();
 FILLCELL_X2 FILLER_24_281 ();
 FILLCELL_X1 FILLER_24_283 ();
 FILLCELL_X2 FILLER_24_301 ();
 FILLCELL_X1 FILLER_24_303 ();
 FILLCELL_X2 FILLER_24_326 ();
 FILLCELL_X1 FILLER_24_328 ();
 FILLCELL_X2 FILLER_24_335 ();
 FILLCELL_X1 FILLER_24_343 ();
 FILLCELL_X2 FILLER_24_347 ();
 FILLCELL_X16 FILLER_24_352 ();
 FILLCELL_X8 FILLER_24_368 ();
 FILLCELL_X2 FILLER_24_376 ();
 FILLCELL_X1 FILLER_24_378 ();
 FILLCELL_X1 FILLER_24_390 ();
 FILLCELL_X2 FILLER_24_417 ();
 FILLCELL_X16 FILLER_25_1 ();
 FILLCELL_X4 FILLER_25_17 ();
 FILLCELL_X1 FILLER_25_21 ();
 FILLCELL_X8 FILLER_25_25 ();
 FILLCELL_X2 FILLER_25_33 ();
 FILLCELL_X8 FILLER_25_40 ();
 FILLCELL_X4 FILLER_25_48 ();
 FILLCELL_X4 FILLER_25_69 ();
 FILLCELL_X2 FILLER_25_73 ();
 FILLCELL_X1 FILLER_25_101 ();
 FILLCELL_X4 FILLER_25_130 ();
 FILLCELL_X2 FILLER_25_141 ();
 FILLCELL_X2 FILLER_25_161 ();
 FILLCELL_X8 FILLER_25_166 ();
 FILLCELL_X8 FILLER_25_185 ();
 FILLCELL_X4 FILLER_25_193 ();
 FILLCELL_X2 FILLER_25_197 ();
 FILLCELL_X1 FILLER_25_199 ();
 FILLCELL_X8 FILLER_25_203 ();
 FILLCELL_X4 FILLER_25_217 ();
 FILLCELL_X2 FILLER_25_231 ();
 FILLCELL_X1 FILLER_25_233 ();
 FILLCELL_X2 FILLER_25_242 ();
 FILLCELL_X16 FILLER_25_248 ();
 FILLCELL_X4 FILLER_25_264 ();
 FILLCELL_X1 FILLER_25_268 ();
 FILLCELL_X8 FILLER_25_298 ();
 FILLCELL_X1 FILLER_25_306 ();
 FILLCELL_X8 FILLER_25_311 ();
 FILLCELL_X1 FILLER_25_319 ();
 FILLCELL_X2 FILLER_25_359 ();
 FILLCELL_X4 FILLER_25_372 ();
 FILLCELL_X2 FILLER_25_376 ();
 FILLCELL_X1 FILLER_25_378 ();
 FILLCELL_X2 FILLER_25_414 ();
 FILLCELL_X2 FILLER_26_1 ();
 FILLCELL_X4 FILLER_26_30 ();
 FILLCELL_X1 FILLER_26_54 ();
 FILLCELL_X4 FILLER_26_67 ();
 FILLCELL_X16 FILLER_26_75 ();
 FILLCELL_X8 FILLER_26_91 ();
 FILLCELL_X1 FILLER_26_99 ();
 FILLCELL_X1 FILLER_26_104 ();
 FILLCELL_X1 FILLER_26_109 ();
 FILLCELL_X1 FILLER_26_116 ();
 FILLCELL_X1 FILLER_26_121 ();
 FILLCELL_X8 FILLER_26_129 ();
 FILLCELL_X4 FILLER_26_141 ();
 FILLCELL_X2 FILLER_26_145 ();
 FILLCELL_X2 FILLER_26_153 ();
 FILLCELL_X8 FILLER_26_163 ();
 FILLCELL_X2 FILLER_26_171 ();
 FILLCELL_X1 FILLER_26_173 ();
 FILLCELL_X8 FILLER_26_185 ();
 FILLCELL_X2 FILLER_26_193 ();
 FILLCELL_X1 FILLER_26_195 ();
 FILLCELL_X4 FILLER_26_215 ();
 FILLCELL_X2 FILLER_26_219 ();
 FILLCELL_X1 FILLER_26_228 ();
 FILLCELL_X2 FILLER_26_232 ();
 FILLCELL_X1 FILLER_26_234 ();
 FILLCELL_X1 FILLER_26_240 ();
 FILLCELL_X8 FILLER_26_249 ();
 FILLCELL_X2 FILLER_26_257 ();
 FILLCELL_X1 FILLER_26_262 ();
 FILLCELL_X8 FILLER_26_267 ();
 FILLCELL_X2 FILLER_26_280 ();
 FILLCELL_X1 FILLER_26_282 ();
 FILLCELL_X16 FILLER_26_286 ();
 FILLCELL_X4 FILLER_26_302 ();
 FILLCELL_X1 FILLER_26_306 ();
 FILLCELL_X8 FILLER_26_311 ();
 FILLCELL_X4 FILLER_26_319 ();
 FILLCELL_X2 FILLER_26_323 ();
 FILLCELL_X1 FILLER_26_325 ();
 FILLCELL_X1 FILLER_26_339 ();
 FILLCELL_X2 FILLER_26_343 ();
 FILLCELL_X1 FILLER_26_377 ();
 FILLCELL_X2 FILLER_26_407 ();
 FILLCELL_X4 FILLER_27_7 ();
 FILLCELL_X2 FILLER_27_11 ();
 FILLCELL_X1 FILLER_27_13 ();
 FILLCELL_X16 FILLER_27_53 ();
 FILLCELL_X4 FILLER_27_69 ();
 FILLCELL_X2 FILLER_27_73 ();
 FILLCELL_X1 FILLER_27_75 ();
 FILLCELL_X4 FILLER_27_79 ();
 FILLCELL_X2 FILLER_27_83 ();
 FILLCELL_X1 FILLER_27_91 ();
 FILLCELL_X8 FILLER_27_96 ();
 FILLCELL_X1 FILLER_27_119 ();
 FILLCELL_X16 FILLER_27_141 ();
 FILLCELL_X16 FILLER_27_174 ();
 FILLCELL_X8 FILLER_27_190 ();
 FILLCELL_X2 FILLER_27_211 ();
 FILLCELL_X1 FILLER_27_220 ();
 FILLCELL_X2 FILLER_27_224 ();
 FILLCELL_X8 FILLER_27_231 ();
 FILLCELL_X4 FILLER_27_239 ();
 FILLCELL_X2 FILLER_27_243 ();
 FILLCELL_X1 FILLER_27_245 ();
 FILLCELL_X2 FILLER_27_266 ();
 FILLCELL_X8 FILLER_27_285 ();
 FILLCELL_X4 FILLER_27_293 ();
 FILLCELL_X1 FILLER_27_297 ();
 FILLCELL_X4 FILLER_27_319 ();
 FILLCELL_X2 FILLER_27_323 ();
 FILLCELL_X2 FILLER_27_334 ();
 FILLCELL_X16 FILLER_27_342 ();
 FILLCELL_X8 FILLER_27_358 ();
 FILLCELL_X1 FILLER_27_366 ();
 FILLCELL_X2 FILLER_27_390 ();
 FILLCELL_X8 FILLER_28_1 ();
 FILLCELL_X2 FILLER_28_9 ();
 FILLCELL_X1 FILLER_28_11 ();
 FILLCELL_X2 FILLER_28_22 ();
 FILLCELL_X2 FILLER_28_42 ();
 FILLCELL_X1 FILLER_28_44 ();
 FILLCELL_X4 FILLER_28_48 ();
 FILLCELL_X1 FILLER_28_52 ();
 FILLCELL_X1 FILLER_28_103 ();
 FILLCELL_X2 FILLER_28_115 ();
 FILLCELL_X2 FILLER_28_124 ();
 FILLCELL_X4 FILLER_28_130 ();
 FILLCELL_X2 FILLER_28_134 ();
 FILLCELL_X4 FILLER_28_142 ();
 FILLCELL_X2 FILLER_28_146 ();
 FILLCELL_X1 FILLER_28_148 ();
 FILLCELL_X8 FILLER_28_181 ();
 FILLCELL_X1 FILLER_28_189 ();
 FILLCELL_X8 FILLER_28_234 ();
 FILLCELL_X2 FILLER_28_242 ();
 FILLCELL_X1 FILLER_28_244 ();
 FILLCELL_X8 FILLER_28_258 ();
 FILLCELL_X4 FILLER_28_266 ();
 FILLCELL_X1 FILLER_28_270 ();
 FILLCELL_X8 FILLER_28_273 ();
 FILLCELL_X1 FILLER_28_281 ();
 FILLCELL_X8 FILLER_28_286 ();
 FILLCELL_X4 FILLER_28_294 ();
 FILLCELL_X1 FILLER_28_318 ();
 FILLCELL_X4 FILLER_28_336 ();
 FILLCELL_X4 FILLER_28_347 ();
 FILLCELL_X2 FILLER_28_351 ();
 FILLCELL_X8 FILLER_28_357 ();
 FILLCELL_X4 FILLER_28_365 ();
 FILLCELL_X2 FILLER_28_375 ();
 FILLCELL_X2 FILLER_28_399 ();
 FILLCELL_X1 FILLER_28_418 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X4 FILLER_29_9 ();
 FILLCELL_X1 FILLER_29_13 ();
 FILLCELL_X1 FILLER_29_32 ();
 FILLCELL_X1 FILLER_29_38 ();
 FILLCELL_X2 FILLER_29_43 ();
 FILLCELL_X2 FILLER_29_52 ();
 FILLCELL_X4 FILLER_29_71 ();
 FILLCELL_X2 FILLER_29_75 ();
 FILLCELL_X1 FILLER_29_77 ();
 FILLCELL_X2 FILLER_29_82 ();
 FILLCELL_X1 FILLER_29_84 ();
 FILLCELL_X2 FILLER_29_91 ();
 FILLCELL_X2 FILLER_29_105 ();
 FILLCELL_X2 FILLER_29_111 ();
 FILLCELL_X1 FILLER_29_113 ();
 FILLCELL_X1 FILLER_29_125 ();
 FILLCELL_X1 FILLER_29_130 ();
 FILLCELL_X2 FILLER_29_155 ();
 FILLCELL_X16 FILLER_29_181 ();
 FILLCELL_X8 FILLER_29_197 ();
 FILLCELL_X4 FILLER_29_205 ();
 FILLCELL_X2 FILLER_29_209 ();
 FILLCELL_X1 FILLER_29_224 ();
 FILLCELL_X1 FILLER_29_228 ();
 FILLCELL_X2 FILLER_29_234 ();
 FILLCELL_X1 FILLER_29_254 ();
 FILLCELL_X2 FILLER_29_262 ();
 FILLCELL_X1 FILLER_29_273 ();
 FILLCELL_X4 FILLER_29_299 ();
 FILLCELL_X2 FILLER_29_303 ();
 FILLCELL_X1 FILLER_29_305 ();
 FILLCELL_X1 FILLER_29_328 ();
 FILLCELL_X1 FILLER_29_336 ();
 FILLCELL_X8 FILLER_29_341 ();
 FILLCELL_X2 FILLER_29_349 ();
 FILLCELL_X2 FILLER_29_357 ();
 FILLCELL_X4 FILLER_29_380 ();
 FILLCELL_X2 FILLER_29_384 ();
 FILLCELL_X1 FILLER_29_386 ();
 FILLCELL_X4 FILLER_29_390 ();
 FILLCELL_X2 FILLER_29_394 ();
 FILLCELL_X1 FILLER_29_396 ();
 FILLCELL_X8 FILLER_29_403 ();
 FILLCELL_X2 FILLER_29_411 ();
 FILLCELL_X2 FILLER_30_1 ();
 FILLCELL_X1 FILLER_30_27 ();
 FILLCELL_X2 FILLER_30_37 ();
 FILLCELL_X2 FILLER_30_43 ();
 FILLCELL_X8 FILLER_30_50 ();
 FILLCELL_X2 FILLER_30_58 ();
 FILLCELL_X1 FILLER_30_93 ();
 FILLCELL_X1 FILLER_30_98 ();
 FILLCELL_X1 FILLER_30_104 ();
 FILLCELL_X4 FILLER_30_112 ();
 FILLCELL_X2 FILLER_30_116 ();
 FILLCELL_X1 FILLER_30_118 ();
 FILLCELL_X4 FILLER_30_126 ();
 FILLCELL_X2 FILLER_30_130 ();
 FILLCELL_X8 FILLER_30_139 ();
 FILLCELL_X4 FILLER_30_147 ();
 FILLCELL_X1 FILLER_30_151 ();
 FILLCELL_X1 FILLER_30_159 ();
 FILLCELL_X32 FILLER_30_163 ();
 FILLCELL_X16 FILLER_30_195 ();
 FILLCELL_X8 FILLER_30_211 ();
 FILLCELL_X2 FILLER_30_219 ();
 FILLCELL_X8 FILLER_30_224 ();
 FILLCELL_X2 FILLER_30_232 ();
 FILLCELL_X1 FILLER_30_252 ();
 FILLCELL_X2 FILLER_30_269 ();
 FILLCELL_X1 FILLER_30_271 ();
 FILLCELL_X1 FILLER_30_276 ();
 FILLCELL_X16 FILLER_30_296 ();
 FILLCELL_X2 FILLER_30_312 ();
 FILLCELL_X1 FILLER_30_314 ();
 FILLCELL_X8 FILLER_30_317 ();
 FILLCELL_X4 FILLER_30_325 ();
 FILLCELL_X1 FILLER_30_329 ();
 FILLCELL_X16 FILLER_30_360 ();
 FILLCELL_X4 FILLER_30_376 ();
 FILLCELL_X1 FILLER_30_380 ();
 FILLCELL_X1 FILLER_30_388 ();
 FILLCELL_X8 FILLER_30_406 ();
 FILLCELL_X4 FILLER_30_414 ();
 FILLCELL_X1 FILLER_30_418 ();
 FILLCELL_X8 FILLER_31_28 ();
 FILLCELL_X2 FILLER_31_36 ();
 FILLCELL_X1 FILLER_31_38 ();
 FILLCELL_X1 FILLER_31_42 ();
 FILLCELL_X8 FILLER_31_69 ();
 FILLCELL_X2 FILLER_31_113 ();
 FILLCELL_X2 FILLER_31_122 ();
 FILLCELL_X1 FILLER_31_124 ();
 FILLCELL_X4 FILLER_31_149 ();
 FILLCELL_X1 FILLER_31_157 ();
 FILLCELL_X32 FILLER_31_162 ();
 FILLCELL_X4 FILLER_31_194 ();
 FILLCELL_X2 FILLER_31_198 ();
 FILLCELL_X1 FILLER_31_204 ();
 FILLCELL_X8 FILLER_31_208 ();
 FILLCELL_X4 FILLER_31_216 ();
 FILLCELL_X1 FILLER_31_220 ();
 FILLCELL_X2 FILLER_31_226 ();
 FILLCELL_X16 FILLER_31_232 ();
 FILLCELL_X8 FILLER_31_248 ();
 FILLCELL_X4 FILLER_31_256 ();
 FILLCELL_X1 FILLER_31_260 ();
 FILLCELL_X4 FILLER_31_266 ();
 FILLCELL_X2 FILLER_31_270 ();
 FILLCELL_X8 FILLER_31_281 ();
 FILLCELL_X2 FILLER_31_289 ();
 FILLCELL_X1 FILLER_31_291 ();
 FILLCELL_X16 FILLER_31_311 ();
 FILLCELL_X4 FILLER_31_327 ();
 FILLCELL_X1 FILLER_31_331 ();
 FILLCELL_X2 FILLER_31_335 ();
 FILLCELL_X8 FILLER_31_340 ();
 FILLCELL_X2 FILLER_31_348 ();
 FILLCELL_X1 FILLER_31_350 ();
 FILLCELL_X16 FILLER_31_354 ();
 FILLCELL_X1 FILLER_31_370 ();
 FILLCELL_X4 FILLER_31_391 ();
 FILLCELL_X2 FILLER_31_404 ();
 FILLCELL_X4 FILLER_31_415 ();
 FILLCELL_X8 FILLER_32_1 ();
 FILLCELL_X4 FILLER_32_9 ();
 FILLCELL_X4 FILLER_32_19 ();
 FILLCELL_X1 FILLER_32_23 ();
 FILLCELL_X1 FILLER_32_33 ();
 FILLCELL_X2 FILLER_32_54 ();
 FILLCELL_X1 FILLER_32_56 ();
 FILLCELL_X8 FILLER_32_62 ();
 FILLCELL_X1 FILLER_32_70 ();
 FILLCELL_X2 FILLER_32_76 ();
 FILLCELL_X2 FILLER_32_91 ();
 FILLCELL_X1 FILLER_32_93 ();
 FILLCELL_X1 FILLER_32_101 ();
 FILLCELL_X2 FILLER_32_116 ();
 FILLCELL_X1 FILLER_32_118 ();
 FILLCELL_X8 FILLER_32_128 ();
 FILLCELL_X2 FILLER_32_136 ();
 FILLCELL_X4 FILLER_32_163 ();
 FILLCELL_X2 FILLER_32_167 ();
 FILLCELL_X16 FILLER_32_172 ();
 FILLCELL_X4 FILLER_32_188 ();
 FILLCELL_X2 FILLER_32_192 ();
 FILLCELL_X4 FILLER_32_213 ();
 FILLCELL_X2 FILLER_32_217 ();
 FILLCELL_X2 FILLER_32_247 ();
 FILLCELL_X1 FILLER_32_258 ();
 FILLCELL_X4 FILLER_32_265 ();
 FILLCELL_X8 FILLER_32_276 ();
 FILLCELL_X2 FILLER_32_306 ();
 FILLCELL_X2 FILLER_32_310 ();
 FILLCELL_X1 FILLER_32_316 ();
 FILLCELL_X2 FILLER_32_341 ();
 FILLCELL_X8 FILLER_32_352 ();
 FILLCELL_X1 FILLER_32_360 ();
 FILLCELL_X4 FILLER_32_365 ();
 FILLCELL_X2 FILLER_32_369 ();
 FILLCELL_X1 FILLER_32_371 ();
 FILLCELL_X2 FILLER_32_404 ();
 FILLCELL_X2 FILLER_32_409 ();
 FILLCELL_X1 FILLER_32_411 ();
 FILLCELL_X4 FILLER_32_415 ();
 FILLCELL_X4 FILLER_33_1 ();
 FILLCELL_X1 FILLER_33_5 ();
 FILLCELL_X2 FILLER_33_9 ();
 FILLCELL_X2 FILLER_33_21 ();
 FILLCELL_X1 FILLER_33_23 ();
 FILLCELL_X8 FILLER_33_34 ();
 FILLCELL_X2 FILLER_33_42 ();
 FILLCELL_X1 FILLER_33_44 ();
 FILLCELL_X2 FILLER_33_60 ();
 FILLCELL_X1 FILLER_33_87 ();
 FILLCELL_X4 FILLER_33_97 ();
 FILLCELL_X2 FILLER_33_120 ();
 FILLCELL_X2 FILLER_33_133 ();
 FILLCELL_X4 FILLER_33_149 ();
 FILLCELL_X2 FILLER_33_153 ();
 FILLCELL_X1 FILLER_33_155 ();
 FILLCELL_X4 FILLER_33_160 ();
 FILLCELL_X2 FILLER_33_164 ();
 FILLCELL_X4 FILLER_33_185 ();
 FILLCELL_X2 FILLER_33_189 ();
 FILLCELL_X1 FILLER_33_191 ();
 FILLCELL_X4 FILLER_33_202 ();
 FILLCELL_X2 FILLER_33_206 ();
 FILLCELL_X1 FILLER_33_208 ();
 FILLCELL_X2 FILLER_33_229 ();
 FILLCELL_X1 FILLER_33_231 ();
 FILLCELL_X2 FILLER_33_264 ();
 FILLCELL_X4 FILLER_33_285 ();
 FILLCELL_X2 FILLER_33_289 ();
 FILLCELL_X1 FILLER_33_291 ();
 FILLCELL_X2 FILLER_33_314 ();
 FILLCELL_X4 FILLER_33_325 ();
 FILLCELL_X1 FILLER_33_331 ();
 FILLCELL_X4 FILLER_33_340 ();
 FILLCELL_X2 FILLER_33_344 ();
 FILLCELL_X8 FILLER_33_363 ();
 FILLCELL_X4 FILLER_33_371 ();
 FILLCELL_X2 FILLER_33_375 ();
 FILLCELL_X8 FILLER_33_410 ();
 FILLCELL_X1 FILLER_33_418 ();
 FILLCELL_X2 FILLER_34_1 ();
 FILLCELL_X2 FILLER_34_43 ();
 FILLCELL_X4 FILLER_34_78 ();
 FILLCELL_X16 FILLER_34_107 ();
 FILLCELL_X8 FILLER_34_123 ();
 FILLCELL_X1 FILLER_34_131 ();
 FILLCELL_X4 FILLER_34_146 ();
 FILLCELL_X2 FILLER_34_159 ();
 FILLCELL_X16 FILLER_34_178 ();
 FILLCELL_X4 FILLER_34_194 ();
 FILLCELL_X1 FILLER_34_198 ();
 FILLCELL_X1 FILLER_34_224 ();
 FILLCELL_X8 FILLER_34_239 ();
 FILLCELL_X2 FILLER_34_247 ();
 FILLCELL_X8 FILLER_34_264 ();
 FILLCELL_X4 FILLER_34_272 ();
 FILLCELL_X4 FILLER_34_279 ();
 FILLCELL_X1 FILLER_34_283 ();
 FILLCELL_X2 FILLER_34_295 ();
 FILLCELL_X32 FILLER_34_339 ();
 FILLCELL_X2 FILLER_34_371 ();
 FILLCELL_X1 FILLER_34_373 ();
 FILLCELL_X1 FILLER_34_388 ();
 FILLCELL_X1 FILLER_34_415 ();
 FILLCELL_X2 FILLER_35_7 ();
 FILLCELL_X1 FILLER_35_9 ();
 FILLCELL_X2 FILLER_35_36 ();
 FILLCELL_X4 FILLER_35_41 ();
 FILLCELL_X1 FILLER_35_48 ();
 FILLCELL_X2 FILLER_35_53 ();
 FILLCELL_X1 FILLER_35_55 ();
 FILLCELL_X1 FILLER_35_62 ();
 FILLCELL_X2 FILLER_35_91 ();
 FILLCELL_X2 FILLER_35_132 ();
 FILLCELL_X1 FILLER_35_134 ();
 FILLCELL_X8 FILLER_35_142 ();
 FILLCELL_X1 FILLER_35_165 ();
 FILLCELL_X8 FILLER_35_177 ();
 FILLCELL_X4 FILLER_35_185 ();
 FILLCELL_X1 FILLER_35_189 ();
 FILLCELL_X8 FILLER_35_218 ();
 FILLCELL_X2 FILLER_35_226 ();
 FILLCELL_X2 FILLER_35_236 ();
 FILLCELL_X2 FILLER_35_248 ();
 FILLCELL_X1 FILLER_35_250 ();
 FILLCELL_X8 FILLER_35_260 ();
 FILLCELL_X4 FILLER_35_268 ();
 FILLCELL_X1 FILLER_35_272 ();
 FILLCELL_X16 FILLER_35_342 ();
 FILLCELL_X8 FILLER_35_358 ();
 FILLCELL_X4 FILLER_35_366 ();
 FILLCELL_X2 FILLER_35_370 ();
 FILLCELL_X2 FILLER_35_404 ();
 FILLCELL_X1 FILLER_35_406 ();
 FILLCELL_X2 FILLER_35_416 ();
 FILLCELL_X1 FILLER_35_418 ();
 FILLCELL_X8 FILLER_36_4 ();
 FILLCELL_X2 FILLER_36_12 ();
 FILLCELL_X2 FILLER_36_62 ();
 FILLCELL_X2 FILLER_36_85 ();
 FILLCELL_X1 FILLER_36_92 ();
 FILLCELL_X2 FILLER_36_113 ();
 FILLCELL_X2 FILLER_36_128 ();
 FILLCELL_X1 FILLER_36_135 ();
 FILLCELL_X8 FILLER_36_143 ();
 FILLCELL_X2 FILLER_36_164 ();
 FILLCELL_X4 FILLER_36_185 ();
 FILLCELL_X2 FILLER_36_189 ();
 FILLCELL_X8 FILLER_36_195 ();
 FILLCELL_X1 FILLER_36_213 ();
 FILLCELL_X16 FILLER_36_234 ();
 FILLCELL_X4 FILLER_36_250 ();
 FILLCELL_X8 FILLER_36_273 ();
 FILLCELL_X2 FILLER_36_281 ();
 FILLCELL_X1 FILLER_36_283 ();
 FILLCELL_X1 FILLER_36_298 ();
 FILLCELL_X8 FILLER_36_311 ();
 FILLCELL_X4 FILLER_36_319 ();
 FILLCELL_X2 FILLER_36_323 ();
 FILLCELL_X1 FILLER_36_325 ();
 FILLCELL_X4 FILLER_36_345 ();
 FILLCELL_X1 FILLER_36_349 ();
 FILLCELL_X4 FILLER_36_361 ();
 FILLCELL_X1 FILLER_36_365 ();
 FILLCELL_X2 FILLER_36_414 ();
 FILLCELL_X2 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_8 ();
 FILLCELL_X8 FILLER_37_40 ();
 FILLCELL_X2 FILLER_37_48 ();
 FILLCELL_X2 FILLER_37_54 ();
 FILLCELL_X1 FILLER_37_67 ();
 FILLCELL_X4 FILLER_37_98 ();
 FILLCELL_X16 FILLER_37_114 ();
 FILLCELL_X4 FILLER_37_130 ();
 FILLCELL_X2 FILLER_37_134 ();
 FILLCELL_X4 FILLER_37_153 ();
 FILLCELL_X1 FILLER_37_157 ();
 FILLCELL_X4 FILLER_37_162 ();
 FILLCELL_X16 FILLER_37_181 ();
 FILLCELL_X4 FILLER_37_197 ();
 FILLCELL_X2 FILLER_37_201 ();
 FILLCELL_X16 FILLER_37_207 ();
 FILLCELL_X8 FILLER_37_223 ();
 FILLCELL_X1 FILLER_37_231 ();
 FILLCELL_X4 FILLER_37_236 ();
 FILLCELL_X8 FILLER_37_246 ();
 FILLCELL_X1 FILLER_37_254 ();
 FILLCELL_X16 FILLER_37_261 ();
 FILLCELL_X2 FILLER_37_280 ();
 FILLCELL_X4 FILLER_37_307 ();
 FILLCELL_X2 FILLER_37_311 ();
 FILLCELL_X1 FILLER_37_313 ();
 FILLCELL_X16 FILLER_37_323 ();
 FILLCELL_X1 FILLER_37_339 ();
 FILLCELL_X1 FILLER_37_357 ();
 FILLCELL_X4 FILLER_37_379 ();
 FILLCELL_X2 FILLER_37_386 ();
 FILLCELL_X1 FILLER_37_388 ();
 FILLCELL_X1 FILLER_37_398 ();
 FILLCELL_X4 FILLER_37_403 ();
 FILLCELL_X2 FILLER_37_407 ();
 FILLCELL_X1 FILLER_37_412 ();
 FILLCELL_X4 FILLER_38_36 ();
 FILLCELL_X2 FILLER_38_40 ();
 FILLCELL_X1 FILLER_38_42 ();
 FILLCELL_X32 FILLER_38_47 ();
 FILLCELL_X4 FILLER_38_79 ();
 FILLCELL_X16 FILLER_38_98 ();
 FILLCELL_X4 FILLER_38_114 ();
 FILLCELL_X2 FILLER_38_118 ();
 FILLCELL_X4 FILLER_38_124 ();
 FILLCELL_X1 FILLER_38_131 ();
 FILLCELL_X1 FILLER_38_135 ();
 FILLCELL_X8 FILLER_38_139 ();
 FILLCELL_X2 FILLER_38_147 ();
 FILLCELL_X1 FILLER_38_158 ();
 FILLCELL_X2 FILLER_38_170 ();
 FILLCELL_X1 FILLER_38_177 ();
 FILLCELL_X2 FILLER_38_197 ();
 FILLCELL_X4 FILLER_38_218 ();
 FILLCELL_X2 FILLER_38_222 ();
 FILLCELL_X2 FILLER_38_248 ();
 FILLCELL_X4 FILLER_38_265 ();
 FILLCELL_X1 FILLER_38_269 ();
 FILLCELL_X2 FILLER_38_289 ();
 FILLCELL_X1 FILLER_38_291 ();
 FILLCELL_X2 FILLER_38_311 ();
 FILLCELL_X4 FILLER_38_342 ();
 FILLCELL_X2 FILLER_38_346 ();
 FILLCELL_X1 FILLER_38_348 ();
 FILLCELL_X1 FILLER_38_356 ();
 FILLCELL_X2 FILLER_38_368 ();
 FILLCELL_X1 FILLER_38_370 ();
 FILLCELL_X2 FILLER_38_382 ();
 FILLCELL_X4 FILLER_38_392 ();
 FILLCELL_X1 FILLER_38_401 ();
 FILLCELL_X2 FILLER_39_10 ();
 FILLCELL_X1 FILLER_39_15 ();
 FILLCELL_X1 FILLER_39_22 ();
 FILLCELL_X4 FILLER_39_46 ();
 FILLCELL_X1 FILLER_39_50 ();
 FILLCELL_X4 FILLER_39_57 ();
 FILLCELL_X2 FILLER_39_61 ();
 FILLCELL_X2 FILLER_39_73 ();
 FILLCELL_X2 FILLER_39_79 ();
 FILLCELL_X1 FILLER_39_81 ();
 FILLCELL_X2 FILLER_39_101 ();
 FILLCELL_X1 FILLER_39_103 ();
 FILLCELL_X1 FILLER_39_134 ();
 FILLCELL_X1 FILLER_39_140 ();
 FILLCELL_X4 FILLER_39_145 ();
 FILLCELL_X1 FILLER_39_153 ();
 FILLCELL_X4 FILLER_39_169 ();
 FILLCELL_X2 FILLER_39_173 ();
 FILLCELL_X8 FILLER_39_185 ();
 FILLCELL_X4 FILLER_39_193 ();
 FILLCELL_X1 FILLER_39_197 ();
 FILLCELL_X1 FILLER_39_208 ();
 FILLCELL_X1 FILLER_39_216 ();
 FILLCELL_X8 FILLER_39_222 ();
 FILLCELL_X1 FILLER_39_230 ();
 FILLCELL_X1 FILLER_39_234 ();
 FILLCELL_X4 FILLER_39_246 ();
 FILLCELL_X1 FILLER_39_250 ();
 FILLCELL_X8 FILLER_39_254 ();
 FILLCELL_X2 FILLER_39_280 ();
 FILLCELL_X2 FILLER_39_301 ();
 FILLCELL_X1 FILLER_39_313 ();
 FILLCELL_X4 FILLER_39_318 ();
 FILLCELL_X1 FILLER_39_322 ();
 FILLCELL_X1 FILLER_39_330 ();
 FILLCELL_X4 FILLER_39_338 ();
 FILLCELL_X1 FILLER_39_342 ();
 FILLCELL_X8 FILLER_39_350 ();
 FILLCELL_X2 FILLER_39_358 ();
 FILLCELL_X1 FILLER_39_360 ();
 FILLCELL_X2 FILLER_39_368 ();
 FILLCELL_X1 FILLER_39_370 ();
 FILLCELL_X1 FILLER_39_398 ();
 FILLCELL_X1 FILLER_39_415 ();
 FILLCELL_X1 FILLER_40_32 ();
 FILLCELL_X2 FILLER_40_35 ();
 FILLCELL_X1 FILLER_40_37 ();
 FILLCELL_X2 FILLER_40_91 ();
 FILLCELL_X1 FILLER_40_93 ();
 FILLCELL_X16 FILLER_40_98 ();
 FILLCELL_X1 FILLER_40_114 ();
 FILLCELL_X4 FILLER_40_122 ();
 FILLCELL_X2 FILLER_40_126 ();
 FILLCELL_X1 FILLER_40_132 ();
 FILLCELL_X1 FILLER_40_143 ();
 FILLCELL_X2 FILLER_40_164 ();
 FILLCELL_X8 FILLER_40_185 ();
 FILLCELL_X4 FILLER_40_193 ();
 FILLCELL_X2 FILLER_40_197 ();
 FILLCELL_X1 FILLER_40_199 ();
 FILLCELL_X2 FILLER_40_210 ();
 FILLCELL_X1 FILLER_40_212 ();
 FILLCELL_X2 FILLER_40_223 ();
 FILLCELL_X1 FILLER_40_225 ();
 FILLCELL_X16 FILLER_40_232 ();
 FILLCELL_X4 FILLER_40_248 ();
 FILLCELL_X1 FILLER_40_252 ();
 FILLCELL_X4 FILLER_40_260 ();
 FILLCELL_X2 FILLER_40_264 ();
 FILLCELL_X1 FILLER_40_266 ();
 FILLCELL_X8 FILLER_40_270 ();
 FILLCELL_X2 FILLER_40_278 ();
 FILLCELL_X2 FILLER_40_288 ();
 FILLCELL_X1 FILLER_40_290 ();
 FILLCELL_X1 FILLER_40_317 ();
 FILLCELL_X1 FILLER_40_339 ();
 FILLCELL_X1 FILLER_40_347 ();
 FILLCELL_X2 FILLER_40_366 ();
 FILLCELL_X1 FILLER_40_368 ();
 FILLCELL_X2 FILLER_40_373 ();
 FILLCELL_X1 FILLER_40_375 ();
 FILLCELL_X1 FILLER_40_392 ();
 FILLCELL_X8 FILLER_40_404 ();
 FILLCELL_X4 FILLER_40_412 ();
 FILLCELL_X2 FILLER_40_416 ();
 FILLCELL_X1 FILLER_40_418 ();
 FILLCELL_X2 FILLER_41_1 ();
 FILLCELL_X1 FILLER_41_3 ();
 FILLCELL_X4 FILLER_41_7 ();
 FILLCELL_X1 FILLER_41_11 ();
 FILLCELL_X2 FILLER_41_15 ();
 FILLCELL_X1 FILLER_41_17 ();
 FILLCELL_X2 FILLER_41_21 ();
 FILLCELL_X2 FILLER_41_26 ();
 FILLCELL_X1 FILLER_41_28 ();
 FILLCELL_X8 FILLER_41_45 ();
 FILLCELL_X4 FILLER_41_53 ();
 FILLCELL_X2 FILLER_41_57 ();
 FILLCELL_X1 FILLER_41_74 ();
 FILLCELL_X1 FILLER_41_78 ();
 FILLCELL_X2 FILLER_41_88 ();
 FILLCELL_X1 FILLER_41_90 ();
 FILLCELL_X8 FILLER_41_113 ();
 FILLCELL_X4 FILLER_41_121 ();
 FILLCELL_X2 FILLER_41_125 ();
 FILLCELL_X4 FILLER_41_153 ();
 FILLCELL_X8 FILLER_41_161 ();
 FILLCELL_X4 FILLER_41_169 ();
 FILLCELL_X1 FILLER_41_173 ();
 FILLCELL_X8 FILLER_41_184 ();
 FILLCELL_X2 FILLER_41_192 ();
 FILLCELL_X1 FILLER_41_197 ();
 FILLCELL_X8 FILLER_41_202 ();
 FILLCELL_X2 FILLER_41_210 ();
 FILLCELL_X1 FILLER_41_226 ();
 FILLCELL_X2 FILLER_41_229 ();
 FILLCELL_X2 FILLER_41_234 ();
 FILLCELL_X1 FILLER_41_236 ();
 FILLCELL_X8 FILLER_41_241 ();
 FILLCELL_X1 FILLER_41_276 ();
 FILLCELL_X4 FILLER_41_285 ();
 FILLCELL_X2 FILLER_41_293 ();
 FILLCELL_X1 FILLER_41_349 ();
 FILLCELL_X2 FILLER_41_358 ();
 FILLCELL_X2 FILLER_41_371 ();
 FILLCELL_X2 FILLER_41_381 ();
 FILLCELL_X1 FILLER_41_383 ();
 FILLCELL_X8 FILLER_42_1 ();
 FILLCELL_X4 FILLER_42_9 ();
 FILLCELL_X16 FILLER_42_32 ();
 FILLCELL_X4 FILLER_42_48 ();
 FILLCELL_X2 FILLER_42_52 ();
 FILLCELL_X16 FILLER_42_83 ();
 FILLCELL_X4 FILLER_42_99 ();
 FILLCELL_X1 FILLER_42_103 ();
 FILLCELL_X8 FILLER_42_121 ();
 FILLCELL_X2 FILLER_42_143 ();
 FILLCELL_X1 FILLER_42_145 ();
 FILLCELL_X1 FILLER_42_150 ();
 FILLCELL_X1 FILLER_42_158 ();
 FILLCELL_X16 FILLER_42_180 ();
 FILLCELL_X4 FILLER_42_196 ();
 FILLCELL_X1 FILLER_42_207 ();
 FILLCELL_X8 FILLER_42_211 ();
 FILLCELL_X1 FILLER_42_219 ();
 FILLCELL_X1 FILLER_42_224 ();
 FILLCELL_X2 FILLER_42_234 ();
 FILLCELL_X16 FILLER_42_240 ();
 FILLCELL_X4 FILLER_42_256 ();
 FILLCELL_X8 FILLER_42_262 ();
 FILLCELL_X2 FILLER_42_270 ();
 FILLCELL_X1 FILLER_42_272 ();
 FILLCELL_X2 FILLER_42_285 ();
 FILLCELL_X8 FILLER_42_325 ();
 FILLCELL_X4 FILLER_42_333 ();
 FILLCELL_X2 FILLER_42_337 ();
 FILLCELL_X1 FILLER_42_339 ();
 FILLCELL_X4 FILLER_42_347 ();
 FILLCELL_X1 FILLER_42_351 ();
 FILLCELL_X8 FILLER_42_359 ();
 FILLCELL_X4 FILLER_42_367 ();
 FILLCELL_X2 FILLER_42_417 ();
 FILLCELL_X2 FILLER_43_1 ();
 FILLCELL_X2 FILLER_43_23 ();
 FILLCELL_X1 FILLER_43_25 ();
 FILLCELL_X4 FILLER_43_29 ();
 FILLCELL_X8 FILLER_43_50 ();
 FILLCELL_X2 FILLER_43_58 ();
 FILLCELL_X4 FILLER_43_100 ();
 FILLCELL_X1 FILLER_43_104 ();
 FILLCELL_X16 FILLER_43_115 ();
 FILLCELL_X1 FILLER_43_131 ();
 FILLCELL_X1 FILLER_43_149 ();
 FILLCELL_X4 FILLER_43_167 ();
 FILLCELL_X2 FILLER_43_190 ();
 FILLCELL_X2 FILLER_43_209 ();
 FILLCELL_X2 FILLER_43_228 ();
 FILLCELL_X1 FILLER_43_230 ();
 FILLCELL_X8 FILLER_43_282 ();
 FILLCELL_X4 FILLER_43_290 ();
 FILLCELL_X2 FILLER_43_305 ();
 FILLCELL_X1 FILLER_43_307 ();
 FILLCELL_X8 FILLER_43_312 ();
 FILLCELL_X4 FILLER_43_320 ();
 FILLCELL_X8 FILLER_43_327 ();
 FILLCELL_X2 FILLER_43_376 ();
 FILLCELL_X8 FILLER_43_400 ();
 FILLCELL_X1 FILLER_43_408 ();
 FILLCELL_X1 FILLER_43_412 ();
 FILLCELL_X8 FILLER_44_1 ();
 FILLCELL_X8 FILLER_44_12 ();
 FILLCELL_X2 FILLER_44_20 ();
 FILLCELL_X1 FILLER_44_22 ();
 FILLCELL_X16 FILLER_44_62 ();
 FILLCELL_X8 FILLER_44_78 ();
 FILLCELL_X4 FILLER_44_86 ();
 FILLCELL_X2 FILLER_44_90 ();
 FILLCELL_X1 FILLER_44_92 ();
 FILLCELL_X4 FILLER_44_117 ();
 FILLCELL_X2 FILLER_44_121 ();
 FILLCELL_X1 FILLER_44_123 ();
 FILLCELL_X8 FILLER_44_143 ();
 FILLCELL_X1 FILLER_44_151 ();
 FILLCELL_X16 FILLER_44_180 ();
 FILLCELL_X8 FILLER_44_196 ();
 FILLCELL_X4 FILLER_44_204 ();
 FILLCELL_X2 FILLER_44_208 ();
 FILLCELL_X4 FILLER_44_212 ();
 FILLCELL_X1 FILLER_44_216 ();
 FILLCELL_X4 FILLER_44_219 ();
 FILLCELL_X2 FILLER_44_223 ();
 FILLCELL_X1 FILLER_44_225 ();
 FILLCELL_X4 FILLER_44_233 ();
 FILLCELL_X1 FILLER_44_237 ();
 FILLCELL_X8 FILLER_44_257 ();
 FILLCELL_X16 FILLER_44_284 ();
 FILLCELL_X2 FILLER_44_300 ();
 FILLCELL_X1 FILLER_44_302 ();
 FILLCELL_X8 FILLER_44_310 ();
 FILLCELL_X2 FILLER_44_318 ();
 FILLCELL_X8 FILLER_44_348 ();
 FILLCELL_X2 FILLER_44_356 ();
 FILLCELL_X1 FILLER_44_361 ();
 FILLCELL_X4 FILLER_44_384 ();
 FILLCELL_X2 FILLER_44_401 ();
 FILLCELL_X1 FILLER_44_403 ();
 FILLCELL_X4 FILLER_44_407 ();
 FILLCELL_X2 FILLER_44_411 ();
 FILLCELL_X8 FILLER_45_1 ();
 FILLCELL_X4 FILLER_45_9 ();
 FILLCELL_X2 FILLER_45_13 ();
 FILLCELL_X1 FILLER_45_15 ();
 FILLCELL_X8 FILLER_45_19 ();
 FILLCELL_X1 FILLER_45_46 ();
 FILLCELL_X8 FILLER_45_50 ();
 FILLCELL_X2 FILLER_45_72 ();
 FILLCELL_X2 FILLER_45_81 ();
 FILLCELL_X4 FILLER_45_94 ();
 FILLCELL_X2 FILLER_45_98 ();
 FILLCELL_X1 FILLER_45_100 ();
 FILLCELL_X8 FILLER_45_110 ();
 FILLCELL_X4 FILLER_45_118 ();
 FILLCELL_X2 FILLER_45_122 ();
 FILLCELL_X1 FILLER_45_137 ();
 FILLCELL_X16 FILLER_45_140 ();
 FILLCELL_X4 FILLER_45_156 ();
 FILLCELL_X4 FILLER_45_169 ();
 FILLCELL_X16 FILLER_45_177 ();
 FILLCELL_X4 FILLER_45_193 ();
 FILLCELL_X1 FILLER_45_197 ();
 FILLCELL_X8 FILLER_45_220 ();
 FILLCELL_X16 FILLER_45_250 ();
 FILLCELL_X4 FILLER_45_266 ();
 FILLCELL_X1 FILLER_45_270 ();
 FILLCELL_X8 FILLER_45_283 ();
 FILLCELL_X4 FILLER_45_291 ();
 FILLCELL_X2 FILLER_45_295 ();
 FILLCELL_X1 FILLER_45_297 ();
 FILLCELL_X1 FILLER_45_304 ();
 FILLCELL_X4 FILLER_45_315 ();
 FILLCELL_X1 FILLER_45_319 ();
 FILLCELL_X4 FILLER_45_336 ();
 FILLCELL_X1 FILLER_45_340 ();
 FILLCELL_X4 FILLER_45_349 ();
 FILLCELL_X1 FILLER_45_353 ();
 FILLCELL_X8 FILLER_45_360 ();
 FILLCELL_X2 FILLER_45_370 ();
 FILLCELL_X4 FILLER_45_381 ();
 FILLCELL_X2 FILLER_45_385 ();
 FILLCELL_X1 FILLER_45_387 ();
 FILLCELL_X4 FILLER_45_391 ();
 FILLCELL_X1 FILLER_45_395 ();
 FILLCELL_X8 FILLER_45_406 ();
 FILLCELL_X2 FILLER_45_414 ();
 FILLCELL_X8 FILLER_46_1 ();
 FILLCELL_X4 FILLER_46_9 ();
 FILLCELL_X2 FILLER_46_13 ();
 FILLCELL_X1 FILLER_46_15 ();
 FILLCELL_X8 FILLER_46_19 ();
 FILLCELL_X1 FILLER_46_30 ();
 FILLCELL_X2 FILLER_46_56 ();
 FILLCELL_X8 FILLER_46_75 ();
 FILLCELL_X2 FILLER_46_83 ();
 FILLCELL_X4 FILLER_46_91 ();
 FILLCELL_X2 FILLER_46_95 ();
 FILLCELL_X8 FILLER_46_101 ();
 FILLCELL_X4 FILLER_46_109 ();
 FILLCELL_X2 FILLER_46_113 ();
 FILLCELL_X8 FILLER_46_135 ();
 FILLCELL_X4 FILLER_46_143 ();
 FILLCELL_X1 FILLER_46_147 ();
 FILLCELL_X4 FILLER_46_154 ();
 FILLCELL_X2 FILLER_46_158 ();
 FILLCELL_X1 FILLER_46_160 ();
 FILLCELL_X8 FILLER_46_185 ();
 FILLCELL_X2 FILLER_46_193 ();
 FILLCELL_X1 FILLER_46_195 ();
 FILLCELL_X2 FILLER_46_218 ();
 FILLCELL_X2 FILLER_46_224 ();
 FILLCELL_X1 FILLER_46_240 ();
 FILLCELL_X4 FILLER_46_249 ();
 FILLCELL_X4 FILLER_46_279 ();
 FILLCELL_X8 FILLER_46_287 ();
 FILLCELL_X4 FILLER_46_295 ();
 FILLCELL_X1 FILLER_46_299 ();
 FILLCELL_X8 FILLER_46_319 ();
 FILLCELL_X1 FILLER_46_327 ();
 FILLCELL_X2 FILLER_46_333 ();
 FILLCELL_X1 FILLER_46_340 ();
 FILLCELL_X1 FILLER_46_356 ();
 FILLCELL_X4 FILLER_46_362 ();
 FILLCELL_X2 FILLER_46_366 ();
 FILLCELL_X4 FILLER_46_388 ();
 FILLCELL_X1 FILLER_46_392 ();
 FILLCELL_X8 FILLER_47_1 ();
 FILLCELL_X2 FILLER_47_9 ();
 FILLCELL_X8 FILLER_47_14 ();
 FILLCELL_X1 FILLER_47_22 ();
 FILLCELL_X32 FILLER_47_43 ();
 FILLCELL_X8 FILLER_47_75 ();
 FILLCELL_X1 FILLER_47_92 ();
 FILLCELL_X16 FILLER_47_99 ();
 FILLCELL_X2 FILLER_47_126 ();
 FILLCELL_X16 FILLER_47_131 ();
 FILLCELL_X2 FILLER_47_147 ();
 FILLCELL_X2 FILLER_47_152 ();
 FILLCELL_X1 FILLER_47_154 ();
 FILLCELL_X4 FILLER_47_157 ();
 FILLCELL_X1 FILLER_47_165 ();
 FILLCELL_X2 FILLER_47_168 ();
 FILLCELL_X4 FILLER_47_172 ();
 FILLCELL_X2 FILLER_47_176 ();
 FILLCELL_X1 FILLER_47_178 ();
 FILLCELL_X1 FILLER_47_184 ();
 FILLCELL_X16 FILLER_47_188 ();
 FILLCELL_X8 FILLER_47_204 ();
 FILLCELL_X4 FILLER_47_212 ();
 FILLCELL_X2 FILLER_47_216 ();
 FILLCELL_X1 FILLER_47_218 ();
 FILLCELL_X4 FILLER_47_223 ();
 FILLCELL_X1 FILLER_47_227 ();
 FILLCELL_X1 FILLER_47_237 ();
 FILLCELL_X16 FILLER_47_250 ();
 FILLCELL_X2 FILLER_47_266 ();
 FILLCELL_X8 FILLER_47_276 ();
 FILLCELL_X2 FILLER_47_284 ();
 FILLCELL_X8 FILLER_47_291 ();
 FILLCELL_X4 FILLER_47_299 ();
 FILLCELL_X2 FILLER_47_303 ();
 FILLCELL_X8 FILLER_47_309 ();
 FILLCELL_X1 FILLER_47_317 ();
 FILLCELL_X16 FILLER_47_321 ();
 FILLCELL_X2 FILLER_47_337 ();
 FILLCELL_X1 FILLER_47_339 ();
 FILLCELL_X1 FILLER_47_351 ();
 FILLCELL_X4 FILLER_47_356 ();
 FILLCELL_X1 FILLER_47_360 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X2 FILLER_48_65 ();
 FILLCELL_X4 FILLER_48_101 ();
 FILLCELL_X1 FILLER_48_105 ();
 FILLCELL_X1 FILLER_48_112 ();
 FILLCELL_X1 FILLER_48_120 ();
 FILLCELL_X2 FILLER_48_128 ();
 FILLCELL_X8 FILLER_48_135 ();
 FILLCELL_X1 FILLER_48_143 ();
 FILLCELL_X2 FILLER_48_179 ();
 FILLCELL_X1 FILLER_48_188 ();
 FILLCELL_X8 FILLER_48_194 ();
 FILLCELL_X2 FILLER_48_202 ();
 FILLCELL_X2 FILLER_48_223 ();
 FILLCELL_X1 FILLER_48_225 ();
 FILLCELL_X8 FILLER_48_247 ();
 FILLCELL_X1 FILLER_48_255 ();
 FILLCELL_X2 FILLER_48_265 ();
 FILLCELL_X1 FILLER_48_267 ();
 FILLCELL_X1 FILLER_48_277 ();
 FILLCELL_X8 FILLER_48_283 ();
 FILLCELL_X8 FILLER_48_305 ();
 FILLCELL_X2 FILLER_48_313 ();
 FILLCELL_X8 FILLER_48_324 ();
 FILLCELL_X4 FILLER_48_332 ();
 FILLCELL_X2 FILLER_48_336 ();
 FILLCELL_X1 FILLER_48_338 ();
 FILLCELL_X8 FILLER_48_348 ();
 FILLCELL_X4 FILLER_48_356 ();
 FILLCELL_X2 FILLER_48_360 ();
 FILLCELL_X8 FILLER_48_376 ();
 FILLCELL_X4 FILLER_48_384 ();
 FILLCELL_X1 FILLER_48_388 ();
 FILLCELL_X1 FILLER_48_418 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X16 FILLER_49_33 ();
 FILLCELL_X2 FILLER_49_49 ();
 FILLCELL_X1 FILLER_49_51 ();
 FILLCELL_X4 FILLER_49_69 ();
 FILLCELL_X2 FILLER_49_90 ();
 FILLCELL_X8 FILLER_49_97 ();
 FILLCELL_X2 FILLER_49_105 ();
 FILLCELL_X2 FILLER_49_111 ();
 FILLCELL_X1 FILLER_49_113 ();
 FILLCELL_X1 FILLER_49_123 ();
 FILLCELL_X16 FILLER_49_128 ();
 FILLCELL_X8 FILLER_49_144 ();
 FILLCELL_X4 FILLER_49_152 ();
 FILLCELL_X1 FILLER_49_156 ();
 FILLCELL_X4 FILLER_49_165 ();
 FILLCELL_X2 FILLER_49_177 ();
 FILLCELL_X16 FILLER_49_202 ();
 FILLCELL_X8 FILLER_49_218 ();
 FILLCELL_X1 FILLER_49_226 ();
 FILLCELL_X2 FILLER_49_246 ();
 FILLCELL_X8 FILLER_49_280 ();
 FILLCELL_X2 FILLER_49_288 ();
 FILLCELL_X1 FILLER_49_290 ();
 FILLCELL_X1 FILLER_49_310 ();
 FILLCELL_X8 FILLER_49_330 ();
 FILLCELL_X2 FILLER_49_338 ();
 FILLCELL_X1 FILLER_49_340 ();
 FILLCELL_X16 FILLER_49_360 ();
 FILLCELL_X4 FILLER_49_397 ();
 FILLCELL_X2 FILLER_49_401 ();
 FILLCELL_X1 FILLER_49_403 ();
 FILLCELL_X2 FILLER_49_416 ();
 FILLCELL_X1 FILLER_49_418 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X4 FILLER_50_65 ();
 FILLCELL_X2 FILLER_50_88 ();
 FILLCELL_X1 FILLER_50_90 ();
 FILLCELL_X8 FILLER_50_97 ();
 FILLCELL_X1 FILLER_50_105 ();
 FILLCELL_X1 FILLER_50_126 ();
 FILLCELL_X4 FILLER_50_132 ();
 FILLCELL_X2 FILLER_50_136 ();
 FILLCELL_X1 FILLER_50_138 ();
 FILLCELL_X1 FILLER_50_147 ();
 FILLCELL_X8 FILLER_50_153 ();
 FILLCELL_X32 FILLER_50_176 ();
 FILLCELL_X32 FILLER_50_208 ();
 FILLCELL_X16 FILLER_50_240 ();
 FILLCELL_X8 FILLER_50_256 ();
 FILLCELL_X2 FILLER_50_264 ();
 FILLCELL_X1 FILLER_50_266 ();
 FILLCELL_X2 FILLER_50_273 ();
 FILLCELL_X4 FILLER_50_294 ();
 FILLCELL_X1 FILLER_50_298 ();
 FILLCELL_X8 FILLER_50_304 ();
 FILLCELL_X4 FILLER_50_312 ();
 FILLCELL_X2 FILLER_50_316 ();
 FILLCELL_X2 FILLER_50_323 ();
 FILLCELL_X4 FILLER_50_329 ();
 FILLCELL_X1 FILLER_50_341 ();
 FILLCELL_X1 FILLER_50_348 ();
 FILLCELL_X1 FILLER_50_353 ();
 FILLCELL_X4 FILLER_50_359 ();
 FILLCELL_X1 FILLER_50_376 ();
 FILLCELL_X1 FILLER_50_386 ();
 FILLCELL_X8 FILLER_50_404 ();
 FILLCELL_X4 FILLER_50_412 ();
 FILLCELL_X2 FILLER_50_416 ();
 FILLCELL_X1 FILLER_50_418 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X16 FILLER_51_65 ();
 FILLCELL_X8 FILLER_51_81 ();
 FILLCELL_X2 FILLER_51_89 ();
 FILLCELL_X4 FILLER_51_102 ();
 FILLCELL_X8 FILLER_51_109 ();
 FILLCELL_X2 FILLER_51_117 ();
 FILLCELL_X2 FILLER_51_128 ();
 FILLCELL_X8 FILLER_51_136 ();
 FILLCELL_X4 FILLER_51_144 ();
 FILLCELL_X2 FILLER_51_154 ();
 FILLCELL_X1 FILLER_51_162 ();
 FILLCELL_X4 FILLER_51_165 ();
 FILLCELL_X1 FILLER_51_169 ();
 FILLCELL_X4 FILLER_51_176 ();
 FILLCELL_X1 FILLER_51_180 ();
 FILLCELL_X32 FILLER_51_184 ();
 FILLCELL_X32 FILLER_51_216 ();
 FILLCELL_X8 FILLER_51_248 ();
 FILLCELL_X4 FILLER_51_256 ();
 FILLCELL_X4 FILLER_51_263 ();
 FILLCELL_X2 FILLER_51_267 ();
 FILLCELL_X4 FILLER_51_272 ();
 FILLCELL_X2 FILLER_51_276 ();
 FILLCELL_X2 FILLER_51_285 ();
 FILLCELL_X2 FILLER_51_290 ();
 FILLCELL_X1 FILLER_51_292 ();
 FILLCELL_X4 FILLER_51_297 ();
 FILLCELL_X2 FILLER_51_315 ();
 FILLCELL_X1 FILLER_51_317 ();
 FILLCELL_X2 FILLER_51_332 ();
 FILLCELL_X1 FILLER_51_351 ();
 FILLCELL_X1 FILLER_51_357 ();
 FILLCELL_X2 FILLER_51_371 ();
 FILLCELL_X2 FILLER_51_383 ();
 FILLCELL_X2 FILLER_51_391 ();
 FILLCELL_X4 FILLER_51_412 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X8 FILLER_52_65 ();
 FILLCELL_X4 FILLER_52_73 ();
 FILLCELL_X8 FILLER_52_96 ();
 FILLCELL_X2 FILLER_52_104 ();
 FILLCELL_X1 FILLER_52_106 ();
 FILLCELL_X4 FILLER_52_117 ();
 FILLCELL_X1 FILLER_52_121 ();
 FILLCELL_X4 FILLER_52_128 ();
 FILLCELL_X2 FILLER_52_132 ();
 FILLCELL_X8 FILLER_52_137 ();
 FILLCELL_X4 FILLER_52_145 ();
 FILLCELL_X4 FILLER_52_152 ();
 FILLCELL_X4 FILLER_52_159 ();
 FILLCELL_X2 FILLER_52_163 ();
 FILLCELL_X1 FILLER_52_165 ();
 FILLCELL_X2 FILLER_52_172 ();
 FILLCELL_X32 FILLER_52_177 ();
 FILLCELL_X32 FILLER_52_209 ();
 FILLCELL_X8 FILLER_52_241 ();
 FILLCELL_X2 FILLER_52_249 ();
 FILLCELL_X4 FILLER_52_268 ();
 FILLCELL_X1 FILLER_52_272 ();
 FILLCELL_X1 FILLER_52_293 ();
 FILLCELL_X1 FILLER_52_300 ();
 FILLCELL_X1 FILLER_52_307 ();
 FILLCELL_X8 FILLER_52_312 ();
 FILLCELL_X1 FILLER_52_320 ();
 FILLCELL_X4 FILLER_52_333 ();
 FILLCELL_X2 FILLER_52_348 ();
 FILLCELL_X1 FILLER_52_350 ();
 FILLCELL_X4 FILLER_52_360 ();
 FILLCELL_X2 FILLER_52_364 ();
 FILLCELL_X1 FILLER_52_370 ();
 FILLCELL_X8 FILLER_52_384 ();
 FILLCELL_X1 FILLER_52_399 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X16 FILLER_53_65 ();
 FILLCELL_X8 FILLER_53_81 ();
 FILLCELL_X2 FILLER_53_89 ();
 FILLCELL_X1 FILLER_53_91 ();
 FILLCELL_X8 FILLER_53_112 ();
 FILLCELL_X4 FILLER_53_120 ();
 FILLCELL_X2 FILLER_53_124 ();
 FILLCELL_X1 FILLER_53_126 ();
 FILLCELL_X2 FILLER_53_130 ();
 FILLCELL_X1 FILLER_53_132 ();
 FILLCELL_X2 FILLER_53_150 ();
 FILLCELL_X1 FILLER_53_152 ();
 FILLCELL_X1 FILLER_53_173 ();
 FILLCELL_X32 FILLER_53_198 ();
 FILLCELL_X32 FILLER_53_230 ();
 FILLCELL_X4 FILLER_53_262 ();
 FILLCELL_X1 FILLER_53_266 ();
 FILLCELL_X8 FILLER_53_284 ();
 FILLCELL_X1 FILLER_53_292 ();
 FILLCELL_X4 FILLER_53_310 ();
 FILLCELL_X1 FILLER_53_314 ();
 FILLCELL_X8 FILLER_53_337 ();
 FILLCELL_X2 FILLER_53_345 ();
 FILLCELL_X8 FILLER_53_375 ();
 FILLCELL_X4 FILLER_53_392 ();
 FILLCELL_X1 FILLER_53_396 ();
 FILLCELL_X16 FILLER_53_400 ();
 FILLCELL_X2 FILLER_53_416 ();
 FILLCELL_X1 FILLER_53_418 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X2 FILLER_54_97 ();
 FILLCELL_X1 FILLER_54_123 ();
 FILLCELL_X1 FILLER_54_143 ();
 FILLCELL_X1 FILLER_54_180 ();
 FILLCELL_X16 FILLER_54_184 ();
 FILLCELL_X4 FILLER_54_200 ();
 FILLCELL_X2 FILLER_54_204 ();
 FILLCELL_X1 FILLER_54_206 ();
 FILLCELL_X2 FILLER_54_210 ();
 FILLCELL_X1 FILLER_54_212 ();
 FILLCELL_X8 FILLER_54_216 ();
 FILLCELL_X4 FILLER_54_224 ();
 FILLCELL_X2 FILLER_54_234 ();
 FILLCELL_X16 FILLER_54_239 ();
 FILLCELL_X8 FILLER_54_255 ();
 FILLCELL_X2 FILLER_54_263 ();
 FILLCELL_X1 FILLER_54_265 ();
 FILLCELL_X1 FILLER_54_269 ();
 FILLCELL_X1 FILLER_54_287 ();
 FILLCELL_X1 FILLER_54_292 ();
 FILLCELL_X1 FILLER_54_312 ();
 FILLCELL_X2 FILLER_54_332 ();
 FILLCELL_X2 FILLER_54_354 ();
 FILLCELL_X1 FILLER_54_356 ();
 FILLCELL_X1 FILLER_54_365 ();
 FILLCELL_X2 FILLER_54_370 ();
 FILLCELL_X8 FILLER_54_376 ();
 FILLCELL_X2 FILLER_54_384 ();
 FILLCELL_X1 FILLER_54_386 ();
 FILLCELL_X8 FILLER_54_408 ();
 FILLCELL_X2 FILLER_54_416 ();
 FILLCELL_X1 FILLER_54_418 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X2 FILLER_55_65 ();
 FILLCELL_X8 FILLER_55_70 ();
 FILLCELL_X4 FILLER_55_78 ();
 FILLCELL_X1 FILLER_55_82 ();
 FILLCELL_X4 FILLER_55_89 ();
 FILLCELL_X2 FILLER_55_93 ();
 FILLCELL_X8 FILLER_55_98 ();
 FILLCELL_X8 FILLER_55_118 ();
 FILLCELL_X4 FILLER_55_126 ();
 FILLCELL_X2 FILLER_55_142 ();
 FILLCELL_X1 FILLER_55_144 ();
 FILLCELL_X2 FILLER_55_178 ();
 FILLCELL_X1 FILLER_55_183 ();
 FILLCELL_X4 FILLER_55_187 ();
 FILLCELL_X1 FILLER_55_191 ();
 FILLCELL_X4 FILLER_55_195 ();
 FILLCELL_X1 FILLER_55_206 ();
 FILLCELL_X2 FILLER_55_210 ();
 FILLCELL_X1 FILLER_55_212 ();
 FILLCELL_X2 FILLER_55_216 ();
 FILLCELL_X1 FILLER_55_218 ();
 FILLCELL_X4 FILLER_55_222 ();
 FILLCELL_X2 FILLER_55_232 ();
 FILLCELL_X1 FILLER_55_234 ();
 FILLCELL_X2 FILLER_55_238 ();
 FILLCELL_X4 FILLER_55_243 ();
 FILLCELL_X2 FILLER_55_247 ();
 FILLCELL_X1 FILLER_55_252 ();
 FILLCELL_X4 FILLER_55_265 ();
 FILLCELL_X2 FILLER_55_275 ();
 FILLCELL_X2 FILLER_55_280 ();
 FILLCELL_X1 FILLER_55_282 ();
 FILLCELL_X2 FILLER_55_289 ();
 FILLCELL_X1 FILLER_55_291 ();
 FILLCELL_X2 FILLER_55_295 ();
 FILLCELL_X1 FILLER_55_297 ();
 FILLCELL_X1 FILLER_55_304 ();
 FILLCELL_X2 FILLER_55_308 ();
 FILLCELL_X1 FILLER_55_313 ();
 FILLCELL_X2 FILLER_55_317 ();
 FILLCELL_X16 FILLER_55_325 ();
 FILLCELL_X4 FILLER_55_341 ();
 FILLCELL_X1 FILLER_55_345 ();
 FILLCELL_X2 FILLER_55_355 ();
 FILLCELL_X1 FILLER_55_357 ();
 FILLCELL_X32 FILLER_55_378 ();
 FILLCELL_X8 FILLER_55_410 ();
 FILLCELL_X1 FILLER_55_418 ();
endmodule
