module johnson_counter (clk,
    enable,
    load_en,
    rst_n,
    count,
    load_val);
 input clk;
 input enable;
 input load_en;
 input rst_n;
 output [3:0] count;
 input [3:0] load_val;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X2 _22_ (.A(enable),
    .Z(_05_));
 OAI21_X1 _23_ (.A(net5),
    .B1(_05_),
    .B2(net6),
    .ZN(_06_));
 BUF_X4 _24_ (.A(load_en),
    .Z(_07_));
 MUX2_X1 _25_ (.A(_00_),
    .B(net1),
    .S(_07_),
    .Z(_08_));
 INV_X1 _26_ (.A(_08_),
    .ZN(_09_));
 AOI21_X1 _27_ (.A(_06_),
    .B1(_09_),
    .B2(_05_),
    .ZN(_01_));
 OAI21_X1 _28_ (.A(net5),
    .B1(_05_),
    .B2(net7),
    .ZN(_10_));
 MUX2_X1 _29_ (.A(net6),
    .B(net2),
    .S(_07_),
    .Z(_11_));
 INV_X1 _30_ (.A(_11_),
    .ZN(_12_));
 AOI21_X1 _31_ (.A(_10_),
    .B1(_12_),
    .B2(_05_),
    .ZN(_02_));
 OAI21_X1 _32_ (.A(net5),
    .B1(_05_),
    .B2(net8),
    .ZN(_13_));
 MUX2_X1 _33_ (.A(net7),
    .B(net3),
    .S(_07_),
    .Z(_14_));
 INV_X1 _34_ (.A(_14_),
    .ZN(_15_));
 AOI21_X1 _35_ (.A(_13_),
    .B1(_15_),
    .B2(_05_),
    .ZN(_03_));
 OAI21_X1 _36_ (.A(net5),
    .B1(net9),
    .B2(_05_),
    .ZN(_16_));
 MUX2_X1 _37_ (.A(net8),
    .B(net4),
    .S(_07_),
    .Z(_17_));
 INV_X1 _38_ (.A(_17_),
    .ZN(_18_));
 AOI21_X1 _39_ (.A(_16_),
    .B1(_18_),
    .B2(_05_),
    .ZN(_04_));
 DFF_X1 \count[0]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net6),
    .QN(_21_));
 DFF_X1 \count[1]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net7),
    .QN(_20_));
 DFF_X1 \count[2]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net8),
    .QN(_19_));
 DFF_X1 \count[3]$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net9),
    .QN(_00_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_91 ();
 BUF_X1 input1 (.A(load_val[0]),
    .Z(net1));
 BUF_X1 input2 (.A(load_val[1]),
    .Z(net2));
 BUF_X1 input3 (.A(load_val[2]),
    .Z(net3));
 BUF_X1 input4 (.A(load_val[3]),
    .Z(net4));
 BUF_X1 input5 (.A(rst_n),
    .Z(net5));
 BUF_X1 output6 (.A(net6),
    .Z(count[0]));
 BUF_X1 output7 (.A(net7),
    .Z(count[1]));
 BUF_X1 output8 (.A(net8),
    .Z(count[2]));
 BUF_X1 output9 (.A(net9),
    .Z(count[3]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X16 FILLER_0_321 ();
 FILLCELL_X4 FILLER_0_337 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X16 FILLER_1_321 ();
 FILLCELL_X4 FILLER_1_337 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X16 FILLER_2_321 ();
 FILLCELL_X4 FILLER_2_337 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X16 FILLER_3_321 ();
 FILLCELL_X4 FILLER_3_337 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X16 FILLER_4_321 ();
 FILLCELL_X4 FILLER_4_337 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X16 FILLER_5_321 ();
 FILLCELL_X4 FILLER_5_337 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X16 FILLER_6_321 ();
 FILLCELL_X4 FILLER_6_337 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X16 FILLER_7_321 ();
 FILLCELL_X4 FILLER_7_337 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X16 FILLER_8_321 ();
 FILLCELL_X4 FILLER_8_337 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X16 FILLER_9_321 ();
 FILLCELL_X4 FILLER_9_337 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X16 FILLER_10_321 ();
 FILLCELL_X4 FILLER_10_337 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X16 FILLER_11_321 ();
 FILLCELL_X4 FILLER_11_337 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X16 FILLER_12_321 ();
 FILLCELL_X4 FILLER_12_337 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X16 FILLER_13_321 ();
 FILLCELL_X4 FILLER_13_337 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X16 FILLER_14_321 ();
 FILLCELL_X4 FILLER_14_337 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X16 FILLER_15_321 ();
 FILLCELL_X4 FILLER_15_337 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X16 FILLER_16_321 ();
 FILLCELL_X4 FILLER_16_337 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X16 FILLER_17_321 ();
 FILLCELL_X4 FILLER_17_337 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X16 FILLER_18_321 ();
 FILLCELL_X4 FILLER_18_337 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X16 FILLER_19_321 ();
 FILLCELL_X4 FILLER_19_337 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X16 FILLER_20_321 ();
 FILLCELL_X4 FILLER_20_337 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X16 FILLER_21_321 ();
 FILLCELL_X4 FILLER_21_337 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X8 FILLER_22_17 ();
 FILLCELL_X1 FILLER_22_25 ();
 FILLCELL_X32 FILLER_22_29 ();
 FILLCELL_X32 FILLER_22_61 ();
 FILLCELL_X32 FILLER_22_93 ();
 FILLCELL_X32 FILLER_22_125 ();
 FILLCELL_X32 FILLER_22_157 ();
 FILLCELL_X8 FILLER_22_189 ();
 FILLCELL_X32 FILLER_22_204 ();
 FILLCELL_X32 FILLER_22_236 ();
 FILLCELL_X32 FILLER_22_268 ();
 FILLCELL_X8 FILLER_22_300 ();
 FILLCELL_X4 FILLER_22_308 ();
 FILLCELL_X2 FILLER_22_312 ();
 FILLCELL_X1 FILLER_22_314 ();
 FILLCELL_X16 FILLER_22_318 ();
 FILLCELL_X4 FILLER_22_334 ();
 FILLCELL_X2 FILLER_22_338 ();
 FILLCELL_X1 FILLER_22_340 ();
 FILLCELL_X16 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_17 ();
 FILLCELL_X32 FILLER_23_22 ();
 FILLCELL_X32 FILLER_23_54 ();
 FILLCELL_X32 FILLER_23_86 ();
 FILLCELL_X32 FILLER_23_118 ();
 FILLCELL_X32 FILLER_23_150 ();
 FILLCELL_X8 FILLER_23_182 ();
 FILLCELL_X2 FILLER_23_190 ();
 FILLCELL_X32 FILLER_23_201 ();
 FILLCELL_X32 FILLER_23_233 ();
 FILLCELL_X32 FILLER_23_265 ();
 FILLCELL_X16 FILLER_23_297 ();
 FILLCELL_X8 FILLER_23_313 ();
 FILLCELL_X1 FILLER_23_321 ();
 FILLCELL_X16 FILLER_23_325 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X16 FILLER_24_129 ();
 FILLCELL_X8 FILLER_24_145 ();
 FILLCELL_X4 FILLER_24_153 ();
 FILLCELL_X2 FILLER_24_157 ();
 FILLCELL_X1 FILLER_24_159 ();
 FILLCELL_X2 FILLER_24_167 ();
 FILLCELL_X32 FILLER_24_199 ();
 FILLCELL_X32 FILLER_24_231 ();
 FILLCELL_X32 FILLER_24_263 ();
 FILLCELL_X32 FILLER_24_295 ();
 FILLCELL_X8 FILLER_24_327 ();
 FILLCELL_X4 FILLER_24_335 ();
 FILLCELL_X2 FILLER_24_339 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X4 FILLER_25_161 ();
 FILLCELL_X4 FILLER_25_182 ();
 FILLCELL_X32 FILLER_25_190 ();
 FILLCELL_X32 FILLER_25_222 ();
 FILLCELL_X32 FILLER_25_254 ();
 FILLCELL_X32 FILLER_25_286 ();
 FILLCELL_X4 FILLER_25_318 ();
 FILLCELL_X2 FILLER_25_322 ();
 FILLCELL_X8 FILLER_25_327 ();
 FILLCELL_X4 FILLER_25_335 ();
 FILLCELL_X2 FILLER_25_339 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X4 FILLER_26_161 ();
 FILLCELL_X1 FILLER_26_165 ();
 FILLCELL_X16 FILLER_26_168 ();
 FILLCELL_X2 FILLER_26_188 ();
 FILLCELL_X1 FILLER_26_190 ();
 FILLCELL_X32 FILLER_26_200 ();
 FILLCELL_X32 FILLER_26_232 ();
 FILLCELL_X32 FILLER_26_264 ();
 FILLCELL_X32 FILLER_26_296 ();
 FILLCELL_X8 FILLER_26_328 ();
 FILLCELL_X4 FILLER_26_336 ();
 FILLCELL_X1 FILLER_26_340 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X4 FILLER_27_161 ();
 FILLCELL_X2 FILLER_27_165 ();
 FILLCELL_X1 FILLER_27_167 ();
 FILLCELL_X32 FILLER_27_176 ();
 FILLCELL_X32 FILLER_27_208 ();
 FILLCELL_X32 FILLER_27_240 ();
 FILLCELL_X32 FILLER_27_272 ();
 FILLCELL_X32 FILLER_27_304 ();
 FILLCELL_X4 FILLER_27_336 ();
 FILLCELL_X1 FILLER_27_340 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X2 FILLER_28_161 ();
 FILLCELL_X1 FILLER_28_180 ();
 FILLCELL_X32 FILLER_28_186 ();
 FILLCELL_X32 FILLER_28_218 ();
 FILLCELL_X32 FILLER_28_250 ();
 FILLCELL_X32 FILLER_28_282 ();
 FILLCELL_X16 FILLER_28_314 ();
 FILLCELL_X8 FILLER_28_330 ();
 FILLCELL_X2 FILLER_28_338 ();
 FILLCELL_X1 FILLER_28_340 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X16 FILLER_29_321 ();
 FILLCELL_X4 FILLER_29_337 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X16 FILLER_30_161 ();
 FILLCELL_X4 FILLER_30_177 ();
 FILLCELL_X32 FILLER_30_185 ();
 FILLCELL_X32 FILLER_30_217 ();
 FILLCELL_X32 FILLER_30_249 ();
 FILLCELL_X32 FILLER_30_281 ();
 FILLCELL_X16 FILLER_30_313 ();
 FILLCELL_X8 FILLER_30_329 ();
 FILLCELL_X4 FILLER_30_337 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X4 FILLER_31_161 ();
 FILLCELL_X2 FILLER_31_165 ();
 FILLCELL_X1 FILLER_31_176 ();
 FILLCELL_X32 FILLER_31_181 ();
 FILLCELL_X32 FILLER_31_213 ();
 FILLCELL_X32 FILLER_31_245 ();
 FILLCELL_X32 FILLER_31_277 ();
 FILLCELL_X32 FILLER_31_309 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X4 FILLER_32_161 ();
 FILLCELL_X4 FILLER_32_169 ();
 FILLCELL_X2 FILLER_32_173 ();
 FILLCELL_X1 FILLER_32_175 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X16 FILLER_32_321 ();
 FILLCELL_X4 FILLER_32_337 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X8 FILLER_33_161 ();
 FILLCELL_X4 FILLER_33_169 ();
 FILLCELL_X2 FILLER_33_173 ();
 FILLCELL_X32 FILLER_33_180 ();
 FILLCELL_X32 FILLER_33_212 ();
 FILLCELL_X32 FILLER_33_244 ();
 FILLCELL_X32 FILLER_33_276 ();
 FILLCELL_X32 FILLER_33_308 ();
 FILLCELL_X1 FILLER_33_340 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X16 FILLER_34_321 ();
 FILLCELL_X4 FILLER_34_337 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X16 FILLER_35_321 ();
 FILLCELL_X4 FILLER_35_337 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X16 FILLER_36_321 ();
 FILLCELL_X4 FILLER_36_337 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X16 FILLER_37_321 ();
 FILLCELL_X4 FILLER_37_337 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X16 FILLER_38_321 ();
 FILLCELL_X4 FILLER_38_337 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X16 FILLER_39_321 ();
 FILLCELL_X4 FILLER_39_337 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X16 FILLER_40_321 ();
 FILLCELL_X4 FILLER_40_337 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X16 FILLER_41_321 ();
 FILLCELL_X4 FILLER_41_337 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X16 FILLER_42_321 ();
 FILLCELL_X4 FILLER_42_337 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X16 FILLER_43_321 ();
 FILLCELL_X4 FILLER_43_337 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X16 FILLER_44_321 ();
 FILLCELL_X4 FILLER_44_337 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X1 FILLER_45_161 ();
 FILLCELL_X2 FILLER_45_165 ();
 FILLCELL_X1 FILLER_45_167 ();
 FILLCELL_X8 FILLER_45_171 ();
 FILLCELL_X1 FILLER_45_179 ();
 FILLCELL_X1 FILLER_45_183 ();
 FILLCELL_X32 FILLER_45_187 ();
 FILLCELL_X32 FILLER_45_219 ();
 FILLCELL_X32 FILLER_45_251 ();
 FILLCELL_X32 FILLER_45_283 ();
 FILLCELL_X16 FILLER_45_315 ();
 FILLCELL_X8 FILLER_45_331 ();
 FILLCELL_X2 FILLER_45_339 ();
endmodule
