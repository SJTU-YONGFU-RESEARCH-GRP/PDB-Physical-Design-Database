module parameterized_sync_reset_counter (clk,
    enable,
    sync_rst,
    tc,
    count);
 input clk;
 input enable;
 input sync_rst;
 output tc;
 output [7:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _34_ (.I(net1),
    .ZN(_08_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _35_ (.A1(net3),
    .A2(_08_),
    .ZN(_09_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _36_ (.A1(net6),
    .A2(net8),
    .A3(net7),
    .A4(net9),
    .Z(_10_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _37_ (.A1(net5),
    .A2(_32_),
    .A3(net10),
    .A4(_10_),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _38_ (.A1(net3),
    .A2(_08_),
    .A3(net2),
    .Z(_11_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _39_ (.A1(net2),
    .A2(_09_),
    .B1(net11),
    .B2(_11_),
    .ZN(_00_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _40_ (.I(net2),
    .ZN(_12_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _41_ (.I0(net4),
    .I1(_33_),
    .S(net1),
    .Z(_13_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _42_ (.A1(_12_),
    .A2(_13_),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _43_ (.A1(_32_),
    .A2(net1),
    .Z(_14_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _44_ (.A1(net5),
    .A2(_14_),
    .ZN(_15_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _45_ (.A1(net2),
    .A2(_15_),
    .ZN(_02_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _46_ (.A1(net10),
    .A2(_10_),
    .Z(_16_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _47_ (.A1(net5),
    .A2(_14_),
    .Z(_17_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _48_ (.A1(net5),
    .A2(net3),
    .A3(net4),
    .A4(net1),
    .Z(_18_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _49_ (.A1(net6),
    .A2(_18_),
    .ZN(_19_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _50_ (.A1(_16_),
    .A2(_17_),
    .B(_19_),
    .C(net2),
    .ZN(_03_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _51_ (.A1(net6),
    .A2(net5),
    .A3(_32_),
    .A4(net1),
    .Z(_20_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _52_ (.A1(net7),
    .A2(_20_),
    .Z(_21_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _53_ (.A1(_12_),
    .A2(_21_),
    .Z(_04_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _54_ (.A1(net6),
    .A2(net7),
    .ZN(_22_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _55_ (.A1(net5),
    .A2(net3),
    .A3(net4),
    .A4(net1),
    .ZN(_23_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _56_ (.A1(_22_),
    .A2(_23_),
    .B(net8),
    .ZN(_24_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _57_ (.A1(net8),
    .A2(_22_),
    .A3(_23_),
    .Z(_25_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _58_ (.A1(_16_),
    .A2(_17_),
    .B1(_24_),
    .B2(_25_),
    .C(net2),
    .ZN(_05_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _59_ (.A1(net6),
    .A2(net8),
    .A3(net7),
    .ZN(_26_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _60_ (.A1(net5),
    .A2(_32_),
    .A3(net1),
    .ZN(_27_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _61_ (.A1(_26_),
    .A2(_27_),
    .B(net9),
    .ZN(_28_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _62_ (.A1(net9),
    .A2(_26_),
    .A3(_27_),
    .Z(_29_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _63_ (.A1(_28_),
    .A2(_29_),
    .B(net2),
    .ZN(_06_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _64_ (.A1(_27_),
    .A2(_23_),
    .ZN(_30_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _65_ (.A1(_10_),
    .A2(_18_),
    .B(net10),
    .ZN(_31_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _66_ (.A1(_16_),
    .A2(_30_),
    .B(_31_),
    .C(net2),
    .ZN(_07_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _67_ (.A(net3),
    .B(net4),
    .CO(_32_),
    .S(_33_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter_reg[0]$_SDFFE_PP0P_  (.D(_00_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net3));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter_reg[1]$_SDFFE_PP0P_  (.D(_01_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter_reg[2]$_SDFFE_PP0P_  (.D(_02_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter_reg[3]$_SDFFE_PP0P_  (.D(_03_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter_reg[4]$_SDFFE_PP0P_  (.D(_04_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter_reg[5]$_SDFFE_PP0P_  (.D(_05_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net8));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter_reg[6]$_SDFFE_PP0P_  (.D(_06_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net9));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter_reg[7]$_SDFFE_PP0P_  (.D(_07_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net10));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_67 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input1 (.I(enable),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input2 (.I(sync_rst),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output3 (.I(net3),
    .Z(count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output4 (.I(net4),
    .Z(count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output5 (.I(net5),
    .Z(count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output6 (.I(net6),
    .Z(count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output7 (.I(net7),
    .Z(count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output8 (.I(net8),
    .Z(count[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output9 (.I(net9),
    .Z(count[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output10 (.I(net10),
    .Z(count[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output11 (.I(net11),
    .Z(tc));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_248 ();
endmodule
