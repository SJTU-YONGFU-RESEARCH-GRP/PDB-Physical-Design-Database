module gpio_controller (clk,
    int_out,
    rst_n,
    gpio_dir,
    gpio_in,
    gpio_out,
    gpio_pins,
    int_clear,
    int_enable,
    int_polarity,
    int_status,
    int_type);
 input clk;
 output int_out;
 input rst_n;
 input [31:0] gpio_dir;
 output [31:0] gpio_in;
 input [31:0] gpio_out;
 inout [31:0] gpio_pins;
 input [31:0] int_clear;
 input [31:0] int_enable;
 input [31:0] int_polarity;
 output [31:0] int_status;
 input [31:0] int_type;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire \gpio_in_prev[0] ;
 wire \gpio_in_prev[10] ;
 wire \gpio_in_prev[11] ;
 wire \gpio_in_prev[12] ;
 wire \gpio_in_prev[13] ;
 wire \gpio_in_prev[14] ;
 wire \gpio_in_prev[15] ;
 wire \gpio_in_prev[16] ;
 wire \gpio_in_prev[17] ;
 wire \gpio_in_prev[18] ;
 wire \gpio_in_prev[19] ;
 wire \gpio_in_prev[1] ;
 wire \gpio_in_prev[20] ;
 wire \gpio_in_prev[21] ;
 wire \gpio_in_prev[22] ;
 wire \gpio_in_prev[23] ;
 wire \gpio_in_prev[24] ;
 wire \gpio_in_prev[25] ;
 wire \gpio_in_prev[26] ;
 wire \gpio_in_prev[27] ;
 wire \gpio_in_prev[28] ;
 wire \gpio_in_prev[29] ;
 wire \gpio_in_prev[2] ;
 wire \gpio_in_prev[30] ;
 wire \gpio_in_prev[31] ;
 wire \gpio_in_prev[3] ;
 wire \gpio_in_prev[4] ;
 wire \gpio_in_prev[5] ;
 wire \gpio_in_prev[6] ;
 wire \gpio_in_prev[7] ;
 wire \gpio_in_prev[8] ;
 wire \gpio_in_prev[9] ;
 wire \gpio_in_sync1[0] ;
 wire \gpio_in_sync1[10] ;
 wire \gpio_in_sync1[11] ;
 wire \gpio_in_sync1[12] ;
 wire \gpio_in_sync1[13] ;
 wire \gpio_in_sync1[14] ;
 wire \gpio_in_sync1[15] ;
 wire \gpio_in_sync1[16] ;
 wire \gpio_in_sync1[17] ;
 wire \gpio_in_sync1[18] ;
 wire \gpio_in_sync1[19] ;
 wire \gpio_in_sync1[1] ;
 wire \gpio_in_sync1[20] ;
 wire \gpio_in_sync1[21] ;
 wire \gpio_in_sync1[22] ;
 wire \gpio_in_sync1[23] ;
 wire \gpio_in_sync1[24] ;
 wire \gpio_in_sync1[25] ;
 wire \gpio_in_sync1[26] ;
 wire \gpio_in_sync1[27] ;
 wire \gpio_in_sync1[28] ;
 wire \gpio_in_sync1[29] ;
 wire \gpio_in_sync1[2] ;
 wire \gpio_in_sync1[30] ;
 wire \gpio_in_sync1[31] ;
 wire \gpio_in_sync1[3] ;
 wire \gpio_in_sync1[4] ;
 wire \gpio_in_sync1[5] ;
 wire \gpio_in_sync1[6] ;
 wire \gpio_in_sync1[7] ;
 wire \gpio_in_sync1[8] ;
 wire \gpio_in_sync1[9] ;
 wire \gpio_in_sync2[0] ;
 wire \gpio_in_sync2[10] ;
 wire \gpio_in_sync2[11] ;
 wire \gpio_in_sync2[12] ;
 wire \gpio_in_sync2[13] ;
 wire \gpio_in_sync2[14] ;
 wire \gpio_in_sync2[15] ;
 wire \gpio_in_sync2[16] ;
 wire \gpio_in_sync2[17] ;
 wire \gpio_in_sync2[18] ;
 wire \gpio_in_sync2[19] ;
 wire \gpio_in_sync2[1] ;
 wire \gpio_in_sync2[20] ;
 wire \gpio_in_sync2[21] ;
 wire \gpio_in_sync2[22] ;
 wire \gpio_in_sync2[23] ;
 wire \gpio_in_sync2[24] ;
 wire \gpio_in_sync2[25] ;
 wire \gpio_in_sync2[26] ;
 wire \gpio_in_sync2[27] ;
 wire \gpio_in_sync2[28] ;
 wire \gpio_in_sync2[29] ;
 wire \gpio_in_sync2[2] ;
 wire \gpio_in_sync2[30] ;
 wire \gpio_in_sync2[31] ;
 wire \gpio_in_sync2[3] ;
 wire \gpio_in_sync2[4] ;
 wire \gpio_in_sync2[5] ;
 wire \gpio_in_sync2[6] ;
 wire \gpio_in_sync2[7] ;
 wire \gpio_in_sync2[8] ;
 wire \gpio_in_sync2[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net227;

 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _212_ (.A1(\gpio_in_sync2[0] ),
    .A2(\gpio_in_prev[0] ),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _213_ (.A1(net130),
    .A2(_032_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _214_ (.A1(\gpio_in_sync2[0] ),
    .A2(net98),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _215_ (.A1(net66),
    .A2(_034_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _216_ (.A1(_033_),
    .A2(_035_),
    .B(net195),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _217_ (.A1(net34),
    .A2(_036_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _218_ (.I(net196),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _219_ (.A1(\gpio_in_prev[10] ),
    .A2(net131),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _220_ (.A1(\gpio_in_sync2[10] ),
    .A2(net99),
    .A3(_038_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _221_ (.I(\gpio_in_prev[10] ),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _222_ (.A1(_040_),
    .A2(net131),
    .B(net99),
    .C(\gpio_in_sync2[10] ),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _223_ (.A1(_039_),
    .A2(_041_),
    .B(net67),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _224_ (.A1(_037_),
    .A2(_042_),
    .B(net35),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _225_ (.I(net197),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _226_ (.A1(\gpio_in_prev[11] ),
    .A2(net132),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _227_ (.A1(\gpio_in_sync2[11] ),
    .A2(net100),
    .A3(_044_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _228_ (.I(\gpio_in_prev[11] ),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _229_ (.A1(_046_),
    .A2(net132),
    .B(net100),
    .C(\gpio_in_sync2[11] ),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _230_ (.A1(_045_),
    .A2(_047_),
    .B(net68),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _231_ (.A1(_043_),
    .A2(_048_),
    .B(net36),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _232_ (.I(net198),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _233_ (.A1(\gpio_in_prev[12] ),
    .A2(net133),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _234_ (.A1(\gpio_in_sync2[12] ),
    .A2(net101),
    .A3(_050_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _235_ (.I(\gpio_in_prev[12] ),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _236_ (.A1(_052_),
    .A2(net133),
    .B(net101),
    .C(\gpio_in_sync2[12] ),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _237_ (.A1(_051_),
    .A2(_053_),
    .B(net69),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _238_ (.A1(_049_),
    .A2(_054_),
    .B(net37),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _239_ (.I(net199),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _240_ (.A1(\gpio_in_prev[13] ),
    .A2(net134),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _241_ (.A1(\gpio_in_sync2[13] ),
    .A2(net102),
    .A3(_056_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _242_ (.I(\gpio_in_prev[13] ),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _243_ (.A1(_058_),
    .A2(net134),
    .B(net102),
    .C(\gpio_in_sync2[13] ),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _244_ (.A1(_057_),
    .A2(_059_),
    .B(net70),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _245_ (.A1(_055_),
    .A2(_060_),
    .B(net38),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _246_ (.I(net200),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _247_ (.A1(net135),
    .A2(\gpio_in_prev[14] ),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _248_ (.A1(\gpio_in_sync2[14] ),
    .A2(net103),
    .A3(_062_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _249_ (.I(\gpio_in_prev[14] ),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _250_ (.A1(net135),
    .A2(_064_),
    .B(\gpio_in_sync2[14] ),
    .C(net103),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _251_ (.A1(_063_),
    .A2(_065_),
    .B(net71),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _252_ (.A1(_061_),
    .A2(_066_),
    .B(net39),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _253_ (.I(net201),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _254_ (.A1(net136),
    .A2(\gpio_in_prev[15] ),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _255_ (.A1(\gpio_in_sync2[15] ),
    .A2(net104),
    .A3(_068_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _256_ (.I(\gpio_in_prev[15] ),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _257_ (.A1(net136),
    .A2(_070_),
    .B(\gpio_in_sync2[15] ),
    .C(net104),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _258_ (.A1(_069_),
    .A2(_071_),
    .B(net72),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _259_ (.A1(_067_),
    .A2(_072_),
    .B(net40),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _260_ (.I(net202),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _261_ (.A1(net137),
    .A2(\gpio_in_prev[16] ),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _262_ (.A1(\gpio_in_sync2[16] ),
    .A2(net105),
    .A3(_074_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _263_ (.I(\gpio_in_prev[16] ),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _264_ (.A1(net137),
    .A2(_076_),
    .B(\gpio_in_sync2[16] ),
    .C(net105),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _265_ (.A1(_075_),
    .A2(_077_),
    .B(net73),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _266_ (.A1(_073_),
    .A2(_078_),
    .B(net41),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _267_ (.A1(\gpio_in_sync2[17] ),
    .A2(\gpio_in_prev[17] ),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _268_ (.A1(net138),
    .A2(_079_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _269_ (.A1(\gpio_in_sync2[17] ),
    .A2(net106),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _270_ (.A1(net74),
    .A2(_081_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _271_ (.A1(_080_),
    .A2(_082_),
    .B(net203),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _272_ (.A1(net42),
    .A2(_083_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _273_ (.A1(\gpio_in_sync2[18] ),
    .A2(\gpio_in_prev[18] ),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _274_ (.A1(net139),
    .A2(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _275_ (.A1(\gpio_in_sync2[18] ),
    .A2(net107),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _276_ (.A1(net75),
    .A2(_086_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _277_ (.A1(_085_),
    .A2(_087_),
    .B(net204),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _278_ (.A1(net43),
    .A2(_088_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _279_ (.A1(\gpio_in_sync2[19] ),
    .A2(\gpio_in_prev[19] ),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _280_ (.A1(net140),
    .A2(_089_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _281_ (.A1(\gpio_in_sync2[19] ),
    .A2(net108),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _282_ (.A1(net76),
    .A2(_091_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _283_ (.A1(_090_),
    .A2(_092_),
    .B(net205),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _284_ (.A1(net44),
    .A2(_093_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _285_ (.A1(\gpio_in_sync2[1] ),
    .A2(\gpio_in_prev[1] ),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _286_ (.A1(net141),
    .A2(_094_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _287_ (.A1(\gpio_in_sync2[1] ),
    .A2(net109),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _288_ (.A1(net77),
    .A2(_096_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _289_ (.A1(_095_),
    .A2(_097_),
    .B(net206),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _290_ (.A1(net45),
    .A2(_098_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _291_ (.A1(\gpio_in_sync2[20] ),
    .A2(\gpio_in_prev[20] ),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _292_ (.A1(net142),
    .A2(_099_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _293_ (.A1(\gpio_in_sync2[20] ),
    .A2(net110),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _294_ (.A1(net78),
    .A2(_101_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _295_ (.A1(_100_),
    .A2(_102_),
    .B(net207),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _296_ (.A1(net46),
    .A2(_103_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _297_ (.A1(\gpio_in_sync2[21] ),
    .A2(\gpio_in_prev[21] ),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _298_ (.A1(net143),
    .A2(_104_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _299_ (.A1(\gpio_in_sync2[21] ),
    .A2(net111),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _300_ (.A1(net79),
    .A2(_106_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _301_ (.A1(_105_),
    .A2(_107_),
    .B(net208),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _302_ (.A1(net47),
    .A2(_108_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _303_ (.A1(\gpio_in_sync2[22] ),
    .A2(\gpio_in_prev[22] ),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _304_ (.A1(net144),
    .A2(_109_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _305_ (.A1(\gpio_in_sync2[22] ),
    .A2(net112),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _306_ (.A1(net80),
    .A2(_111_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _307_ (.A1(_110_),
    .A2(_112_),
    .B(net209),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _308_ (.A1(net48),
    .A2(_113_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _309_ (.A1(\gpio_in_sync2[23] ),
    .A2(\gpio_in_prev[23] ),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _310_ (.A1(net145),
    .A2(_114_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _311_ (.A1(\gpio_in_sync2[23] ),
    .A2(net113),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _312_ (.A1(net81),
    .A2(_116_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _313_ (.A1(_115_),
    .A2(_117_),
    .B(net210),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _314_ (.A1(net49),
    .A2(_118_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _315_ (.A1(\gpio_in_sync2[24] ),
    .A2(\gpio_in_prev[24] ),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _316_ (.A1(net146),
    .A2(_119_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _317_ (.A1(\gpio_in_sync2[24] ),
    .A2(net114),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _318_ (.A1(net82),
    .A2(_121_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _319_ (.A1(_120_),
    .A2(_122_),
    .B(net211),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _320_ (.A1(net50),
    .A2(_123_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _321_ (.A1(\gpio_in_sync2[25] ),
    .A2(\gpio_in_prev[25] ),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _322_ (.A1(net147),
    .A2(_124_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _323_ (.A1(\gpio_in_sync2[25] ),
    .A2(net115),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _324_ (.A1(net83),
    .A2(_126_),
    .Z(_127_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _325_ (.A1(_125_),
    .A2(_127_),
    .B(net212),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _326_ (.A1(net51),
    .A2(_128_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _327_ (.A1(\gpio_in_sync2[26] ),
    .A2(\gpio_in_prev[26] ),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _328_ (.A1(net148),
    .A2(_129_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _329_ (.A1(\gpio_in_sync2[26] ),
    .A2(net116),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _330_ (.A1(net84),
    .A2(_131_),
    .Z(_132_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _331_ (.A1(_130_),
    .A2(_132_),
    .B(net213),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _332_ (.A1(net52),
    .A2(_133_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _333_ (.A1(\gpio_in_sync2[27] ),
    .A2(\gpio_in_prev[27] ),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _334_ (.A1(net149),
    .A2(_134_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _335_ (.A1(\gpio_in_sync2[27] ),
    .A2(net117),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _336_ (.A1(net85),
    .A2(_136_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _337_ (.A1(_135_),
    .A2(_137_),
    .B(net214),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _338_ (.A1(net53),
    .A2(_138_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _339_ (.A1(\gpio_in_sync2[28] ),
    .A2(\gpio_in_prev[28] ),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _340_ (.A1(net150),
    .A2(_139_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _341_ (.A1(\gpio_in_sync2[28] ),
    .A2(net118),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _342_ (.A1(net86),
    .A2(_141_),
    .Z(_142_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _343_ (.A1(_140_),
    .A2(_142_),
    .B(net215),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _344_ (.A1(net54),
    .A2(_143_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _345_ (.A1(\gpio_in_sync2[29] ),
    .A2(\gpio_in_prev[29] ),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _346_ (.A1(net151),
    .A2(_144_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _347_ (.A1(\gpio_in_sync2[29] ),
    .A2(net119),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _348_ (.A1(net87),
    .A2(_146_),
    .Z(_147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _349_ (.A1(_145_),
    .A2(_147_),
    .B(net216),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _350_ (.A1(net55),
    .A2(_148_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _351_ (.A1(\gpio_in_sync2[2] ),
    .A2(\gpio_in_prev[2] ),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _352_ (.A1(net152),
    .A2(_149_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _353_ (.A1(\gpio_in_sync2[2] ),
    .A2(net120),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _354_ (.A1(net88),
    .A2(_151_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _355_ (.A1(_150_),
    .A2(_152_),
    .B(net217),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _356_ (.A1(net56),
    .A2(_153_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _357_ (.A1(\gpio_in_sync2[30] ),
    .A2(\gpio_in_prev[30] ),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _358_ (.A1(net153),
    .A2(_154_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _359_ (.A1(\gpio_in_sync2[30] ),
    .A2(net121),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _360_ (.A1(net89),
    .A2(_156_),
    .Z(_157_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _361_ (.A1(_155_),
    .A2(_157_),
    .B(net218),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _362_ (.A1(net57),
    .A2(_158_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _363_ (.A1(\gpio_in_sync2[31] ),
    .A2(\gpio_in_prev[31] ),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _364_ (.A1(net154),
    .A2(_159_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _365_ (.A1(\gpio_in_sync2[31] ),
    .A2(net122),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _366_ (.A1(net90),
    .A2(_161_),
    .Z(_162_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _367_ (.A1(_160_),
    .A2(_162_),
    .B(net219),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _368_ (.A1(net58),
    .A2(_163_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _369_ (.A1(\gpio_in_sync2[3] ),
    .A2(\gpio_in_prev[3] ),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _370_ (.A1(net155),
    .A2(_164_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _371_ (.A1(\gpio_in_sync2[3] ),
    .A2(net123),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _372_ (.A1(net91),
    .A2(_166_),
    .Z(_167_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _373_ (.A1(_165_),
    .A2(_167_),
    .B(net220),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _374_ (.A1(net59),
    .A2(_168_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _375_ (.A1(\gpio_in_sync2[4] ),
    .A2(\gpio_in_prev[4] ),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _376_ (.A1(net156),
    .A2(_169_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _377_ (.A1(\gpio_in_sync2[4] ),
    .A2(net124),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _378_ (.A1(net92),
    .A2(_171_),
    .Z(_172_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _379_ (.A1(_170_),
    .A2(_172_),
    .B(net221),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _380_ (.A1(net60),
    .A2(_173_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _381_ (.A1(\gpio_in_sync2[5] ),
    .A2(\gpio_in_prev[5] ),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _382_ (.A1(net157),
    .A2(_174_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _383_ (.A1(\gpio_in_sync2[5] ),
    .A2(net125),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _384_ (.A1(net93),
    .A2(_176_),
    .Z(_177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _385_ (.A1(_175_),
    .A2(_177_),
    .B(net222),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _386_ (.A1(net61),
    .A2(_178_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _387_ (.A1(\gpio_in_sync2[6] ),
    .A2(\gpio_in_prev[6] ),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _388_ (.A1(net158),
    .A2(_179_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _389_ (.A1(\gpio_in_sync2[6] ),
    .A2(net126),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _390_ (.A1(net94),
    .A2(_181_),
    .Z(_182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _391_ (.A1(_180_),
    .A2(_182_),
    .B(net223),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _392_ (.A1(net62),
    .A2(_183_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _393_ (.I(net224),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _394_ (.A1(net159),
    .A2(\gpio_in_prev[7] ),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _395_ (.A1(\gpio_in_sync2[7] ),
    .A2(net127),
    .A3(_185_),
    .Z(_186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _396_ (.I(\gpio_in_prev[7] ),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _397_ (.A1(net159),
    .A2(_187_),
    .B(\gpio_in_sync2[7] ),
    .C(net127),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _398_ (.A1(_186_),
    .A2(_188_),
    .B(net95),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _399_ (.A1(_184_),
    .A2(_189_),
    .B(net63),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _400_ (.I(net225),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _401_ (.A1(net160),
    .A2(\gpio_in_prev[8] ),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _402_ (.A1(\gpio_in_sync2[8] ),
    .A2(net128),
    .A3(_191_),
    .Z(_192_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _403_ (.I(\gpio_in_prev[8] ),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _404_ (.A1(net160),
    .A2(_193_),
    .B(\gpio_in_sync2[8] ),
    .C(net128),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _405_ (.A1(_192_),
    .A2(_194_),
    .B(net96),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _406_ (.A1(_190_),
    .A2(_195_),
    .B(net64),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _407_ (.I(net226),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _408_ (.A1(net161),
    .A2(\gpio_in_prev[9] ),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _409_ (.A1(\gpio_in_sync2[9] ),
    .A2(net129),
    .A3(_197_),
    .Z(_198_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _410_ (.I(\gpio_in_prev[9] ),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _411_ (.A1(net161),
    .A2(_199_),
    .B(\gpio_in_sync2[9] ),
    .C(net129),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _412_ (.A1(_198_),
    .A2(_200_),
    .B(net97),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _413_ (.A1(_196_),
    .A2(_201_),
    .B(net65),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _414_ (.A1(net203),
    .A2(net207),
    .A3(net210),
    .A4(net209),
    .Z(_202_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _415_ (.A1(net202),
    .A2(net205),
    .A3(net204),
    .A4(net208),
    .Z(_203_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _416_ (.A1(net212),
    .A2(net215),
    .A3(net219),
    .A4(net218),
    .Z(_204_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _417_ (.A1(net211),
    .A2(net214),
    .A3(net213),
    .A4(net216),
    .Z(_205_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _418_ (.A1(_202_),
    .A2(_203_),
    .A3(_204_),
    .A4(_205_),
    .Z(_206_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _419_ (.A1(net222),
    .A2(net221),
    .A3(net224),
    .A4(net200),
    .Z(_207_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _420_ (.A1(net206),
    .A2(net195),
    .A3(net220),
    .A4(net217),
    .Z(_208_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _421_ (.A1(net223),
    .A2(net199),
    .A3(net198),
    .A4(net201),
    .Z(_209_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _422_ (.A1(net226),
    .A2(net225),
    .A3(net197),
    .A4(net196),
    .Z(_210_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _423_ (.A1(_207_),
    .A2(_208_),
    .A3(_209_),
    .A4(_210_),
    .Z(_211_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _424_ (.A1(_206_),
    .A2(_211_),
    .Z(net194));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _425_ (.I(net2),
    .Z(net162));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _426_ (.I(net13),
    .Z(net173));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _427_ (.I(net24),
    .Z(net184));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _428_ (.I(net27),
    .Z(net187));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _429_ (.I(net28),
    .Z(net188));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _430_ (.I(net29),
    .Z(net189));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _431_ (.I(net30),
    .Z(net190));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _432_ (.I(net31),
    .Z(net191));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _433_ (.I(net32),
    .Z(net192));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _434_ (.I(net33),
    .Z(net193));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _435_ (.I(net3),
    .Z(net163));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _436_ (.I(net4),
    .Z(net164));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _437_ (.I(net5),
    .Z(net165));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _438_ (.I(net6),
    .Z(net166));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _439_ (.I(net7),
    .Z(net167));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _440_ (.I(net8),
    .Z(net168));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _441_ (.I(net9),
    .Z(net169));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _442_ (.I(net10),
    .Z(net170));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _443_ (.I(net11),
    .Z(net171));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _444_ (.I(net12),
    .Z(net172));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _445_ (.I(net14),
    .Z(net174));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _446_ (.I(net15),
    .Z(net175));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _447_ (.I(net16),
    .Z(net176));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _448_ (.I(net17),
    .Z(net177));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _449_ (.I(net18),
    .Z(net178));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _450_ (.I(net19),
    .Z(net179));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _451_ (.I(net20),
    .Z(net180));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _452_ (.I(net21),
    .Z(net181));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _453_ (.I(net22),
    .Z(net182));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _454_ (.I(net23),
    .Z(net183));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _455_ (.I(net25),
    .Z(net185));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _456_ (.I(net26),
    .Z(net186));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _457_ (.I(net2),
    .Z(gpio_pins[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _458_ (.I(net13),
    .Z(gpio_pins[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _459_ (.I(net24),
    .Z(gpio_pins[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _460_ (.I(net27),
    .Z(gpio_pins[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _461_ (.I(net28),
    .Z(gpio_pins[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _462_ (.I(net29),
    .Z(gpio_pins[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _463_ (.I(net30),
    .Z(gpio_pins[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _464_ (.I(net31),
    .Z(gpio_pins[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _465_ (.I(net32),
    .Z(gpio_pins[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _466_ (.I(net33),
    .Z(gpio_pins[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _467_ (.I(net3),
    .Z(gpio_pins[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _468_ (.I(net4),
    .Z(gpio_pins[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _469_ (.I(net5),
    .Z(gpio_pins[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _470_ (.I(net6),
    .Z(gpio_pins[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _471_ (.I(net7),
    .Z(gpio_pins[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _472_ (.I(net8),
    .Z(gpio_pins[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _473_ (.I(net9),
    .Z(gpio_pins[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _474_ (.I(net10),
    .Z(gpio_pins[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _475_ (.I(net11),
    .Z(gpio_pins[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _476_ (.I(net12),
    .Z(gpio_pins[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _477_ (.I(net14),
    .Z(gpio_pins[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _478_ (.I(net15),
    .Z(gpio_pins[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _479_ (.I(net16),
    .Z(gpio_pins[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _480_ (.I(net17),
    .Z(gpio_pins[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _481_ (.I(net18),
    .Z(gpio_pins[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _482_ (.I(net19),
    .Z(gpio_pins[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _483_ (.I(net20),
    .Z(gpio_pins[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _484_ (.I(net21),
    .Z(gpio_pins[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _485_ (.I(net22),
    .Z(gpio_pins[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _486_ (.I(net23),
    .Z(gpio_pins[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _487_ (.I(net25),
    .Z(gpio_pins[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _488_ (.I(net26),
    .Z(gpio_pins[31]));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[0]$_DFF_PN0_  (.D(\gpio_in_sync2[0] ),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\gpio_in_prev[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[10]$_DFF_PN0_  (.D(\gpio_in_sync2[10] ),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\gpio_in_prev[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[11]$_DFF_PN0_  (.D(\gpio_in_sync2[11] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\gpio_in_prev[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[12]$_DFF_PN0_  (.D(\gpio_in_sync2[12] ),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\gpio_in_prev[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[13]$_DFF_PN0_  (.D(\gpio_in_sync2[13] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_prev[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[14]$_DFF_PN0_  (.D(\gpio_in_sync2[14] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_prev[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[15]$_DFF_PN0_  (.D(\gpio_in_sync2[15] ),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\gpio_in_prev[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[16]$_DFF_PN0_  (.D(\gpio_in_sync2[16] ),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\gpio_in_prev[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[17]$_DFF_PN0_  (.D(\gpio_in_sync2[17] ),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\gpio_in_prev[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[18]$_DFF_PN0_  (.D(\gpio_in_sync2[18] ),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\gpio_in_prev[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[19]$_DFF_PN0_  (.D(\gpio_in_sync2[19] ),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\gpio_in_prev[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[1]$_DFF_PN0_  (.D(\gpio_in_sync2[1] ),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\gpio_in_prev[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[20]$_DFF_PN0_  (.D(\gpio_in_sync2[20] ),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\gpio_in_prev[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[21]$_DFF_PN0_  (.D(\gpio_in_sync2[21] ),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\gpio_in_prev[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[22]$_DFF_PN0_  (.D(\gpio_in_sync2[22] ),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\gpio_in_prev[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[23]$_DFF_PN0_  (.D(\gpio_in_sync2[23] ),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\gpio_in_prev[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[24]$_DFF_PN0_  (.D(\gpio_in_sync2[24] ),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\gpio_in_prev[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[25]$_DFF_PN0_  (.D(\gpio_in_sync2[25] ),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\gpio_in_prev[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[26]$_DFF_PN0_  (.D(\gpio_in_sync2[26] ),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\gpio_in_prev[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[27]$_DFF_PN0_  (.D(\gpio_in_sync2[27] ),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\gpio_in_prev[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[28]$_DFF_PN0_  (.D(\gpio_in_sync2[28] ),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\gpio_in_prev[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[29]$_DFF_PN0_  (.D(\gpio_in_sync2[29] ),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\gpio_in_prev[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[2]$_DFF_PN0_  (.D(\gpio_in_sync2[2] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\gpio_in_prev[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[30]$_DFF_PN0_  (.D(\gpio_in_sync2[30] ),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\gpio_in_prev[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[31]$_DFF_PN0_  (.D(\gpio_in_sync2[31] ),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\gpio_in_prev[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[3]$_DFF_PN0_  (.D(\gpio_in_sync2[3] ),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\gpio_in_prev[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[4]$_DFF_PN0_  (.D(\gpio_in_sync2[4] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_prev[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[5]$_DFF_PN0_  (.D(\gpio_in_sync2[5] ),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\gpio_in_prev[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[6]$_DFF_PN0_  (.D(\gpio_in_sync2[6] ),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\gpio_in_prev[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[7]$_DFF_PN0_  (.D(\gpio_in_sync2[7] ),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\gpio_in_prev[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[8]$_DFF_PN0_  (.D(\gpio_in_sync2[8] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\gpio_in_prev[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_prev[9]$_DFF_PN0_  (.D(\gpio_in_sync2[9] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\gpio_in_prev[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[0]$_DFF_PN0_  (.D(net2),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync1[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[10]$_DFF_PN0_  (.D(net3),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync1[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[11]$_DFF_PN0_  (.D(net4),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync1[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[12]$_DFF_PN0_  (.D(net5),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\gpio_in_sync1[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[13]$_DFF_PN0_  (.D(net6),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync1[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[14]$_DFF_PN0_  (.D(net7),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync1[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[15]$_DFF_PN0_  (.D(net8),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync1[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[16]$_DFF_PN0_  (.D(net9),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\gpio_in_sync1[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[17]$_DFF_PN0_  (.D(net10),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\gpio_in_sync1[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[18]$_DFF_PN0_  (.D(net11),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\gpio_in_sync1[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[19]$_DFF_PN0_  (.D(net12),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\gpio_in_sync1[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[1]$_DFF_PN0_  (.D(net13),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\gpio_in_sync1[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[20]$_DFF_PN0_  (.D(net14),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync1[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[21]$_DFF_PN0_  (.D(net15),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\gpio_in_sync1[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[22]$_DFF_PN0_  (.D(net16),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\gpio_in_sync1[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[23]$_DFF_PN0_  (.D(net17),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\gpio_in_sync1[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[24]$_DFF_PN0_  (.D(net18),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\gpio_in_sync1[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[25]$_DFF_PN0_  (.D(net19),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync1[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[26]$_DFF_PN0_  (.D(net20),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\gpio_in_sync1[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[27]$_DFF_PN0_  (.D(net21),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync1[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[28]$_DFF_PN0_  (.D(net22),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync1[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[29]$_DFF_PN0_  (.D(net23),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\gpio_in_sync1[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[2]$_DFF_PN0_  (.D(net24),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\gpio_in_sync1[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[30]$_DFF_PN0_  (.D(net25),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\gpio_in_sync1[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[31]$_DFF_PN0_  (.D(net26),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync1[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[3]$_DFF_PN0_  (.D(net27),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\gpio_in_sync1[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[4]$_DFF_PN0_  (.D(net28),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync1[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[5]$_DFF_PN0_  (.D(net29),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\gpio_in_sync1[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[6]$_DFF_PN0_  (.D(net30),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\gpio_in_sync1[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[7]$_DFF_PN0_  (.D(net31),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\gpio_in_sync1[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[8]$_DFF_PN0_  (.D(net32),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync1[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync1[9]$_DFF_PN0_  (.D(net33),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\gpio_in_sync1[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[0]$_DFF_PN0_  (.D(\gpio_in_sync1[0] ),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\gpio_in_sync2[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[10]$_DFF_PN0_  (.D(\gpio_in_sync1[10] ),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(\gpio_in_sync2[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[11]$_DFF_PN0_  (.D(\gpio_in_sync1[11] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync2[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[12]$_DFF_PN0_  (.D(\gpio_in_sync1[12] ),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(\gpio_in_sync2[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[13]$_DFF_PN0_  (.D(\gpio_in_sync1[13] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync2[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[14]$_DFF_PN0_  (.D(\gpio_in_sync1[14] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync2[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[15]$_DFF_PN0_  (.D(\gpio_in_sync1[15] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync2[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[16]$_DFF_PN0_  (.D(\gpio_in_sync1[16] ),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\gpio_in_sync2[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[17]$_DFF_PN0_  (.D(\gpio_in_sync1[17] ),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\gpio_in_sync2[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[18]$_DFF_PN0_  (.D(\gpio_in_sync1[18] ),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\gpio_in_sync2[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[19]$_DFF_PN0_  (.D(\gpio_in_sync1[19] ),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(\gpio_in_sync2[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[1]$_DFF_PN0_  (.D(\gpio_in_sync1[1] ),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\gpio_in_sync2[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[20]$_DFF_PN0_  (.D(\gpio_in_sync1[20] ),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync2[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[21]$_DFF_PN0_  (.D(\gpio_in_sync1[21] ),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(\gpio_in_sync2[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[22]$_DFF_PN0_  (.D(\gpio_in_sync1[22] ),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(\gpio_in_sync2[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[23]$_DFF_PN0_  (.D(\gpio_in_sync1[23] ),
    .RN(net1),
    .CLK(clknet_4_9_0_clk),
    .Q(\gpio_in_sync2[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[24]$_DFF_PN0_  (.D(\gpio_in_sync1[24] ),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\gpio_in_sync2[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[25]$_DFF_PN0_  (.D(\gpio_in_sync1[25] ),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync2[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[26]$_DFF_PN0_  (.D(\gpio_in_sync1[26] ),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync2[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[27]$_DFF_PN0_  (.D(\gpio_in_sync1[27] ),
    .RN(net1),
    .CLK(clknet_4_12_0_clk),
    .Q(\gpio_in_sync2[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[28]$_DFF_PN0_  (.D(\gpio_in_sync1[28] ),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync2[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[29]$_DFF_PN0_  (.D(\gpio_in_sync1[29] ),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(\gpio_in_sync2[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[2]$_DFF_PN0_  (.D(\gpio_in_sync1[2] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\gpio_in_sync2[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[30]$_DFF_PN0_  (.D(\gpio_in_sync1[30] ),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(\gpio_in_sync2[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[31]$_DFF_PN0_  (.D(\gpio_in_sync1[31] ),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(\gpio_in_sync2[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[3]$_DFF_PN0_  (.D(\gpio_in_sync1[3] ),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\gpio_in_sync2[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[4]$_DFF_PN0_  (.D(\gpio_in_sync1[4] ),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(\gpio_in_sync2[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[5]$_DFF_PN0_  (.D(\gpio_in_sync1[5] ),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(\gpio_in_sync2[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[6]$_DFF_PN0_  (.D(\gpio_in_sync1[6] ),
    .RN(net1),
    .CLK(clknet_4_3_0_clk),
    .Q(\gpio_in_sync2[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[7]$_DFF_PN0_  (.D(\gpio_in_sync1[7] ),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(\gpio_in_sync2[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[8]$_DFF_PN0_  (.D(\gpio_in_sync1[8] ),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(\gpio_in_sync2[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gpio_in_sync2[9]$_DFF_PN0_  (.D(\gpio_in_sync1[9] ),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(\gpio_in_sync2[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(net195));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[10]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net196));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[11]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net197));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[12]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net198));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[13]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(net199));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[14]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_4_0_0_clk),
    .Q(net200));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[15]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(net201));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[16]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(net202));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[17]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(net203));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[18]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(net204));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[19]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(net205));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[1]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(net206));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[20]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(net207));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[21]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_4_14_0_clk),
    .Q(net208));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[22]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(net209));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[23]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_4_11_0_clk),
    .Q(net210));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[24]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(net211));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[25]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(net212));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[26]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(net213));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[27]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_4_15_0_clk),
    .Q(net214));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[28]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(net215));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[29]$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_4_13_0_clk),
    .Q(net216));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[2]$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_4_6_0_clk),
    .Q(net217));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[30]$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_4_10_0_clk),
    .Q(net218));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[31]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_4_8_0_clk),
    .Q(net219));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[3]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_4_4_0_clk),
    .Q(net220));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[4]$_DFFE_PN0P_  (.D(_026_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(net221));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[5]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(net222));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[6]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_4_2_0_clk),
    .Q(net223));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[7]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_4_1_0_clk),
    .Q(net224));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[8]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_4_5_0_clk),
    .Q(net225));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \int_status_reg[9]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_4_7_0_clk),
    .Q(net226));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 hold1 (.I(net227),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_91 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_92 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_93 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_94 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_95 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_96 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_97 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_98 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_99 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_139 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(gpio_out[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(gpio_out[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(gpio_out[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(gpio_out[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(gpio_out[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(gpio_out[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(gpio_out[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(gpio_out[16]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(gpio_out[17]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(gpio_out[18]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(gpio_out[19]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(gpio_out[1]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(gpio_out[20]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(gpio_out[21]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(gpio_out[22]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(gpio_out[23]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(gpio_out[24]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(gpio_out[25]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(gpio_out[26]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(gpio_out[27]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(gpio_out[28]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(gpio_out[29]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(gpio_out[2]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(gpio_out[30]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(gpio_out[31]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(gpio_out[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(gpio_out[4]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(gpio_out[5]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(gpio_out[6]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(gpio_out[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(gpio_out[8]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(gpio_out[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input33 (.I(int_clear[0]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(int_clear[10]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(int_clear[11]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(int_clear[12]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(int_clear[13]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(int_clear[14]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input39 (.I(int_clear[15]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input40 (.I(int_clear[16]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(int_clear[17]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(int_clear[18]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(int_clear[19]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input44 (.I(int_clear[1]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(int_clear[20]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input46 (.I(int_clear[21]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input47 (.I(int_clear[22]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(int_clear[23]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(int_clear[24]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input50 (.I(int_clear[25]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input51 (.I(int_clear[26]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(int_clear[27]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(int_clear[28]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input54 (.I(int_clear[29]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input55 (.I(int_clear[2]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input56 (.I(int_clear[30]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input57 (.I(int_clear[31]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input58 (.I(int_clear[3]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input59 (.I(int_clear[4]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input60 (.I(int_clear[5]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input61 (.I(int_clear[6]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input62 (.I(int_clear[7]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input63 (.I(int_clear[8]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input64 (.I(int_clear[9]),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input65 (.I(int_enable[0]),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input66 (.I(int_enable[10]),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input67 (.I(int_enable[11]),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input68 (.I(int_enable[12]),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input69 (.I(int_enable[13]),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input70 (.I(int_enable[14]),
    .Z(net71));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input71 (.I(int_enable[15]),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input72 (.I(int_enable[16]),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input73 (.I(int_enable[17]),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input74 (.I(int_enable[18]),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input75 (.I(int_enable[19]),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input76 (.I(int_enable[1]),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input77 (.I(int_enable[20]),
    .Z(net78));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input78 (.I(int_enable[21]),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input79 (.I(int_enable[22]),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input80 (.I(int_enable[23]),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input81 (.I(int_enable[24]),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input82 (.I(int_enable[25]),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input83 (.I(int_enable[26]),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input84 (.I(int_enable[27]),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input85 (.I(int_enable[28]),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input86 (.I(int_enable[29]),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input87 (.I(int_enable[2]),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input88 (.I(int_enable[30]),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input89 (.I(int_enable[31]),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input90 (.I(int_enable[3]),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input91 (.I(int_enable[4]),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input92 (.I(int_enable[5]),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input93 (.I(int_enable[6]),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input94 (.I(int_enable[7]),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input95 (.I(int_enable[8]),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input96 (.I(int_enable[9]),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input97 (.I(int_polarity[0]),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input98 (.I(int_polarity[10]),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input99 (.I(int_polarity[11]),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input100 (.I(int_polarity[12]),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input101 (.I(int_polarity[13]),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input102 (.I(int_polarity[14]),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input103 (.I(int_polarity[15]),
    .Z(net104));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input104 (.I(int_polarity[16]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input105 (.I(int_polarity[17]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input106 (.I(int_polarity[18]),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input107 (.I(int_polarity[19]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input108 (.I(int_polarity[1]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input109 (.I(int_polarity[20]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input110 (.I(int_polarity[21]),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input111 (.I(int_polarity[22]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input112 (.I(int_polarity[23]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input113 (.I(int_polarity[24]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input114 (.I(int_polarity[25]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input115 (.I(int_polarity[26]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input116 (.I(int_polarity[27]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input117 (.I(int_polarity[28]),
    .Z(net118));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input118 (.I(int_polarity[29]),
    .Z(net119));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input119 (.I(int_polarity[2]),
    .Z(net120));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input120 (.I(int_polarity[30]),
    .Z(net121));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input121 (.I(int_polarity[31]),
    .Z(net122));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input122 (.I(int_polarity[3]),
    .Z(net123));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input123 (.I(int_polarity[4]),
    .Z(net124));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input124 (.I(int_polarity[5]),
    .Z(net125));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input125 (.I(int_polarity[6]),
    .Z(net126));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input126 (.I(int_polarity[7]),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input127 (.I(int_polarity[8]),
    .Z(net128));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input128 (.I(int_polarity[9]),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input129 (.I(int_type[0]),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input130 (.I(int_type[10]),
    .Z(net131));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input131 (.I(int_type[11]),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input132 (.I(int_type[12]),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input133 (.I(int_type[13]),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input134 (.I(int_type[14]),
    .Z(net135));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input135 (.I(int_type[15]),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input136 (.I(int_type[16]),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input137 (.I(int_type[17]),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input138 (.I(int_type[18]),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input139 (.I(int_type[19]),
    .Z(net140));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input140 (.I(int_type[1]),
    .Z(net141));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input141 (.I(int_type[20]),
    .Z(net142));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input142 (.I(int_type[21]),
    .Z(net143));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input143 (.I(int_type[22]),
    .Z(net144));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input144 (.I(int_type[23]),
    .Z(net145));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input145 (.I(int_type[24]),
    .Z(net146));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input146 (.I(int_type[25]),
    .Z(net147));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input147 (.I(int_type[26]),
    .Z(net148));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input148 (.I(int_type[27]),
    .Z(net149));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input149 (.I(int_type[28]),
    .Z(net150));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input150 (.I(int_type[29]),
    .Z(net151));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input151 (.I(int_type[2]),
    .Z(net152));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input152 (.I(int_type[30]),
    .Z(net153));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input153 (.I(int_type[31]),
    .Z(net154));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input154 (.I(int_type[3]),
    .Z(net155));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input155 (.I(int_type[4]),
    .Z(net156));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input156 (.I(int_type[5]),
    .Z(net157));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input157 (.I(int_type[6]),
    .Z(net158));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input158 (.I(int_type[7]),
    .Z(net159));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input159 (.I(int_type[8]),
    .Z(net160));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input160 (.I(int_type[9]),
    .Z(net161));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output161 (.I(net162),
    .Z(gpio_in[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output162 (.I(net163),
    .Z(gpio_in[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output163 (.I(net164),
    .Z(gpio_in[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output164 (.I(net165),
    .Z(gpio_in[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output165 (.I(net166),
    .Z(gpio_in[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output166 (.I(net167),
    .Z(gpio_in[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output167 (.I(net168),
    .Z(gpio_in[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output168 (.I(net169),
    .Z(gpio_in[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output169 (.I(net170),
    .Z(gpio_in[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output170 (.I(net171),
    .Z(gpio_in[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output171 (.I(net172),
    .Z(gpio_in[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output172 (.I(net173),
    .Z(gpio_in[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output173 (.I(net174),
    .Z(gpio_in[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output174 (.I(net175),
    .Z(gpio_in[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output175 (.I(net176),
    .Z(gpio_in[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output176 (.I(net177),
    .Z(gpio_in[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output177 (.I(net178),
    .Z(gpio_in[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output178 (.I(net179),
    .Z(gpio_in[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output179 (.I(net180),
    .Z(gpio_in[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output180 (.I(net181),
    .Z(gpio_in[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output181 (.I(net182),
    .Z(gpio_in[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output182 (.I(net183),
    .Z(gpio_in[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output183 (.I(net184),
    .Z(gpio_in[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output184 (.I(net185),
    .Z(gpio_in[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output185 (.I(net186),
    .Z(gpio_in[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output186 (.I(net187),
    .Z(gpio_in[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output187 (.I(net188),
    .Z(gpio_in[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output188 (.I(net189),
    .Z(gpio_in[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output189 (.I(net190),
    .Z(gpio_in[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output190 (.I(net191),
    .Z(gpio_in[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output191 (.I(net192),
    .Z(gpio_in[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output192 (.I(net193),
    .Z(gpio_in[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output193 (.I(net194),
    .Z(int_out));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output194 (.I(net195),
    .Z(int_status[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output195 (.I(net196),
    .Z(int_status[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output196 (.I(net197),
    .Z(int_status[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output197 (.I(net198),
    .Z(int_status[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output198 (.I(net199),
    .Z(int_status[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output199 (.I(net200),
    .Z(int_status[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output200 (.I(net201),
    .Z(int_status[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output201 (.I(net202),
    .Z(int_status[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output202 (.I(net203),
    .Z(int_status[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output203 (.I(net204),
    .Z(int_status[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output204 (.I(net205),
    .Z(int_status[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output205 (.I(net206),
    .Z(int_status[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output206 (.I(net207),
    .Z(int_status[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output207 (.I(net208),
    .Z(int_status[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output208 (.I(net209),
    .Z(int_status[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output209 (.I(net210),
    .Z(int_status[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output210 (.I(net211),
    .Z(int_status[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output211 (.I(net212),
    .Z(int_status[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output212 (.I(net213),
    .Z(int_status[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output213 (.I(net214),
    .Z(int_status[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output214 (.I(net215),
    .Z(int_status[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output215 (.I(net216),
    .Z(int_status[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output216 (.I(net217),
    .Z(int_status[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output217 (.I(net218),
    .Z(int_status[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output218 (.I(net219),
    .Z(int_status[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output219 (.I(net220),
    .Z(int_status[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output220 (.I(net221),
    .Z(int_status[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output221 (.I(net222),
    .Z(int_status[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output222 (.I(net223),
    .Z(int_status[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output223 (.I(net224),
    .Z(int_status[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output224 (.I(net225),
    .Z(int_status[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output225 (.I(net226),
    .Z(int_status[9]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_8_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_9_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_10_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_11_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_12_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_13_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_14_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_4_15_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload0 (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload1 (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload2 (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload3 (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload4 (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload5 (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload6 (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload7 (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload8 (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload9 (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload10 (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload11 (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload12 (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload13 (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload14 (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net227));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_11 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_422 ();
endmodule
