
* cell parameterized_freq_divider
* pin duty_cycle[2]
* pin divide_value[12]
* pin divide_value[11]
* pin divide_value[10]
* pin divide_value[9]
* pin duty_cycle[3]
* pin divide_value[2]
* pin divide_value[3]
* pin divide_value[5]
* pin divide_value[7]
* pin duty_cycle[1]
* pin divide_value[6]
* pin divide_value[4]
* pin divide_value[8]
* pin divide_value[0]
* pin divide_value[13]
* pin duty_cycle[0]
* pin divide_value[1]
* pin enable
* pin clk_in
* pin rst_n
* pin PWELL
* pin NWELL
* pin divide_value[14]
* pin duty_cycle[4]
* pin duty_cycle[5]
* pin divide_value[15]
* pin duty_cycle[6]
* pin clk_out
.SUBCKT parameterized_freq_divider 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
+ 19 20 21 25 44 2885 2886 2887 2888 2889 2890
* net 1 duty_cycle[2]
* net 2 divide_value[12]
* net 3 divide_value[11]
* net 4 divide_value[10]
* net 5 divide_value[9]
* net 6 duty_cycle[3]
* net 7 divide_value[2]
* net 8 divide_value[3]
* net 9 divide_value[5]
* net 10 divide_value[7]
* net 11 duty_cycle[1]
* net 12 divide_value[6]
* net 13 divide_value[4]
* net 14 divide_value[8]
* net 15 divide_value[0]
* net 16 divide_value[13]
* net 17 duty_cycle[0]
* net 18 divide_value[1]
* net 19 enable
* net 20 clk_in
* net 21 rst_n
* net 25 PWELL
* net 44 NWELL
* net 2885 divide_value[14]
* net 2886 duty_cycle[4]
* net 2887 duty_cycle[5]
* net 2888 divide_value[15]
* net 2889 duty_cycle[6]
* net 2890 clk_out
* cell instance $2 r0 *1 356.06,1.4
X$2 1 25 44 22 BUF_X2
* cell instance $8 r0 *1 358.34,1.4
X$8 2 25 44 34 BUF_X2
* cell instance $14 r0 *1 361.57,1.4
X$14 3 25 44 26 CLKBUF_X3
* cell instance $20 r0 *1 367.84,1.4
X$20 4 25 44 32 CLKBUF_X3
* cell instance $26 r0 *1 370.12,1.4
X$26 5 25 44 23 CLKBUF_X3
* cell instance $32 r0 *1 377.34,1.4
X$32 6 25 44 38 BUF_X2
* cell instance $38 m0 *1 400.33,4.2
X$38 7 25 44 186 CLKBUF_X3
* cell instance $44 r0 *1 400.9,1.4
X$44 8 25 44 24 CLKBUF_X3
* cell instance $50 m0 *1 401.47,4.2
X$50 9 25 44 48 CLKBUF_X3
* cell instance $57 r0 *1 399.57,1.4
X$57 10 44 39 25 BUF_X4
* cell instance $63 r0 *1 398.81,1.4
X$63 11 25 44 42 BUF_X2
* cell instance $68 r0 *1 402.8,1.4
X$68 12 25 44 40 CLKBUF_X3
* cell instance $74 r0 *1 403.94,1.4
X$74 13 25 44 90 BUF_X1
* cell instance $80 r0 *1 404.7,1.4
X$80 14 25 44 49 BUF_X1
* cell instance $86 r0 *1 408.31,1.4
X$86 15 25 44 201 BUF_X2
* cell instance $93 r0 *1 405.27,1.4
X$93 16 25 44 31 BUF_X1
* cell instance $99 r0 *1 406.22,1.4
X$99 17 25 44 27 CLKBUF_X3
* cell instance $105 r0 *1 409.07,1.4
X$105 18 25 44 28 BUF_X2
* cell instance $110 r0 *1 413.82,1.4
X$110 19 25 44 29 BUF_X1
* cell instance $120 r0 *1 421.23,1.4
X$120 20 44 30 25 BUF_X4
* cell instance $122 r0 *1 423.51,1.4
X$122 25 43 44 21 BUF_X8
* cell instance $135 m0 *1 383.99,12.6
X$135 22 24 44 25 222 AND2_X1
* cell instance $137 m0 *1 383.61,4.2
X$137 22 25 44 35 BUF_X2
* cell instance $141 r0 *1 336.49,9.8
X$141 22 60 44 25 183 AND2_X1
* cell instance $145 r0 *1 392.16,21
X$145 22 301 44 25 535 AND2_X1
* cell instance $148 m0 *1 334.4,21
X$148 22 189 44 25 381 AND2_X1
* cell instance $150 r0 *1 334.78,15.4
X$150 22 158 44 25 293 AND2_X1
* cell instance $153 r0 *1 386.65,21
X$153 467 38 22 25 44 443 OR3_X1
* cell instance $155 r0 *1 389.5,21
X$155 22 186 44 25 442 AND2_X1
* cell instance $178 m0 *1 351.69,4.2
X$178 36 23 44 25 99 AND2_X1
* cell instance $180 m0 *1 388.36,4.2
X$180 49 23 25 44 50 NOR2_X1
* cell instance $182 m0 *1 387.98,12.6
X$182 23 254 44 25 250 XNOR2_X1
* cell instance $184 m0 *1 385.7,7
X$184 32 23 41 176 25 44 151 OR4_X1
* cell instance $187 r0 *1 348.65,9.8
X$187 23 123 25 44 199 NAND2_X1
* cell instance $189 m0 *1 348.46,21
X$189 323 23 44 25 407 AND2_X1
* cell instance $192 r0 *1 364.8,7
X$192 33 23 44 25 178 AND2_X1
* cell instance $194 m0 *1 352.45,15.4
X$194 167 23 44 25 214 AND2_X1
* cell instance $196 m0 *1 369.93,21
X$196 213 23 44 25 368 AND2_X1
* cell instance $199 m0 *1 364.99,4.2
X$199 35 23 44 25 64 AND2_X1
* cell instance $217 m0 *1 401.47,26.6
X$217 24 534 44 25 500 XNOR2_X1
* cell instance $220 m0 *1 392.16,26.6
X$220 24 213 25 44 618 NAND2_X1
* cell instance $223 r0 *1 381.33,4.2
X$223 38 24 44 25 121 AND2_X1
* cell instance $225 m0 *1 398.62,18.2
X$225 24 186 25 44 265 OR2_X1
* cell instance $227 m0 *1 375.25,26.6
X$227 513 24 44 25 533 AND2_X1
* cell instance $230 r0 *1 378.67,9.8
X$230 167 24 44 25 182 AND2_X1
* cell instance $233 m0 *1 374.49,9.8
X$233 123 24 44 25 180 AND2_X1
* cell instance $235 r0 *1 388.55,21
X$235 42 24 44 25 466 AND2_X1
* cell instance $236 m0 *1 381.52,107.8
X$236 2791 2347 2346 44 2810 25 NOR3_X2
* cell instance $238 m0 *1 382.85,107.8
X$238 2346 2347 2791 25 44 2808 OR3_X2
* cell instance $241 m0 *1 387.79,107.8
X$241 2751 2776 25 44 2562 OR2_X1
* cell instance $244 m0 *1 390.83,107.8
X$244 2562 2593 25 44 2812 NAND2_X1
* cell instance $246 m0 *1 391.59,107.8
X$246 2751 2593 25 44 2813 OR2_X1
* cell instance $249 r0 *1 381.33,107.8
X$249 764 2294 2808 44 2806 25 OAI21_X1
* cell instance $251 r0 *1 382.47,107.8
X$251 25 2593 2810 1884 2811 44 AOI21_X4
* cell instance $254 r0 *1 385.51,107.8
X$254 25 2808 2776 764 2793 2294 44 OAI211_X4
* cell instance $258 r0 *1 391.21,107.8
X$258 2812 2813 2792 44 25 2779 OAI21_X2
* cell instance $259 r0 *1 392.54,107.8
X$259 2793 44 2307 25 BUF_X4
* cell instance $260 m0 *1 395.2,107.8
X$260 25 2814 2815 2582 2752 2785 44 AOI22_X4
* cell instance $261 m0 *1 393.49,107.8
X$261 2422 2015 2307 2592 25 2785 44 NAND4_X2
* cell instance $264 m0 *1 399.38,107.8
X$264 757 2331 25 44 2773 NAND2_X2
* cell instance $270 r0 *1 395.2,107.8
X$270 2685 2369 2423 44 25 2815 OAI21_X2
* cell instance $271 r0 *1 396.53,107.8
X$271 2793 25 44 2348 INV_X4
* cell instance $274 r0 *1 398.05,107.8
X$274 2348 2331 2754 25 44 NOR2_X4
* cell instance $275 r0 *1 399.76,107.8
X$275 2754 2832 25 44 2753 NAND2_X1
* cell instance $277 r0 *1 400.71,107.8
X$277 2307 2685 25 44 2816 NAND2_X2
* cell instance $278 m0 *1 402.04,107.8
X$278 25 2794 2816 2773 2771 2689 44 OAI22_X4
* cell instance $279 m0 *1 401.47,107.8
X$279 2816 2755 25 44 2729 NOR2_X1
* cell instance $280 m0 *1 405.27,107.8
X$280 2794 2685 25 44 2795 NOR2_X1
* cell instance $282 r0 *1 401.66,107.8
X$282 2422 2755 25 44 2794 XNOR2_X2
* cell instance $283 r0 *1 403.56,107.8
X$283 2773 2689 25 44 2821 NOR2_X2
* cell instance $284 r0 *1 404.51,107.8
X$284 25 2796 2795 2756 2850 2685 44 AOI22_X4
* cell instance $286 m0 *1 406.22,107.8
X$286 2779 2797 25 2486 44 NAND2_X4
* cell instance $287 m0 *1 408.12,107.8
X$287 2797 2779 44 25 2780 AND2_X1
* cell instance $289 m0 *1 409.07,107.8
X$289 2809 2779 25 44 2629 OR2_X1
* cell instance $293 m0 *1 412.3,107.8
X$293 2780 44 2018 25 BUF_X4
* cell instance $296 m0 *1 415.34,107.8
X$296 2758 2757 1951 2771 1364 2019 25 44 OAI221_X2
* cell instance $301 r0 *1 408.31,107.8
X$301 2527 2529 2809 2836 25 2628 44 NAND4_X2
* cell instance $302 r0 *1 410.02,107.8
X$302 2413 2654 25 44 2828 NOR2_X1
* cell instance $305 m0 *1 419.52,107.8
X$305 2761 2000 2021 25 44 2759 NOR3_X1
* cell instance $308 m0 *1 420.47,107.8
X$308 25 2762 2000 2021 1999 44 AOI21_X4
* cell instance $310 m0 *1 423.13,107.8
X$310 2047 2073 25 44 2801 NOR2_X1
* cell instance $312 m0 *1 423.89,107.8
X$312 2782 2801 2734 44 25 2800 OAI21_X2
* cell instance $316 r0 *1 420.85,107.8
X$316 639 2796 2807 44 2799 25 OAI21_X1
* cell instance $317 r0 *1 421.61,107.8
X$317 639 2796 2807 25 44 2798 OR3_X1
* cell instance $318 r0 *1 422.56,107.8
X$318 2798 2799 1364 25 44 2734 NAND3_X2
* cell instance $321 r0 *1 424.46,107.8
X$321 2799 2798 44 25 2563 AND2_X2
* cell instance $324 m0 *1 425.6,107.8
X$324 2800 2019 2763 44 25 2567 OAI21_X4
* cell instance $491 m0 *1 391.02,105
X$491 1625 2591 2623 44 25 2676 OAI21_X2
* cell instance $497 r0 *1 391.02,105
X$497 757 2751 25 44 2777 NOR2_X1
* cell instance $498 r0 *1 391.59,105
X$498 2777 2593 2792 44 25 2228 OAI21_X4
* cell instance $501 r0 *1 395.2,105
X$501 2307 2692 2676 44 25 2814 AND3_X1
* cell instance $503 r0 *1 396.53,105
X$503 2692 2331 2307 25 2752 44 AOI21_X2
* cell instance $505 m0 *1 397.29,105
X$505 2676 2692 1885 25 44 2650 NAND3_X2
* cell instance $511 m0 *1 399.19,105
X$511 2773 2753 2688 2689 2599 2693 44 25 AOI221_X2
* cell instance $515 m0 *1 403.56,105
X$515 2691 2690 1885 44 2748 25 NOR3_X2
* cell instance $516 m0 *1 404.89,105
X$516 2691 2690 25 44 2730 NOR2_X1
* cell instance $517 m0 *1 405.46,105
X$517 2730 2756 1885 44 25 2732 MUX2_X2
* cell instance $520 m0 *1 409.45,105
X$520 25 2757 2486 2086 1952 44 AOI21_X4
* cell instance $523 m0 *1 413.63,105
X$523 2134 2731 2379 2732 2733 2772 44 25 AOI221_X2
* cell instance $524 m0 *1 415.72,105
X$524 25 2732 2733 2153 2731 2134 44 AOI22_X4
* cell instance $527 r0 *1 399,105
X$527 25 2692 2754 2689 2755 2656 44 NAND4_X4
* cell instance $528 r0 *1 402.42,105
X$528 2755 2422 25 44 2778 NOR2_X1
* cell instance $529 r0 *1 402.99,105
X$529 2778 2273 2652 44 25 2784 OAI21_X2
* cell instance $530 r0 *1 404.32,105
X$530 2652 2273 25 44 2796 NOR2_X2
* cell instance $531 r0 *1 405.27,105
X$531 25 2758 2748 1885 2756 44 AOI21_X4
* cell instance $535 r0 *1 411.73,105
X$535 2653 2529 2780 44 2698 25 NOR3_X2
* cell instance $537 r0 *1 413.44,105
X$537 2018 2413 2068 44 25 2733 OAI21_X2
* cell instance $539 r0 *1 414.96,105
X$539 25 2758 2757 2771 2074 1951 44 OAI22_X4
* cell instance $541 r0 *1 418.38,105
X$541 2772 44 2000 25 BUF_X4
* cell instance $543 r0 *1 419.9,105
X$543 2759 2760 25 44 2770 NOR2_X1
* cell instance $545 m0 *1 420.09,105
X$545 2770 2532 25 44 2735 NOR2_X1
* cell instance $546 m0 *1 423.7,105
X$546 2074 2428 2762 44 2747 25 OAI21_X1
* cell instance $547 m0 *1 424.46,105
X$547 2747 2761 44 2736 25 XOR2_X2
* cell instance $550 r0 *1 420.47,105
X$550 2021 2699 25 44 2781 NOR2_X1
* cell instance $552 r0 *1 421.23,105
X$552 2760 2759 2781 25 44 2701 OR3_X1
* cell instance $553 r0 *1 422.18,105
X$553 25 2782 2762 2761 2734 2745 44 NAND4_X4
* cell instance $554 r0 *1 425.6,105
X$554 2761 2762 2763 25 44 2764 OR3_X2
* cell instance $556 m0 *1 430.16,105
X$556 2745 2764 44 25 2661 AND2_X2
* cell instance $557 m0 *1 428.07,105
X$557 1948 1949 2043 2764 2745 2710 44 25 AOI221_X2
* cell instance $563 r0 *1 429.21,105
X$563 2764 2745 25 2658 44 NAND2_X4
* cell instance $567 r0 *1 435.1,105
X$567 2704 2658 2735 25 44 2766 OR3_X1
* cell instance $568 m0 *1 435.86,105
X$568 2704 44 2539 25 BUF_X4
* cell instance $569 m0 *1 435.29,105
X$569 2043 2658 25 44 2703 NAND2_X1
* cell instance $572 m0 *1 438.14,105
X$572 25 2539 2740 2661 2538 2606 44 OAI211_X4
* cell instance $574 m0 *1 442.89,105
X$574 2631 2567 2737 44 25 2765 AND3_X1
* cell instance $575 m0 *1 443.84,105
X$575 2736 2539 25 44 2737 NOR2_X1
* cell instance $576 m0 *1 444.41,105
X$576 2567 2631 25 44 2738 NAND2_X1
* cell instance $579 r0 *1 436.43,105
X$579 2735 2704 2658 44 25 1562 OAI21_X2
* cell instance $580 r0 *1 437.76,105
X$580 2766 1562 25 44 2239 NAND2_X2
* cell instance $585 r0 *1 444.41,105
X$585 2239 2765 2736 2738 2202 44 25 AOI211_X2
* cell instance $587 m0 *1 445.36,105
X$587 2737 2738 2736 25 44 2319 MUX2_X1
* cell instance $746 m0 *1 419.33,40.6
X$746 921 922 923 25 44 935 NOR3_X1
* cell instance $747 m0 *1 418.76,40.6
X$747 881 940 25 44 880 NOR2_X1
* cell instance $749 m0 *1 420.28,40.6
X$749 935 923 921 25 917 44 AOI21_X2
* cell instance $750 m0 *1 421.61,40.6
X$750 924 919 917 25 848 44 AOI21_X1
* cell instance $751 m0 *1 422.37,40.6
X$751 969 924 917 930 44 25 814 AND4_X1
* cell instance $752 m0 *1 423.51,40.6
X$752 927 882 44 25 926 XNOR2_X1
* cell instance $753 m0 *1 424.65,40.6
X$753 992 25 44 927 INV_X1
* cell instance $754 m0 *1 425.03,40.6
X$754 927 880 25 44 884 NOR2_X1
* cell instance $755 m0 *1 425.6,40.6
X$755 883 884 929 25 44 930 MUX2_X1
* cell instance $812 m0 *1 388.93,40.6
X$812 781 874 948 44 25 949 HA_X1
* cell instance $815 m0 *1 393.3,40.6
X$815 950 887 1257 44 25 913 HA_X1
* cell instance $819 m0 *1 407.55,40.6
X$819 944 879 916 25 44 841 NAND3_X1
* cell instance $820 m0 *1 408.31,40.6
X$820 879 916 842 25 44 813 NAND3_X1
* cell instance $822 m0 *1 409.26,40.6
X$822 944 879 916 842 25 44 943 NAND4_X1
* cell instance $825 m0 *1 411.16,40.6
X$825 924 917 943 44 25 844 AND3_X1
* cell instance $826 m0 *1 412.11,40.6
X$826 917 25 44 817 INV_X1
* cell instance $831 r0 *1 389.12,40.6
X$831 948 913 949 863 25 44 789 AOI211_X4
* cell instance $835 r0 *1 401.85,40.6
X$835 915 971 44 25 945 XNOR2_X1
* cell instance $838 r0 *1 403.94,40.6
X$838 967 878 915 25 44 983 OR3_X1
* cell instance $839 r0 *1 404.89,40.6
X$839 878 44 981 25 BUF_X4
* cell instance $841 r0 *1 406.6,40.6
X$841 944 947 945 25 812 44 AOI21_X2
* cell instance $844 r0 *1 414.2,40.6
X$844 968 918 25 44 842 OR2_X1
* cell instance $845 r0 *1 414.96,40.6
X$845 918 968 25 44 919 NOR2_X1
* cell instance $846 m0 *1 417.62,40.6
X$846 940 939 25 44 921 OR2_X1
* cell instance $847 m0 *1 415.15,40.6
X$847 922 940 881 44 25 878 OAI21_X4
* cell instance $851 r0 *1 416.48,40.6
X$851 920 967 25 44 939 NOR2_X1
* cell instance $855 r0 *1 418.38,40.6
X$855 939 989 25 44 881 OR2_X1
* cell instance $859 r0 *1 423.13,40.6
X$859 925 880 926 25 44 924 MUX2_X1
* cell instance $862 r0 *1 426.17,40.6
X$862 928 883 25 44 929 NAND2_X1
* cell instance $976 m0 *1 332.31,23.8
X$976 431 25 44 430 INV_X1
* cell instance $981 m0 *1 335.16,23.8
X$981 432 25 44 486 INV_X1
* cell instance $984 m0 *1 337.82,23.8
X$984 467 34 44 25 433 AND2_X1
* cell instance $987 m0 *1 346.18,23.8
X$987 434 25 44 435 INV_X1
* cell instance $992 r0 *1 332.31,23.8
X$992 467 60 44 25 504 AND2_X1
* cell instance $997 r0 *1 338.2,23.8
X$997 25 485 523 525 487 486 44 FA_X1
* cell instance $1000 r0 *1 341.43,23.8
X$1000 26 323 25 44 524 NAND2_X1
* cell instance $1002 r0 *1 343.52,23.8
X$1002 468 25 44 506 INV_X1
* cell instance $1005 r0 *1 345.8,23.8
X$1005 435 469 526 44 25 541 HA_X1
* cell instance $1007 m0 *1 350.93,23.8
X$1007 450 408 470 44 25 436 HA_X1
* cell instance $1012 m0 *1 356.82,23.8
X$1012 452 25 44 489 INV_X1
* cell instance $1013 m0 *1 357.2,23.8
X$1013 25 392 490 530 454 437 44 FA_X1
* cell instance $1016 m0 *1 363.47,23.8
X$1016 48 323 25 44 492 NAND2_X1
* cell instance $1023 r0 *1 352.26,23.8
X$1023 470 44 528 25 BUF_X4
* cell instance $1025 r0 *1 356.63,23.8
X$1025 489 490 564 44 25 510 HA_X1
* cell instance $1033 r0 *1 362.52,23.8
X$1033 25 493 471 512 492 472 44 FA_X1
* cell instance $1036 r0 *1 368.79,23.8
X$1036 494 25 44 544 INV_X1
* cell instance $1040 r0 *1 373.35,23.8
X$1040 473 25 44 532 INV_X1
* cell instance $1041 r0 *1 373.73,23.8
X$1041 25 474 568 514 459 220 44 FA_X1
* cell instance $1042 m0 *1 376.01,23.8
X$1042 186 323 25 44 459 NAND2_X1
* cell instance $1047 m0 *1 380.57,23.8
X$1047 25 440 438 463 462 439 44 FA_X1
* cell instance $1048 m0 *1 383.61,23.8
X$1048 25 464 496 441 463 318 44 FA_X1
* cell instance $1050 m0 *1 387.41,23.8
X$1050 25 442 464 515 466 465 44 FA_X1
* cell instance $1059 r0 *1 379.62,23.8
X$1059 25 496 475 476 438 411 44 FA_X1
* cell instance $1060 r0 *1 382.66,23.8
X$1060 467 291 44 25 440 AND2_X1
* cell instance $1064 r0 *1 392.92,23.8
X$1064 42 291 44 25 516 AND2_X1
* cell instance $1068 m0 *1 399.19,23.8
X$1068 47 415 44 25 458 XNOR2_X1
* cell instance $1071 r0 *1 400.71,23.8
X$1071 501 25 44 499 INV_X1
* cell instance $1072 m0 *1 400.9,23.8
X$1072 457 456 416 44 413 25 OAI21_X1
* cell instance $1076 m0 *1 404.89,23.8
X$1076 424 444 451 44 455 25 OAI21_X1
* cell instance $1081 r0 *1 401.09,23.8
X$1081 480 458 501 44 25 457 HA_X1
* cell instance $1082 r0 *1 402.99,23.8
X$1082 499 455 498 25 456 44 AOI21_X1
* cell instance $1083 r0 *1 403.75,23.8
X$1083 478 500 451 44 25 497 HA_X1
* cell instance $1084 r0 *1 405.65,23.8
X$1084 497 25 44 498 INV_X1
* cell instance $1088 r0 *1 410.97,23.8
X$1088 196 57 160 159 25 44 477 NOR4_X1
* cell instance $1090 m0 *1 411.35,23.8
X$1090 229 168 132 54 25 44 495 NOR4_X1
* cell instance $1093 m0 *1 417.05,23.8
X$1093 335 376 44 25 303 AND2_X1
* cell instance $1095 m0 *1 420.85,23.8
X$1095 396 445 44 25 302 AND2_X1
* cell instance $1096 m0 *1 421.61,23.8
X$1096 445 336 25 44 447 NAND2_X1
* cell instance $1100 m0 *1 426.93,23.8
X$1100 446 447 44 25 448 XNOR2_X1
* cell instance $1112 r0 *1 411.92,23.8
X$1112 495 477 491 488 25 44 419 NAND4_X1
* cell instance $1114 r0 *1 415.91,23.8
X$1114 478 25 44 479 BUF_X1
* cell instance $1115 r0 *1 416.48,23.8
X$1115 376 481 479 480 25 44 491 NOR4_X1
* cell instance $1119 r0 *1 419.52,23.8
X$1119 397 25 44 481 BUF_X1
* cell instance $1122 r0 *1 420.66,23.8
X$1122 418 480 479 481 44 25 445 AND4_X1
* cell instance $1124 r0 *1 421.99,23.8
X$1124 336 481 479 25 44 484 NAND3_X1
* cell instance $1126 r0 *1 422.94,23.8
X$1126 482 484 44 25 517 XNOR2_X1
* cell instance $1127 r0 *1 424.08,23.8
X$1127 25 30 483 43 446 396 44 DFFR_X2
* cell instance $1129 r0 *1 428.45,23.8
X$1129 448 195 25 44 483 NOR2_X1
* cell instance $2007 m0 *1 359.67,99.4
X$2007 2553 2573 25 44 2621 NOR2_X1
* cell instance $2010 m0 *1 360.43,99.4
X$2010 2573 2553 25 44 2487 OR2_X1
* cell instance $2013 m0 *1 362.9,99.4
X$2013 2680 2414 2584 44 25 2576 AND3_X1
* cell instance $2017 r0 *1 359.67,99.4
X$2017 2621 2462 44 25 2640 AND2_X1
* cell instance $2022 r0 *1 361.95,99.4
X$2022 2458 25 44 2641 BUF_X2
* cell instance $2023 r0 *1 362.71,99.4
X$2023 2621 2414 25 44 2668 XNOR2_X2
* cell instance $2025 r0 *1 364.99,99.4
X$2025 2641 2487 1842 25 44 2705 NAND3_X1
* cell instance $2028 r0 *1 366.89,99.4
X$2028 2517 1581 25 44 2642 NAND2_X1
* cell instance $2029 m0 *1 367.46,99.4
X$2029 1512 2401 2146 25 2622 44 AOI21_X2
* cell instance $2032 r0 *1 367.46,99.4
X$2032 2517 763 25 44 2643 NAND2_X1
* cell instance $2033 r0 *1 368.03,99.4
X$2033 2622 763 25 44 2644 NOR2_X1
* cell instance $2036 m0 *1 369.17,99.4
X$2036 2146 2585 25 44 2495 XNOR2_X2
* cell instance $2040 m0 *1 390.07,99.4
X$2040 2331 2591 2623 44 25 2597 OAI21_X2
* cell instance $2042 m0 *1 392.16,99.4
X$2042 2549 2649 1625 25 44 2594 NAND3_X2
* cell instance $2044 m0 *1 396.53,99.4
X$2044 2592 2015 2676 2348 25 44 2625 AOI211_X4
* cell instance $2046 m0 *1 399.38,99.4
X$2046 2597 2307 25 44 2598 NOR2_X1
* cell instance $2052 r0 *1 377.15,99.4
X$2052 2588 2343 25 44 2645 NOR2_X2
* cell instance $2056 r0 *1 380.57,99.4
X$2056 2589 2415 25 44 2671 NAND2_X1
* cell instance $2060 r0 *1 384.75,99.4
X$2060 2064 2063 2671 44 2646 25 OAI21_X1
* cell instance $2063 r0 *1 386.08,99.4
X$2063 2017 2065 2586 25 44 2647 NAND3_X1
* cell instance $2067 r0 *1 390.83,99.4
X$2067 2591 2623 2422 25 44 NOR2_X4
* cell instance $2073 r0 *1 398.43,99.4
X$2073 2650 2624 2721 2678 1765 2151 25 44 OAI221_X2
* cell instance $2076 r0 *1 401.66,99.4
X$2076 2349 2381 2595 44 25 2677 AND3_X2
* cell instance $2077 r0 *1 402.8,99.4
X$2077 2595 2381 2349 25 44 2652 NAND3_X2
* cell instance $2081 r0 *1 406.22,99.4
X$2081 25 2627 2626 2675 2486 1765 44 AOI22_X4
* cell instance $2083 m0 *1 406.41,99.4
X$2083 2639 2529 25 44 2600 NAND2_X2
* cell instance $2088 r0 *1 410.78,99.4
X$2088 2639 44 2527 25 BUF_X4
* cell instance $2089 m0 *1 410.97,99.4
X$2089 25 2228 2067 2628 2629 2620 44 NAND4_X4
* cell instance $2092 m0 *1 414.58,99.4
X$2092 2629 2628 2530 25 44 2638 NAND3_X1
* cell instance $2094 r0 *1 412.11,99.4
X$2094 25 2602 2626 2655 2656 44 AOI21_X4
* cell instance $2096 m0 *1 418.19,99.4
X$2096 2603 2530 25 2073 44 NAND2_X4
* cell instance $2097 m0 *1 415.72,99.4
X$2097 25 2603 2620 2602 2601 44 AOI21_X4
* cell instance $2098 m0 *1 419.9,99.4
X$2098 2638 25 44 2604 INV_X1
* cell instance $2103 m0 *1 428.83,99.4
X$2103 1948 1949 25 44 2432 NAND2_X2
* cell instance $2105 r0 *1 417.62,99.4
X$2105 2530 2603 44 25 2672 AND2_X1
* cell instance $2106 r0 *1 418.38,99.4
X$2106 2672 44 2021 25 BUF_X4
* cell instance $2108 r0 *1 419.9,99.4
X$2108 2630 25 44 729 INV_X4
* cell instance $2109 r0 *1 420.85,99.4
X$2109 2630 44 1932 25 BUF_X4
* cell instance $2113 r0 *1 424.65,99.4
X$2113 1932 2734 25 44 2564 OR2_X1
* cell instance $2116 r0 *1 427.12,99.4
X$2116 2379 1932 25 44 2433 XNOR2_X2
* cell instance $2119 r0 *1 429.59,99.4
X$2119 2702 2669 25 44 2277 NAND2_X1
* cell instance $2121 m0 *1 430.16,99.4
X$2121 2563 2433 2503 44 25 2632 AND3_X1
* cell instance $2122 m0 *1 431.11,99.4
X$2122 25 2632 2215 1892 2432 2633 44 AND4_X4
* cell instance $2126 m0 *1 436.05,99.4
X$2126 25 2353 2631 2043 2633 2637 44 NOR4_X4
* cell instance $2128 m0 *1 440.99,99.4
X$2128 25 1893 44 2538 BUF_X8
* cell instance $2130 r0 *1 430.35,99.4
X$2130 2661 2657 2317 44 2669 25 OAI21_X1
* cell instance $2131 r0 *1 431.11,99.4
X$2131 2632 2215 1892 2432 25 44 2657 NAND4_X1
* cell instance $2135 r0 *1 433.39,99.4
X$2135 25 2606 2633 2539 2658 2044 44 NAND4_X4
* cell instance $2137 r0 *1 437.57,99.4
X$2137 2658 2633 2631 44 25 2518 OAI21_X2
* cell instance $2139 r0 *1 439.28,99.4
X$2139 2606 2661 25 44 2170 NOR2_X2
* cell instance $2140 r0 *1 440.23,99.4
X$2140 2660 2567 25 44 2608 NOR2_X1
* cell instance $2142 r0 *1 441.18,99.4
X$2142 2660 2634 2667 25 44 2664 MUX2_X1
* cell instance $2143 r0 *1 442.51,99.4
X$2143 2539 2635 25 44 2667 OR2_X1
* cell instance $2144 r0 *1 443.27,99.4
X$2144 2635 2661 25 44 2662 NOR2_X1
* cell instance $2145 m0 *1 444.03,99.4
X$2145 2635 2567 25 44 2570 NAND2_X1
* cell instance $2196 r0 *1 443.84,99.4
X$2196 2634 2662 2633 2631 2636 25 44 OAI211_X2
* cell instance $2197 r0 *1 445.55,99.4
X$2197 2663 2664 2636 25 44 2512 NAND3_X1
* cell instance $2199 r0 *1 446.69,99.4
X$2199 2636 2664 2663 44 25 2474 AND3_X1
* cell instance $2382 m0 *1 369.74,51.8
X$2382 1209 1020 1208 25 1269 44 NAND3_X4
* cell instance $2383 r0 *1 369.74,51.8
X$2383 1248 1209 1020 1208 25 1357 44 NAND4_X2
* cell instance $2386 r0 *1 372.4,51.8
X$2386 1292 1061 1358 44 1301 25 NOR3_X2
* cell instance $2387 m0 *1 373.92,51.8
X$2387 978 870 1253 1211 1250 25 44 OAI211_X2
* cell instance $2388 m0 *1 372.59,51.8
X$2388 1250 1251 1210 44 25 1270 OAI21_X2
* cell instance $2392 r0 *1 374.49,51.8
X$2392 1253 1211 25 44 1311 NOR2_X2
* cell instance $2393 r0 *1 375.44,51.8
X$2393 25 1211 1152 1271 1112 44 NOR3_X4
* cell instance $2395 m0 *1 377.53,51.8
X$2395 1153 1064 1154 25 44 1248 OR3_X2
* cell instance $2396 m0 *1 378.86,51.8
X$2396 25 1153 1064 1154 1241 44 NOR3_X4
* cell instance $2401 m0 *1 386.08,51.8
X$2401 1158 1212 25 44 1272 XNOR2_X2
* cell instance $2402 m0 *1 384.18,51.8
X$2402 1255 1155 25 44 1425 XNOR2_X2
* cell instance $2406 r0 *1 384.18,51.8
X$2406 25 1361 1273 1301 1295 44 AOI21_X4
* cell instance $2411 m0 *1 390.64,51.8
X$2411 1274 1065 44 25 1114 AND2_X1
* cell instance $2412 r0 *1 390.64,51.8
X$2412 1065 1274 25 44 1273 NAND2_X1
* cell instance $2414 r0 *1 391.59,51.8
X$2414 1273 1213 25 44 1316 NAND2_X1
* cell instance $2415 m0 *1 392.35,51.8
X$2415 1159 1213 1214 25 44 1215 NAND3_X2
* cell instance $2416 m0 *1 391.78,51.8
X$2416 1213 1214 25 44 1157 NAND2_X1
* cell instance $2419 m0 *1 394.44,51.8
X$2419 1213 1159 25 44 1275 XNOR2_X2
* cell instance $2420 m0 *1 394.06,51.8
X$2420 1257 25 44 1213 INV_X1
* cell instance $2425 r0 *1 399,51.8
X$2425 1358 25 44 1317 INV_X2
* cell instance $2427 m0 *1 399,51.8
X$2427 1275 25 44 967 CLKBUF_X3
* cell instance $2429 m0 *1 400.9,51.8
X$2429 981 967 25 44 1276 NOR2_X1
* cell instance $2430 m0 *1 401.47,51.8
X$2430 915 1277 1216 44 1259 25 OAI21_X1
* cell instance $2432 m0 *1 402.42,51.8
X$2432 1217 915 982 25 44 1216 NAND3_X1
* cell instance $2433 m0 *1 403.18,51.8
X$2433 751 1100 25 44 1217 NOR2_X1
* cell instance $2436 r0 *1 401.09,51.8
X$2436 1276 1386 1217 25 1277 44 AOI21_X1
* cell instance $2437 r0 *1 401.85,51.8
X$2437 1217 1276 915 1274 1317 44 25 1069 OAI221_X1
* cell instance $2439 r0 *1 403.37,51.8
X$2439 987 1025 44 25 1279 XNOR2_X1
* cell instance $2440 m0 *1 404.32,51.8
X$2440 1279 751 1100 44 1278 25 NOR3_X2
* cell instance $2445 r0 *1 404.7,51.8
X$2445 1025 981 967 44 1318 25 NOR3_X2
* cell instance $2447 m0 *1 407.74,51.8
X$2447 1366 1025 981 25 44 1219 NOR3_X1
* cell instance $2448 m0 *1 406.79,51.8
X$2448 982 981 1218 25 44 1262 OR3_X1
* cell instance $2451 m0 *1 409.45,51.8
X$2451 1220 1222 1254 25 44 NOR2_X4
* cell instance $2454 m0 *1 412.11,51.8
X$2454 1222 633 25 44 1074 XNOR2_X2
* cell instance $2455 m0 *1 414.01,51.8
X$2455 1300 1162 1299 25 44 1369 MUX2_X1
* cell instance $2456 m0 *1 415.34,51.8
X$2456 1221 1281 1220 25 44 1298 NOR3_X1
* cell instance $2460 r0 *1 409.26,51.8
X$2460 1280 1386 25 44 1366 NOR2_X1
* cell instance $2461 r0 *1 409.83,51.8
X$2461 1280 982 25 44 987 NAND2_X2
* cell instance $2465 r0 *1 413.25,51.8
X$2465 1320 1319 1258 25 44 1075 MUX2_X1
* cell instance $2466 r0 *1 414.58,51.8
X$2466 1074 1321 25 44 1299 NOR2_X1
* cell instance $2469 r0 *1 415.72,51.8
X$2469 1368 1319 1369 25 920 44 AOI21_X2
* cell instance $2470 r0 *1 417.05,51.8
X$2470 1281 1163 1389 44 1362 25 OAI21_X1
* cell instance $2472 m0 *1 419.71,51.8
X$2472 1256 633 1297 25 1221 44 AOI21_X2
* cell instance $2476 m0 *1 421.99,51.8
X$2476 1282 25 44 1297 INV_X1
* cell instance $2479 r0 *1 421.23,51.8
X$2479 1191 25 44 1281 INV_X2
* cell instance $2480 r0 *1 421.8,51.8
X$2480 25 1323 1282 1283 1365 1284 44 OAI22_X4
* cell instance $2481 m0 *1 422.94,51.8
X$2481 1223 1222 25 44 1283 NAND2_X2
* cell instance $2483 m0 *1 423.89,51.8
X$2483 1283 1284 25 44 1256 NOR2_X1
* cell instance $2486 m0 *1 424.84,51.8
X$2486 25 1165 1294 1222 1164 44 AOI21_X4
* cell instance $2488 r0 *1 425.22,51.8
X$2488 1362 1354 44 883 25 XOR2_X2
* cell instance $2490 m0 *1 427.88,51.8
X$2490 1286 25 44 1294 INV_X1
* cell instance $2495 m0 *1 440.61,51.8
X$2495 1228 1227 1229 25 1287 44 AOI21_X2
* cell instance $2499 r0 *1 427.69,51.8
X$2499 1325 25 44 1328 INV_X1
* cell instance $2500 r0 *1 428.07,51.8
X$2500 1285 1328 1119 1286 25 44 1224 AOI22_X1
* cell instance $2501 r0 *1 429.02,51.8
X$2501 1122 1293 1325 25 1284 44 AOI21_X2
* cell instance $2502 r0 *1 430.35,51.8
X$2502 1285 1325 25 44 1356 NOR2_X1
* cell instance $2503 r0 *1 430.92,51.8
X$2503 1286 1119 25 44 1331 NAND2_X1
* cell instance $2507 r0 *1 433.58,51.8
X$2507 1348 1173 44 1293 25 XOR2_X2
* cell instance $2510 r0 *1 439.09,51.8
X$2510 1227 1032 1082 44 25 1345 OAI21_X2
* cell instance $2512 r0 *1 440.61,51.8
X$2512 1229 1227 25 44 1334 NAND2_X1
* cell instance $2513 r0 *1 441.18,51.8
X$2513 1342 1444 1172 25 1337 44 AOI21_X1
* cell instance $2515 m0 *1 444.79,51.8
X$2515 1230 999 725 25 44 1288 NAND3_X1
* cell instance $2517 m0 *1 445.55,51.8
X$2517 25 1032 1228 1290 1128 44 AOI21_X4
* cell instance $2520 m0 *1 454.29,51.8
X$2520 1130 1230 1179 1231 25 44 1232 NAND4_X1
* cell instance $2523 m0 *1 456.19,51.8
X$2523 1230 1130 44 25 1131 XNOR2_X1
* cell instance $2574 r0 *1 444.98,51.8
X$2574 1288 1289 25 44 1342 NAND2_X1
* cell instance $2575 r0 *1 445.55,51.8
X$2575 1288 1289 1089 25 44 1445 NAND3_X1
* cell instance $2578 r0 *1 446.88,51.8
X$2578 725 1174 1340 25 44 1289 OR3_X1
* cell instance $2583 r0 *1 453.34,51.8
X$2583 1179 725 25 44 1338 NOR2_X1
* cell instance $2771 m0 *1 448.21,63
X$2771 1716 1573 25 44 1574 XNOR2_X2
* cell instance $2775 m0 *1 451.82,63
X$2775 1566 1621 25 44 1485 XNOR2_X2
* cell instance $2777 r0 *1 448.02,63
X$2777 1617 1659 1672 25 44 1085 OR3_X2
* cell instance $2780 r0 *1 449.73,63
X$2780 1657 1617 1666 25 1671 44 AOI21_X1
* cell instance $2783 r0 *1 452.39,63
X$2783 1894 1482 1529 25 1621 44 AOI21_X2
* cell instance $2786 m0 *1 454.1,63
X$2786 1563 680 1569 25 44 1666 MUX2_X1
* cell instance $2787 m0 *1 456.19,63
X$2787 1620 1567 1564 1568 1531 1563 44 25 AOI221_X2
* cell instance $2788 m0 *1 458.28,63
X$2788 1565 1527 1618 25 44 1567 NAND3_X1
* cell instance $2791 m0 *1 459.99,63
X$2791 1566 1487 25 44 1619 OR2_X1
* cell instance $2798 r0 *1 456.95,63
X$2798 1717 1395 1333 1490 44 1564 25 NOR4_X2
* cell instance $2799 r0 *1 458.66,63
X$2799 1660 1333 25 44 1530 NOR2_X1
* cell instance $2800 r0 *1 459.23,63
X$2800 1664 25 44 1617 CLKBUF_X3
* cell instance $2802 r0 *1 460.56,63
X$2802 1663 1662 1530 1439 1661 1619 25 44 1664 OAI33_X1
* cell instance $6782 r0 *1 631.75,211.4
X$6782 25 2891 44 598 BUF_X8
* cell instance $19571 m0 *1 809.59,376.6
X$19571 2891 25 44 2890 BUF_X1
* cell instance $29992 m0 *1 363.85,105
X$29992 2144 2358 44 25 2739 AND2_X1
* cell instance $29994 m0 *1 364.8,105
X$29994 25 1842 2739 2802 2666 2144 44 AOI22_X4
* cell instance $30025 r0 *1 368.41,105
X$30025 2666 2726 25 44 2774 OR2_X1
* cell instance $30028 r0 *1 372.4,105
X$30028 2728 1625 25 44 2775 NOR2_X1
* cell instance $30032 r0 *1 375.44,105
X$30032 2749 2728 2725 44 2788 25 OAI21_X1
* cell instance $30035 m0 *1 376.77,105
X$30035 2750 2727 2302 2670 25 2742 44 NAND4_X2
* cell instance $30037 r0 *1 376.96,105
X$30037 2302 2727 2750 2670 44 25 2776 AND4_X2
* cell instance $30038 r0 *1 378.29,105
X$30038 2750 2727 25 44 2751 NAND2_X1
* cell instance $30041 r0 *1 379.81,105
X$30041 2749 2728 2767 44 2783 25 OAI21_X1
* cell instance $30042 m0 *1 380.57,105
X$30042 2728 2586 1884 25 2746 44 AOI21_X1
* cell instance $30049 r0 *1 381.14,105
X$30049 2767 2302 25 44 2768 NAND2_X1
* cell instance $30051 r0 *1 382.47,105
X$30051 2783 2064 2768 44 25 2769 OAI21_X2
* cell instance $30054 m0 *1 386.27,105
X$30054 2586 2714 25 44 2688 XNOR2_X2
* cell instance $30058 r0 *1 387.03,105
X$30058 2715 2769 2591 2623 25 44 2831 NOR4_X1
* cell instance $30060 r0 *1 388.36,105
X$30060 1625 44 2685 25 BUF_X4
* cell instance $30194 m0 *1 366.13,107.8
X$30194 2679 2725 44 25 2803 AND2_X1
* cell instance $30195 m0 *1 366.89,107.8
X$30195 25 2749 2803 2824 2802 2774 44 AOI22_X4
* cell instance $30197 m0 *1 373.16,107.8
X$30197 2725 2586 2775 25 2787 44 AOI21_X1
* cell instance $30226 r0 *1 369.36,107.8
X$30226 2666 764 25 44 2786 NOR2_X1
* cell instance $30227 r0 *1 369.93,107.8
X$30227 2786 2679 2804 2666 2144 2789 44 25 AOI221_X2
* cell instance $30230 r0 *1 372.59,107.8
X$30230 1884 2679 25 44 2804 NOR2_X1
* cell instance $30232 r0 *1 373.35,107.8
X$30232 2725 2679 25 44 2817 NOR2_X1
* cell instance $30234 m0 *1 374.49,107.8
X$30234 2767 2680 25 44 2826 NAND2_X1
* cell instance $30236 m0 *1 375.06,107.8
X$30236 2787 2680 25 44 2791 NAND2_X1
* cell instance $30243 r0 *1 375.25,107.8
X$30243 2787 1884 2818 25 44 2805 MUX2_X1
* cell instance $30245 r0 *1 376.77,107.8
X$30245 2805 2742 25 44 2790 NAND2_X1
* cell instance $30247 r0 *1 377.72,107.8
X$30247 2805 2790 2789 44 25 2797 MUX2_X2
* cell instance $30249 r0 *1 379.62,107.8
X$30249 2806 2789 2790 25 2809 44 AOI21_X2
* cell instance $30435 m0 *1 386.27,113.4
X$30435 2852 2853 2851 44 25 2860 AND3_X1
* cell instance $30437 m0 *1 387.22,113.4
X$30437 2852 2851 2853 25 2859 44 AOI21_X1
* cell instance $30438 m0 *1 387.98,113.4
X$30438 2851 2853 2852 25 44 2847 NAND3_X1
* cell instance $30441 m0 *1 390.07,113.4
X$30441 2861 2755 2860 2863 2859 2862 44 25 AOI221_X2
* cell instance $30453 m0 *1 397.29,113.4
X$30453 2862 44 2529 25 BUF_X4
* cell instance $30455 m0 *1 398.62,113.4
X$30455 2855 2854 2856 2720 44 25 2865 AND4_X1
* cell instance $30456 m0 *1 399.76,113.4
X$30456 2331 757 25 44 2837 XNOR2_X2
* cell instance $30457 m0 *1 401.66,113.4
X$30457 2816 2422 2755 25 2876 44 AOI21_X1
* cell instance $30458 m0 *1 402.42,113.4
X$30458 2855 2333 2677 25 2857 44 AOI21_X2
* cell instance $30459 m0 *1 403.75,113.4
X$30459 2595 2837 44 25 2866 AND2_X1
* cell instance $30463 r0 *1 397.1,113.4
X$30463 25 2856 2720 2855 2854 2836 44 NAND4_X4
* cell instance $30467 m0 *1 408.69,113.4
X$30467 2865 639 2527 44 2849 25 OAI21_X1
* cell instance $30469 m0 *1 409.83,113.4
X$30469 2722 2527 2018 25 44 2858 NAND3_X2
* cell instance $30470 m0 *1 411.92,113.4
X$30470 2858 2529 2086 25 2864 44 AOI21_X2
* cell instance $30473 m0 *1 416.1,113.4
X$30473 2839 44 1951 25 BUF_X4
* cell instance $30474 m0 *1 413.63,113.4
X$30474 25 1999 2864 1951 2871 44 AOI21_X4
* cell instance $30756 m0 *1 372.21,110.6
X$30756 2775 2586 25 44 2829 NAND2_X1
* cell instance $30757 m0 *1 372.78,110.6
X$30757 2586 2775 44 25 2825 AND2_X1
* cell instance $30759 m0 *1 373.73,110.6
X$30759 2825 1884 2826 2776 2827 44 25 AOI211_X2
* cell instance $30760 m0 *1 375.44,110.6
X$30760 2820 2819 2788 44 25 2818 AND3_X1
* cell instance $30761 m0 *1 376.39,110.6
X$30761 2819 2820 2824 25 2294 44 NAND3_X4
* cell instance $30762 m0 *1 378.86,110.6
X$30762 2820 2819 2824 44 25 2811 AND3_X1
* cell instance $30763 m0 *1 379.81,110.6
X$30763 2331 2711 2684 44 25 2820 OAI21_X4
* cell instance $30792 r0 *1 372.59,110.6
X$30792 764 2829 2817 2742 2853 25 44 OAI211_X2
* cell instance $30796 r0 *1 376.39,110.6
X$30796 2819 2824 44 25 2840 AND2_X1
* cell instance $30797 r0 *1 377.15,110.6
X$30797 1884 2820 2742 2840 2851 25 44 OAI211_X2
* cell instance $30798 r0 *1 378.86,110.6
X$30798 2824 2819 25 44 2841 NAND2_X1
* cell instance $30801 r0 *1 381.71,110.6
X$30801 2842 764 2776 2841 2843 44 25 AOI211_X2
* cell instance $30802 m0 *1 382.85,110.6
X$30802 2711 2684 25 44 2830 NOR2_X1
* cell instance $30808 m0 *1 391.97,110.6
X$30808 2015 2616 2422 2592 44 25 2792 AND4_X2
* cell instance $30809 m0 *1 393.3,110.6
X$30809 2592 2015 25 44 2832 NAND2_X1
* cell instance $30812 m0 *1 397.67,110.6
X$30812 2423 2369 2594 25 44 2854 OR3_X2
* cell instance $30816 r0 *1 383.42,110.6
X$30816 2830 2685 25 44 2842 NOR2_X1
* cell instance $30819 r0 *1 384.56,110.6
X$30819 2843 2827 2715 2769 44 25 2845 OAI22_X2
* cell instance $30822 r0 *1 386.84,110.6
X$30822 2715 2769 25 44 2852 NOR2_X1
* cell instance $30823 r0 *1 387.41,110.6
X$30823 2616 2831 44 25 2861 AND2_X1
* cell instance $30825 r0 *1 388.36,110.6
X$30825 2831 2616 25 44 2846 NAND2_X1
* cell instance $30828 r0 *1 389.88,110.6
X$30828 2792 2845 2846 2832 2847 2654 25 44 OAI221_X2
* cell instance $30831 r0 *1 392.54,110.6
X$30831 2592 2422 2616 2015 25 44 2863 NAND4_X1
* cell instance $30834 r0 *1 394.63,110.6
X$30834 2369 2423 2755 25 44 NOR2_X4
* cell instance $30837 r0 *1 397.48,110.6
X$30837 2689 2423 2369 44 25 2855 OAI21_X2
* cell instance $30839 r0 *1 399.19,110.6
X$30839 757 2685 25 44 2856 NAND2_X1
* cell instance $30840 r0 *1 399.76,110.6
X$30840 2832 757 25 44 2833 NOR2_X1
* cell instance $30841 r0 *1 400.33,110.6
X$30841 2689 2833 44 25 2838 XNOR2_X1
* cell instance $30844 r0 *1 402.04,110.6
X$30844 2689 2755 25 44 2834 XNOR2_X2
* cell instance $30845 m0 *1 403.18,110.6
X$30845 25 2731 2821 2754 2834 44 AOI21_X4
* cell instance $30851 r0 *1 403.94,110.6
X$30851 2834 2333 2677 25 2850 44 AOI21_X2
* cell instance $30853 r0 *1 405.65,110.6
X$30853 2857 2018 2068 25 2835 44 AOI21_X1
* cell instance $30854 r0 *1 406.41,110.6
X$30854 2884 2835 2086 2486 2844 25 44 OAI211_X2
* cell instance $30857 r0 *1 408.69,110.6
X$30857 2836 2486 25 44 2848 NAND2_X1
* cell instance $30859 r0 *1 409.45,110.6
X$30859 2527 2848 2849 44 2760 25 OAI21_X1
* cell instance $30861 r0 *1 410.59,110.6
X$30861 2582 2844 25 44 2761 XNOR2_X2
* cell instance $30863 m0 *1 411.35,110.6
X$30863 25 2858 2828 2875 2047 2134 44 OAI22_X4
* cell instance $30869 r0 *1 413.44,110.6
X$30869 2018 2695 2068 44 25 2839 OAI21_X2
* cell instance $30872 r0 *1 415.34,110.6
X$30872 2839 25 44 2134 INV_X4
* cell instance $30876 r0 *1 417.62,110.6
X$30876 2838 25 44 2807 INV_X1
* cell instance $30877 r0 *1 418,110.6
X$30877 2134 44 639 25 BUF_X4
* cell instance $30879 m0 *1 420.47,110.6
X$30879 639 2837 2807 25 44 2823 OR3_X1
* cell instance $30881 m0 *1 421.42,110.6
X$30881 639 2807 2837 44 2822 25 OAI21_X1
* cell instance $30882 m0 *1 422.18,110.6
X$30882 2073 2822 2823 25 2763 44 AOI21_X2
* cell instance $30884 m0 *1 423.7,110.6
X$30884 2823 2822 44 25 2782 AND2_X1
* cell instance $31204 m0 *1 403.18,116.2
X$31204 2836 2582 2653 25 44 2879 NAND3_X1
* cell instance $31246 r0 *1 403.94,116.2
X$31246 2876 2821 25 44 2880 NOR2_X1
* cell instance $31247 m0 *1 405.65,116.2
X$31247 2226 2333 2866 44 25 2869 AND3_X1
* cell instance $31248 m0 *1 404.32,116.2
X$31248 2866 2333 2226 25 44 2867 NAND3_X2
* cell instance $31249 m0 *1 406.6,116.2
X$31249 2784 2877 2869 2868 2878 25 44 OAI211_X2
* cell instance $31250 m0 *1 408.31,116.2
X$31250 2865 2722 2527 25 44 2877 NOR3_X1
* cell instance $31251 m0 *1 409.07,116.2
X$31251 2865 2527 25 44 2870 NAND2_X1
* cell instance $31254 r0 *1 404.89,116.2
X$31254 2821 2876 25 44 2868 OR2_X1
* cell instance $31257 r0 *1 406.22,116.2
X$31257 2867 2880 25 44 2884 NAND2_X1
* cell instance $31260 r0 *1 407.36,116.2
X$31260 2868 2869 2784 44 2883 25 OAI21_X1
* cell instance $31262 r0 *1 408.5,116.2
X$31262 2870 2878 2882 2872 2871 25 44 OAI211_X2
* cell instance $31264 m0 *1 410.02,116.2
X$31264 2722 2653 25 44 2872 NAND2_X1
* cell instance $31265 m0 *1 410.78,116.2
X$31265 2836 2653 25 44 2873 NOR2_X1
* cell instance $31267 m0 *1 411.54,116.2
X$31267 2582 2527 25 44 2874 NOR2_X1
* cell instance $31283 r0 *1 410.78,116.2
X$31283 2881 2873 2883 2874 2875 44 25 AOI211_X2
* cell instance $31570 m0 *1 403.37,119
X$31570 2879 2857 2867 2880 2881 44 25 AOI211_X2
* cell instance $31572 m0 *1 405.84,119
X$31572 2857 2880 2867 25 2882 44 AOI21_X1
* cell instance $34582 m0 *1 165.3,203
X$34582 25 1003 44 2889 BUF_X8
* cell instance $35268 m0 *1 165.11,191.8
X$35268 25 786 44 2885 BUF_X8
* cell instance $35284 r0 *1 169.48,191.8
X$35284 25 727 44 2886 BUF_X8
* cell instance $38685 m0 *1 167.01,194.6
X$38685 25 819 44 2887 BUF_X8
* cell instance $38791 r0 *1 175.56,194.6
X$38791 25 1037 44 2888 BUF_X8
* cell instance $41647 m0 *1 352.26,85.4
X$41647 25 2264 2259 2093 2238 44 AOI21_X4
* cell instance $41648 m0 *1 354.73,85.4
X$41648 2238 2093 2259 2055 2237 2260 44 25 AOI221_X2
* cell instance $41650 m0 *1 357.58,85.4
X$41650 2055 25 44 1879 INV_X4
* cell instance $41654 m0 *1 363.28,85.4
X$41654 2261 2213 2262 44 25 2256 OAI21_X4
* cell instance $41655 m0 *1 365.75,85.4
X$41655 2262 2261 2264 25 44 2267 NAND3_X1
* cell instance $41678 r0 *1 350.36,85.4
X$41678 1669 2006 25 44 2297 NOR2_X1
* cell instance $41682 r0 *1 352.26,85.4
X$41682 2055 44 1759 25 BUF_X4
* cell instance $41685 r0 *1 354.73,85.4
X$41685 2006 2169 2323 44 25 2324 OAI21_X2
* cell instance $41686 r0 *1 356.06,85.4
X$41686 1669 1667 25 44 2323 NOR2_X1
* cell instance $41688 r0 *1 357.01,85.4
X$41688 2324 1879 2337 25 44 NOR2_X4
* cell instance $41691 r0 *1 359.67,85.4
X$41691 1879 44 877 25 BUF_X4
* cell instance $41694 r0 *1 361.38,85.4
X$41694 25 2222 2103 2223 2414 2101 44 OAI211_X4
* cell instance $41695 r0 *1 364.61,85.4
X$41695 2263 2184 2101 2264 2339 2340 44 25 AOI221_X2
* cell instance $41697 r0 *1 366.89,85.4
X$41697 2298 2101 1748 2265 44 2325 25 NOR4_X2
* cell instance $41698 m0 *1 367.84,85.4
X$41698 1728 1799 2265 25 44 NOR2_X4
* cell instance $41700 m0 *1 369.55,85.4
X$41700 2287 44 2146 25 BUF_X4
* cell instance $41703 m0 *1 377.72,85.4
X$41703 2256 2249 44 25 2302 AND2_X2
* cell instance $41704 m0 *1 378.67,85.4
X$41704 25 2269 2290 2327 2289 44 AOI21_X4
* cell instance $41705 m0 *1 381.14,85.4
X$41705 2249 2256 25 2347 44 NAND2_X4
* cell instance $41712 r0 *1 371.45,85.4
X$41712 2266 2326 25 44 2298 NAND2_X2
* cell instance $41713 r0 *1 372.4,85.4
X$41713 1625 2266 2326 25 2299 44 AOI21_X1
* cell instance $41715 r0 *1 373.35,85.4
X$41715 2266 2326 1411 25 44 2300 NAND3_X1
* cell instance $41716 r0 *1 374.11,85.4
X$41716 1411 44 2331 25 BUF_X4
* cell instance $41719 r0 *1 378.86,85.4
X$41719 1737 2268 25 44 2327 NOR2_X2
* cell instance $41720 r0 *1 379.81,85.4
X$41720 2101 2103 1907 44 2301 25 NOR3_X2
* cell instance $41724 r0 *1 383.8,85.4
X$41724 2012 2302 44 25 2364 AND2_X1
* cell instance $41725 r0 *1 384.56,85.4
X$41725 2302 2012 25 44 2303 NAND2_X1
* cell instance $41726 r0 *1 385.13,85.4
X$41726 2216 2012 25 44 2344 NOR2_X1
* cell instance $41727 r0 *1 385.7,85.4
X$41727 2012 2216 25 44 2304 OR2_X1
* cell instance $41729 m0 *1 386.27,85.4
X$41729 2059 1461 25 44 2329 NAND2_X1
* cell instance $41732 r0 *1 386.65,85.4
X$41732 2188 1498 25 44 2376 NOR2_X1
* cell instance $41734 r0 *1 387.98,85.4
X$41734 2345 2305 2329 1333 1426 2188 25 44 2306 OAI33_X1
* cell instance $41735 m0 *1 388.17,85.4
X$41735 2216 2012 25 44 2270 NAND2_X1
* cell instance $41737 m0 *1 388.74,85.4
X$41737 2270 2059 1415 25 44 2292 NAND3_X2
* cell instance $41741 m0 *1 394.06,85.4
X$41741 2064 2063 2187 44 2420 25 OAI21_X1
* cell instance $41742 m0 *1 394.82,85.4
X$41742 2188 2294 2295 44 25 2296 OAI21_X2
* cell instance $41748 r0 *1 393.49,85.4
X$41748 2271 2065 2017 25 2368 44 AOI21_X2
* cell instance $41751 m0 *1 398.24,85.4
X$41751 25 2135 2296 1083 2307 2272 44 NAND4_X4
* cell instance $41754 m0 *1 403.18,85.4
X$41754 2272 2220 2225 25 2273 44 NAND3_X4
* cell instance $41756 m0 *1 406.41,85.4
X$41756 2220 2272 44 25 2309 AND2_X1
* cell instance $41757 m0 *1 407.17,85.4
X$41757 2225 2272 25 44 2274 NAND2_X2
* cell instance $41762 m0 *1 413.63,85.4
X$41762 2293 1426 25 44 2275 NOR2_X2
* cell instance $41763 m0 *1 414.58,85.4
X$41763 25 2312 2274 2275 1951 44 AOI21_X4
* cell instance $41764 m0 *1 417.05,85.4
X$41764 2275 25 44 2291 INV_X1
* cell instance $41771 r0 *1 400.33,85.4
X$41771 2307 1927 2110 25 2381 44 NAND3_X4
* cell instance $41775 r0 *1 406.41,85.4
X$41775 2309 2310 1686 2225 25 2308 44 NAND4_X2
* cell instance $41779 r0 *1 412.3,85.4
X$41779 25 1426 2293 2311 2334 44 NOR3_X4
* cell instance $41780 r0 *1 414.96,85.4
X$41780 2274 25 44 2311 INV_X2
* cell instance $41783 r0 *1 417.24,85.4
X$41783 1461 2351 2312 44 25 2314 OAI21_X4
* cell instance $41785 r0 *1 420.47,85.4
X$41785 2313 2230 25 44 2332 NAND2_X1
* cell instance $41788 r0 *1 424.46,85.4
X$41788 2116 2314 25 44 2330 NOR2_X2
* cell instance $41789 r0 *1 425.41,85.4
X$41789 2315 2116 2314 44 2400 25 NOR3_X2
* cell instance $41790 m0 *1 426.36,85.4
X$41790 1498 2197 2157 25 2276 44 AOI21_X2
* cell instance $41792 m0 *1 427.69,85.4
X$41792 2288 2276 2158 25 2328 44 AOI21_X2
* cell instance $41793 m0 *1 429.02,85.4
X$41793 2277 2317 2067 25 44 2075 NAND3_X1
* cell instance $41794 m0 *1 429.78,85.4
X$41794 2277 2286 25 44 2131 NAND2_X2
* cell instance $41798 r0 *1 426.74,85.4
X$41798 2314 2116 2315 25 44 2316 OR3_X1
* cell instance $41800 m0 *1 433.58,85.4
X$41800 1893 2023 2276 25 44 2242 NAND3_X1
* cell instance $41802 m0 *1 434.34,85.4
X$41802 2286 2317 2044 25 44 2280 NAND3_X1
* cell instance $41808 r0 *1 434.15,85.4
X$41808 2044 2317 2286 44 25 2320 AND3_X2
* cell instance $41810 r0 *1 436.05,85.4
X$41810 1947 2637 2506 44 25 1863 OAI21_X4
* cell instance $41812 m0 *1 444.22,85.4
X$41812 2280 2233 2318 25 44 2208 MUX2_X1
* cell instance $41813 m0 *1 440.8,85.4
X$41813 25 2278 1863 1775 2279 2318 44 NOR4_X4
* cell instance $41817 m0 *1 449.54,85.4
X$41817 25 1863 1775 2279 2281 44 NOR3_X4
* cell instance $41818 m0 *1 452.2,85.4
X$41818 2284 2281 44 2282 25 XOR2_X2
* cell instance $41819 m0 *1 453.91,85.4
X$41819 2229 2285 2282 2233 2235 2321 25 44 2080 OAI33_X1
* cell instance $41820 m0 *1 455.24,85.4
X$41820 1898 2285 1416 44 25 1718 MUX2_X2
* cell instance $41821 m0 *1 456.95,85.4
X$41821 2284 2322 25 44 1528 XNOR2_X2
* cell instance $41873 r0 *1 446.31,85.4
X$41873 2319 2233 2320 2239 25 44 2207 OR4_X1
* cell instance $41877 r0 *1 449.92,85.4
X$41877 2396 44 1857 25 BUF_X4
* cell instance $41881 r0 *1 452.58,85.4
X$41881 25 2229 2281 2235 2322 2233 44 OAI22_X4
* cell instance $41882 r0 *1 455.81,85.4
X$41882 2321 1898 25 44 2283 NOR2_X1
* cell instance $41886 r0 *1 457.71,85.4
X$41886 2322 2284 44 1779 25 XOR2_X2
* cell instance $42144 r0 *1 350.17,88.2
X$42144 1740 2006 25 44 2370 NOR2_X1
* cell instance $42145 m0 *1 351.31,88.2
X$42145 2297 2335 2055 44 25 2338 MUX2_X2
* cell instance $42146 m0 *1 350.36,88.2
X$42146 1667 2141 2370 44 25 2335 AND3_X1
* cell instance $42147 m0 *1 353.02,88.2
X$42147 2005 2141 1759 44 2336 25 OAI21_X1
* cell instance $42149 m0 *1 353.97,88.2
X$42149 877 2006 2005 25 2355 44 AOI21_X2
* cell instance $42154 r0 *1 352.26,88.2
X$42154 2398 2006 2336 25 2371 44 AOI21_X2
* cell instance $42155 r0 *1 353.59,88.2
X$42155 2457 877 2006 25 44 2398 NOR3_X1
* cell instance $42158 r0 *1 355.3,88.2
X$42158 1669 2355 25 44 2459 XNOR2_X2
* cell instance $42160 m0 *1 358.15,88.2
X$42160 2337 2338 2356 2182 2008 2358 25 44 2458 OAI33_X1
* cell instance $42164 m0 *1 360.43,88.2
X$42164 2337 2338 25 44 2339 NOR2_X2
* cell instance $42168 r0 *1 358.91,88.2
X$42168 2222 2338 2337 44 25 2183 OAI21_X2
* cell instance $42172 r0 *1 362.71,88.2
X$42172 2145 1876 1581 44 2358 25 NOR3_X2
* cell instance $42174 m0 *1 363.28,88.2
X$42174 2461 2339 25 44 2261 NOR2_X2
* cell instance $42177 r0 *1 364.04,88.2
X$42177 2145 1876 2517 25 44 NOR2_X4
* cell instance $42180 r0 *1 367.65,88.2
X$42180 2401 2146 2185 25 44 2372 NAND3_X2
* cell instance $42181 r0 *1 368.98,88.2
X$42181 2103 1581 25 44 2443 NAND2_X2
* cell instance $42183 m0 *1 371.64,88.2
X$42183 2298 1625 25 44 2341 NOR2_X1
* cell instance $42185 m0 *1 372.21,88.2
X$42185 2341 2299 2340 44 25 2415 MUX2_X2
* cell instance $42188 m0 *1 376.01,88.2
X$42188 2298 2331 25 44 2360 NAND2_X1
* cell instance $42189 m0 *1 374.3,88.2
X$42189 2300 2360 2340 44 25 2343 MUX2_X2
* cell instance $42192 r0 *1 374.68,88.2
X$42192 2298 2340 25 44 2494 XNOR2_X2
* cell instance $42194 m0 *1 377.15,88.2
X$42194 2268 44 763 25 BUF_X4
* cell instance $42199 m0 *1 379.62,88.2
X$42199 25 2588 2301 2289 2251 44 AOI21_X4
* cell instance $42200 m0 *1 383.61,88.2
X$42200 2364 2065 2363 2344 2405 2366 44 25 AOI221_X2
* cell instance $42201 m0 *1 385.7,88.2
X$42201 2304 2345 2305 25 44 2363 NOR3_X1
* cell instance $42205 r0 *1 380.76,88.2
X$42205 2302 2404 2403 44 25 2063 OAI21_X4
* cell instance $42206 r0 *1 383.23,88.2
X$42206 2403 2404 25 44 2405 NOR2_X1
* cell instance $42207 r0 *1 383.8,88.2
X$42207 2304 2373 2303 2064 2407 2412 25 44 OAI221_X2
* cell instance $42208 r0 *1 385.89,88.2
X$42208 2344 2374 2406 25 44 2407 NAND3_X1
* cell instance $42209 r0 *1 386.65,88.2
X$42209 2376 2374 2375 25 2411 44 AOI21_X2
* cell instance $42210 m0 *1 387.03,88.2
X$42210 25 2346 2409 2347 2292 2367 44 NOR4_X4
* cell instance $42215 r0 *1 388.17,88.2
X$42215 2418 2377 25 44 2409 NOR2_X2
* cell instance $42216 r0 *1 389.12,88.2
X$42216 2346 2409 2347 2292 25 44 2421 OR4_X1
* cell instance $42217 r0 *1 390.26,88.2
X$42217 1360 2411 2419 25 2378 44 AOI21_X2
* cell instance $42218 m0 *1 391.78,88.2
X$42218 25 2366 2378 2367 2369 2368 44 OAI211_X4
* cell instance $42222 m0 *1 396.72,88.2
X$42222 2307 44 1885 25 BUF_X4
* cell instance $42224 m0 *1 398.81,88.2
X$42224 2189 2348 25 44 2349 NAND2_X2
* cell instance $42229 r0 *1 394.06,88.2
X$42229 1360 44 2379 25 BUF_X4
* cell instance $42232 r0 *1 397.29,88.2
X$42232 2348 44 757 25 BUF_X4
* cell instance $42233 r0 *1 398.62,88.2
X$42233 2422 2189 2307 44 2380 25 NOR3_X2
* cell instance $42235 m0 *1 400.33,88.2
X$42235 2348 1927 2110 25 2451 44 AOI21_X2
* cell instance $42240 m0 *1 404.13,88.2
X$42240 2381 2349 25 44 2293 NAND2_X2
* cell instance $42243 m0 *1 406.03,88.2
X$42243 2333 2226 25 44 2350 NAND2_X1
* cell instance $42247 r0 *1 404.13,88.2
X$42247 2349 2381 44 25 2226 AND2_X2
* cell instance $42250 m0 *1 407.93,88.2
X$42250 1802 2068 2310 2350 25 44 2361 OR4_X1
* cell instance $42251 m0 *1 406.98,88.2
X$42251 2350 2310 2068 1802 25 44 2365 NOR4_X1
* cell instance $42253 m0 *1 409.83,88.2
X$42253 2310 2018 25 44 2362 NAND2_X1
* cell instance $42258 r0 *1 407.55,88.2
X$42258 2310 2068 2018 25 44 2382 NAND3_X1
* cell instance $42260 r0 *1 408.5,88.2
X$42260 2365 2383 2413 44 25 2384 MUX2_X2
* cell instance $42262 r0 *1 410.97,88.2
X$42262 2361 2362 2413 44 25 2426 MUX2_X2
* cell instance $42264 r0 *1 413.44,88.2
X$42264 2427 2384 2334 1951 2408 44 25 AOI211_X2
* cell instance $42266 r0 *1 415.34,88.2
X$42266 2334 25 44 2410 INV_X1
* cell instance $42267 m0 *1 415.53,88.2
X$42267 2334 1951 25 2197 44 NAND2_X4
* cell instance $42272 r0 *1 415.91,88.2
X$42272 2410 2134 2351 25 44 NOR2_X4
* cell instance $42273 r0 *1 417.62,88.2
X$42273 2312 2453 2195 2385 44 25 2452 OAI22_X2
* cell instance $42274 m0 *1 418.57,88.2
X$42274 2195 2312 2351 44 25 2359 OAI21_X2
* cell instance $42278 m0 *1 426.17,88.2
X$42278 2330 2288 2389 2352 2316 2429 25 44 OAI221_X2
* cell instance $42281 r0 *1 419.33,88.2
X$42281 2157 2408 2132 2386 25 44 2402 AOI22_X2
* cell instance $42282 r0 *1 421.04,88.2
X$42282 2132 2386 2197 2157 2387 44 25 AOI211_X2
* cell instance $42283 r0 *1 422.75,88.2
X$42283 2132 2157 2197 25 2388 44 AOI21_X2
* cell instance $42284 r0 *1 424.08,88.2
X$42284 2359 2386 729 44 2352 25 NOR3_X2
* cell instance $42285 r0 *1 425.41,88.2
X$42285 2386 729 1364 25 44 2399 NAND3_X2
* cell instance $42287 r0 *1 427.12,88.2
X$42287 2352 2389 25 44 2390 NOR2_X2
* cell instance $42290 r0 *1 431.3,88.2
X$42290 2431 2399 2023 2276 25 44 2537 AOI22_X2
* cell instance $42293 m0 *1 434.72,88.2
X$42293 1893 1976 2198 44 25 2357 OAI21_X2
* cell instance $42296 m0 *1 438.52,88.2
X$42296 2357 2390 44 2284 25 XOR2_X2
* cell instance $42301 r0 *1 436.24,88.2
X$42301 1893 2390 25 44 2481 NAND2_X1
* cell instance $42304 r0 *1 439.09,88.2
X$42304 2357 2390 2229 25 44 2441 NAND3_X1
* cell instance $42308 m0 *1 445.36,88.2
X$42308 2202 2320 25 2235 44 NAND2_X4
* cell instance $42311 m0 *1 447.26,88.2
X$42311 2392 2354 1416 2318 25 2035 44 NAND4_X2
* cell instance $42316 r0 *1 445.74,88.2
X$42316 2320 2202 44 25 2392 AND2_X1
* cell instance $42317 r0 *1 446.5,88.2
X$42317 2202 2320 2434 2391 25 44 2395 NAND4_X1
* cell instance $42320 r0 *1 449.16,88.2
X$42320 2475 2397 2393 44 25 2396 AND3_X1
* cell instance $42323 m0 *1 450.11,88.2
X$42323 2235 2354 25 44 2285 NOR2_X1
* cell instance $42326 r0 *1 451.06,88.2
X$42326 552 2395 1416 44 25 1490 MUX2_X2
* cell instance $42327 r0 *1 452.77,88.2
X$42327 25 1566 2477 2437 2394 44 AOI21_X4
* cell instance $42328 m0 *1 454.86,88.2
X$42328 1416 2284 25 44 2321 OR2_X1
* cell instance $42329 m0 *1 454.1,88.2
X$42329 2285 2321 25 44 2394 OR2_X1
* cell instance $42639 r0 *1 351.31,79.8
X$42639 25 2259 1959 2143 2142 44 AOI21_X4
* cell instance $42641 m0 *1 351.88,79.8
X$42641 2120 1747 1639 1798 25 44 2119 NAND4_X1
* cell instance $42642 m0 *1 353.59,79.8
X$42642 1798 1639 1747 2120 44 25 2169 AND4_X1
* cell instance $42647 r0 *1 354.16,79.8
X$42647 1959 25 44 2211 INV_X1
* cell instance $42649 m0 *1 357.58,79.8
X$42649 2091 44 2144 25 BUF_X4
* cell instance $42653 r0 *1 357.58,79.8
X$42653 2092 1667 1879 25 2172 44 AOI21_X1
* cell instance $42654 r0 *1 358.34,79.8
X$42654 2092 1695 25 44 2182 NOR2_X1
* cell instance $42655 r0 *1 358.91,79.8
X$42655 2183 1801 1959 25 44 1646 NAND3_X2
* cell instance $42656 m0 *1 360.24,79.8
X$42656 25 2123 2052 1512 2094 2222 44 NAND4_X4
* cell instance $42658 m0 *1 363.66,79.8
X$42658 2052 2123 2094 25 44 2095 NAND3_X1
* cell instance $42660 m0 *1 364.61,79.8
X$42660 2052 2094 25 44 2185 NAND2_X2
* cell instance $42668 r0 *1 363.66,79.8
X$42668 2145 2144 1876 44 2171 25 NOR3_X2
* cell instance $42671 r0 *1 365.56,79.8
X$42671 2096 1411 25 44 1748 NAND2_X2
* cell instance $42672 r0 *1 366.51,79.8
X$42672 25 2171 2146 2054 2223 2148 44 OAI211_X4
* cell instance $42673 m0 *1 369.17,79.8
X$42673 2053 2097 2147 1747 25 44 2125 AOI22_X2
* cell instance $42675 m0 *1 370.88,79.8
X$42675 2097 1962 1801 44 25 2148 MUX2_X2
* cell instance $42676 m0 *1 372.59,79.8
X$42676 2085 2099 2125 2129 2401 44 25 AOI211_X2
* cell instance $42677 m0 *1 374.3,79.8
X$42677 1908 1759 25 44 2098 NOR2_X1
* cell instance $42678 m0 *1 374.87,79.8
X$42678 2098 2130 2148 2054 1970 2342 25 44 OAI221_X2
* cell instance $42681 r0 *1 370.12,79.8
X$42681 2042 1411 2096 2010 44 25 2097 AND4_X1
* cell instance $42683 r0 *1 371.64,79.8
X$42683 2096 2042 25 44 2147 NAND2_X2
* cell instance $42685 m0 *1 377.53,79.8
X$42685 2100 44 2101 25 BUF_X4
* cell instance $42691 m0 *1 381.52,79.8
X$42691 1993 2056 2105 2106 2289 44 25 AOI211_X2
* cell instance $42692 m0 *1 380.76,79.8
X$42692 1735 2103 2096 25 44 2102 NAND3_X1
* cell instance $42693 m0 *1 383.23,79.8
X$42693 2106 2105 44 25 2175 AND2_X1
* cell instance $42696 r0 *1 380.95,79.8
X$42696 2102 2175 2104 1907 2103 2101 25 44 2149 OAI33_X1
* cell instance $42698 m0 *1 385.32,79.8
X$42698 2058 2013 1461 2059 25 2216 44 NAND4_X2
* cell instance $42700 m0 *1 387.03,79.8
X$42700 2058 2013 25 44 2188 NAND2_X2
* cell instance $42706 m0 *1 390.64,79.8
X$42706 2017 2048 25 2061 44 NAND2_X4
* cell instance $42709 m0 *1 394.25,79.8
X$42709 2062 1831 25 44 2133 NAND2_X1
* cell instance $42713 r0 *1 395.39,79.8
X$42713 2188 2065 2150 44 25 2219 OAI21_X2
* cell instance $42714 m0 *1 396.15,79.8
X$42714 25 2135 2107 2061 2133 44 AOI21_X4
* cell instance $42717 r0 *1 396.72,79.8
X$42717 2150 2061 2133 25 44 2189 MUX2_X1
* cell instance $42719 r0 *1 398.43,79.8
X$42719 2177 2059 1083 44 2255 25 OAI21_X1
* cell instance $42721 m0 *1 399,79.8
X$42721 2108 2065 2017 25 2177 44 AOI21_X1
* cell instance $42722 m0 *1 400.52,79.8
X$42722 1765 2111 2109 44 25 2110 OAI21_X2
* cell instance $42728 m0 *1 407.55,79.8
X$42728 1887 2112 1802 44 2138 25 NOR3_X2
* cell instance $42729 m0 *1 406.79,79.8
X$42729 1846 2194 1626 25 44 2140 NAND3_X1
* cell instance $42733 m0 *1 409.26,79.8
X$42733 2140 2069 1539 2139 2195 44 25 AOI211_X2
* cell instance $42734 m0 *1 411.73,79.8
X$42734 25 2113 2138 1386 2132 2114 44 OAI211_X4
* cell instance $42735 m0 *1 414.96,79.8
X$42735 2113 1846 1386 2114 2137 25 44 OAI211_X2
* cell instance $42738 m0 *1 418.38,79.8
X$42738 1846 2134 25 44 2071 NAND2_X1
* cell instance $42745 r0 *1 410.97,79.8
X$42745 25 2114 2152 2086 2178 44 AOI21_X4
* cell instance $42746 r0 *1 413.44,79.8
X$42746 1848 2068 25 44 2178 NOR2_X1
* cell instance $42749 r0 *1 415.91,79.8
X$42749 2112 2193 639 44 25 2156 OAI21_X2
* cell instance $42750 r0 *1 417.24,79.8
X$42750 2021 1999 2134 2154 2153 1909 44 25 AOI221_X2
* cell instance $42751 r0 *1 419.33,79.8
X$42751 2154 2153 2137 1999 2021 2158 44 25 AOI221_X2
* cell instance $42754 r0 *1 421.99,79.8
X$42754 2194 1501 25 44 2176 NAND2_X1
* cell instance $42756 r0 *1 422.75,79.8
X$42756 2155 2156 1501 25 44 2161 NAND3_X1
* cell instance $42759 r0 *1 426.74,79.8
X$42759 2176 2157 2197 25 2115 44 AOI21_X1
* cell instance $42760 r0 *1 427.5,79.8
X$42760 2197 2157 25 44 2159 NAND2_X1
* cell instance $42761 m0 *1 427.88,79.8
X$42761 2115 1081 2116 44 25 2160 OAI21_X2
* cell instance $42763 m0 *1 429.21,79.8
X$42763 2161 2116 2159 1081 25 44 2199 NOR4_X1
* cell instance $42766 m0 *1 434.72,79.8
X$42766 2044 2128 44 25 1580 AND2_X1
* cell instance $42769 r0 *1 428.07,79.8
X$42769 2158 1083 25 44 2174 NAND2_X1
* cell instance $42770 r0 *1 428.64,79.8
X$42770 1081 2159 2116 2161 44 2173 25 OR4_X2
* cell instance $42771 r0 *1 429.97,79.8
X$42771 2159 2174 44 25 2162 XNOR2_X1
* cell instance $42772 r0 *1 431.11,79.8
X$42772 2043 1081 2160 2173 2430 44 25 AOI211_X2
* cell instance $42776 r0 *1 436.43,79.8
X$42776 2043 1976 1081 25 44 2212 NOR3_X1
* cell instance $42777 r0 *1 437.19,79.8
X$42777 2162 2212 25 44 2163 NAND2_X1
* cell instance $42779 r0 *1 437.95,79.8
X$42779 551 2163 2201 2170 2164 2210 25 44 OAI221_X2
* cell instance $42780 m0 *1 439.09,79.8
X$42780 1333 1168 2209 25 44 1937 OR3_X2
* cell instance $42785 m0 *1 447.26,79.8
X$42785 2127 2124 25 44 2128 XOR2_X1
* cell instance $42786 m0 *1 448.4,79.8
X$42786 2127 2122 1857 44 25 2026 OAI21_X2
* cell instance $42788 m0 *1 450.49,79.8
X$42788 1482 1529 1978 2118 2079 2124 44 25 AOI221_X2
* cell instance $42794 r0 *1 447.07,79.8
X$42794 2207 2203 44 25 2127 AND2_X1
* cell instance $42795 r0 *1 447.83,79.8
X$42795 1539 2235 2233 44 25 1861 OAI21_X2
* cell instance $42798 r0 *1 452.96,79.8
X$42798 2167 2168 44 1985 25 XOR2_X2
* cell instance $42799 m0 *1 454.67,79.8
X$42799 2080 1777 44 25 2122 AND2_X1
* cell instance $42802 r0 *1 454.67,79.8
X$42802 2168 2167 25 44 1449 XNOR2_X2
* cell instance $42803 m0 *1 456,79.8
X$42803 1777 1482 2121 25 2117 44 AOI21_X1
* cell instance $42805 m0 *1 456.76,79.8
X$42805 1857 25 44 2118 INV_X1
* cell instance $42806 m0 *1 457.14,79.8
X$42806 1941 1528 2118 44 2121 25 OAI21_X1
* cell instance $42812 r0 *1 458.66,79.8
X$42812 2165 1490 1777 25 2166 44 AOI21_X1
* cell instance $42814 m0 *1 459.04,79.8
X$42814 2118 2166 1528 44 25 2081 OAI21_X2
* cell instance $42863 r0 *1 459.42,79.8
X$42863 1941 25 44 2165 INV_X1
* cell instance $43100 m0 *1 349.22,82.6
X$43100 1740 2090 1667 44 25 2179 OAI21_X2
* cell instance $43101 m0 *1 350.55,82.6
X$43101 1740 2005 25 44 2236 NAND2_X1
* cell instance $43102 m0 *1 351.12,82.6
X$43102 2090 2119 2236 25 2237 44 AOI21_X1
* cell instance $43104 m0 *1 352.07,82.6
X$43104 25 2211 2179 2050 2238 44 NOR3_X4
* cell instance $43105 m0 *1 354.73,82.6
X$43105 2050 2179 1959 25 44 2180 NOR3_X1
* cell instance $43127 r0 *1 350.17,82.6
X$43127 25 2142 1669 2006 2005 44 AOI21_X4
* cell instance $43129 r0 *1 352.83,82.6
X$43129 2143 2142 1959 25 44 2221 NAND3_X2
* cell instance $43131 r0 *1 354.35,82.6
X$43131 2211 2050 2179 44 25 2181 OAI21_X2
* cell instance $43133 r0 *1 355.87,82.6
X$43133 1899 2240 25 44 2249 NOR2_X2
* cell instance $43134 m0 *1 356.06,82.6
X$43134 2180 877 2003 25 44 2240 NOR3_X1
* cell instance $43137 m0 *1 357.01,82.6
X$43137 2003 877 2180 25 44 2186 OR3_X2
* cell instance $43140 r0 *1 358.34,82.6
X$43140 2181 2144 1801 2221 2356 25 44 OAI211_X2
* cell instance $43141 m0 *1 358.72,82.6
X$43141 2181 1801 2221 44 25 2213 OAI21_X2
* cell instance $43145 m0 *1 364.61,82.6
X$43145 2095 2213 2096 44 2184 25 OAI21_X1
* cell instance $43155 r0 *1 362.9,82.6
X$43155 2222 2223 2101 44 25 2262 OAI21_X2
* cell instance $43159 r0 *1 365.56,82.6
X$43159 2172 2244 2243 44 2263 25 OAI21_X1
* cell instance $43161 r0 *1 366.51,82.6
X$43161 1907 1512 25 44 2243 NOR2_X1
* cell instance $43164 r0 *1 367.65,82.6
X$43164 1728 1799 1411 44 2244 25 OAI21_X1
* cell instance $43167 r0 *1 368.98,82.6
X$43167 1799 1728 25 44 2287 OR2_X1
* cell instance $43169 r0 *1 370.5,82.6
X$43169 2010 1879 2147 25 44 2266 OR3_X2
* cell instance $43170 r0 *1 371.64,82.6
X$43170 2010 2147 877 44 25 2326 OAI21_X2
* cell instance $43175 r0 *1 378.67,82.6
X$43175 2101 2103 25 44 2290 NOR2_X1
* cell instance $43177 m0 *1 381.14,82.6
X$43177 2267 2186 25 44 2057 NAND2_X2
* cell instance $43178 m0 *1 379.43,82.6
X$43178 1802 1360 2096 25 44 NOR2_X4
* cell instance $43183 r0 *1 379.81,82.6
X$43183 1737 2268 1907 44 2251 25 NOR3_X2
* cell instance $43189 m0 *1 389.31,82.6
X$43189 1416 2216 2012 25 2217 44 AOI21_X1
* cell instance $43191 r0 *1 389.31,82.6
X$43191 2216 764 25 44 2254 NOR2_X1
* cell instance $43192 r0 *1 389.88,82.6
X$43192 2012 2254 25 44 2220 XNOR2_X2
* cell instance $43194 m0 *1 391.21,82.6
X$43194 2048 44 2065 25 BUF_X4
* cell instance $43195 m0 *1 393.3,82.6
X$43195 2217 2062 1831 25 44 2271 NAND3_X1
* cell instance $43197 m0 *1 394.25,82.6
X$43197 1831 2062 2217 44 25 2187 AND3_X1
* cell instance $43201 m0 *1 397.67,82.6
X$43201 2219 25 44 2257 INV_X1
* cell instance $43204 m0 *1 399,82.6
X$43204 25 1885 2135 1461 2219 2190 44 NAND4_X4
* cell instance $43210 r0 *1 395.39,82.6
X$43210 2064 2063 2059 44 2295 25 OAI21_X1
* cell instance $43212 r0 *1 396.53,82.6
X$43212 2295 2188 1426 25 44 2224 NOR3_X1
* cell instance $43213 r0 *1 397.29,82.6
X$43213 2348 2257 2224 2255 2188 2225 44 25 AOI221_X2
* cell instance $43216 r0 *1 402.61,82.6
X$43216 2220 2272 2225 44 25 2258 AND3_X1
* cell instance $43217 r0 *1 403.56,82.6
X$43217 2258 44 2333 25 BUF_X4
* cell instance $43218 m0 *1 406.22,82.6
X$43218 2190 2220 44 2112 25 XOR2_X2
* cell instance $43219 m0 *1 404.32,82.6
X$43219 2220 2190 25 44 2194 XNOR2_X2
* cell instance $43224 r0 *1 406.03,82.6
X$43224 2225 2226 1461 25 44 2193 NAND3_X2
* cell instance $43228 r0 *1 408.69,82.6
X$43228 1415 44 2229 25 BUF_X4
* cell instance $43229 m0 *1 410.02,82.6
X$43229 2087 2191 1848 2018 44 25 2152 OAI22_X2
* cell instance $43232 r0 *1 410.02,82.6
X$43232 2256 1860 25 44 2227 NAND2_X1
* cell instance $43235 m0 *1 412.11,82.6
X$43235 744 2186 2192 25 2247 44 AOI21_X1
* cell instance $43236 m0 *1 415.91,82.6
X$43236 2193 639 2112 25 44 2253 NOR3_X1
* cell instance $43238 m0 *1 416.86,82.6
X$43238 2193 25 44 2218 INV_X1
* cell instance $43239 m0 *1 417.24,82.6
X$43239 2218 1951 2194 25 44 2155 NAND3_X2
* cell instance $43240 m0 *1 418.57,82.6
X$43240 2194 2218 1951 25 2196 44 AOI21_X1
* cell instance $43243 r0 *1 412.11,82.6
X$43243 2228 2227 2067 44 2192 25 OAI21_X1
* cell instance $43244 r0 *1 412.87,82.6
X$43244 2227 2228 25 44 2250 NOR2_X1
* cell instance $43247 r0 *1 415.15,82.6
X$43247 2311 2291 2134 44 25 2157 OAI21_X4
* cell instance $43249 r0 *1 418.38,82.6
X$43249 2253 2196 2229 44 2315 25 OAI21_X1
* cell instance $43251 r0 *1 419.52,82.6
X$43251 2252 2230 1860 25 44 2200 NAND3_X1
* cell instance $43252 r0 *1 420.28,82.6
X$43252 2332 2250 25 44 2022 NOR2_X2
* cell instance $43253 r0 *1 421.23,82.6
X$43253 2230 2248 2044 2247 44 25 1825 AND4_X1
* cell instance $43255 r0 *1 422.56,82.6
X$43255 2155 2156 2229 25 44 2288 NAND3_X2
* cell instance $43256 m0 *1 422.94,82.6
X$43256 2155 2156 25 44 2246 NAND2_X1
* cell instance $43263 r0 *1 425.03,82.6
X$43263 2246 2330 25 44 2232 XNOR2_X2
* cell instance $43265 m0 *1 426.17,82.6
X$43265 2197 2157 2176 2158 1083 2214 44 25 AOI221_X2
* cell instance $43266 m0 *1 428.45,82.6
X$43266 1083 1892 2214 2199 2198 25 44 OAI211_X2
* cell instance $43267 m0 *1 430.16,82.6
X$43267 2160 2173 25 44 2215 NAND2_X2
* cell instance $43273 r0 *1 434.15,82.6
X$43273 2077 2245 44 25 2231 XNOR2_X1
* cell instance $43274 m0 *1 434.72,82.6
X$43274 2231 2200 25 44 1992 NOR2_X1
* cell instance $43277 m0 *1 436.05,82.6
X$43277 2200 2131 25 44 2206 NOR2_X1
* cell instance $43278 m0 *1 436.62,82.6
X$43278 2353 2162 25 44 2201 OR2_X1
* cell instance $43280 m0 *1 437.57,82.6
X$43280 2212 2162 25 44 2164 OR2_X1
* cell instance $43281 m0 *1 438.33,82.6
X$43281 2170 2201 2164 44 2209 25 OAI21_X1
* cell instance $43283 m0 *1 439.28,82.6
X$43283 2210 44 1775 25 BUF_X4
* cell instance $43289 r0 *1 439.47,82.6
X$43289 2232 2242 25 44 2168 XNOR2_X2
* cell instance $43292 r0 *1 443.08,82.6
X$43292 2232 1190 25 44 2279 NAND2_X2
* cell instance $43294 m0 *1 444.22,82.6
X$43294 2208 2202 25 44 2076 NAND2_X1
* cell instance $43296 m0 *1 444.79,82.6
X$43296 2202 2208 44 25 2077 AND2_X2
* cell instance $43299 r0 *1 444.79,82.6
X$43299 2241 2280 2239 44 25 1673 OAI21_X2
* cell instance $43300 r0 *1 446.12,82.6
X$43300 2233 2319 25 44 2241 NOR2_X1
* cell instance $43302 m0 *1 447.07,82.6
X$43302 2206 2203 2207 25 44 2078 NAND3_X2
* cell instance $43306 r0 *1 447.07,82.6
X$43306 2319 2233 2239 44 2203 25 OAI21_X1
* cell instance $43308 m0 *1 450.49,82.6
X$43308 1775 1863 1333 44 2204 25 NOR3_X2
* cell instance $43312 m0 *1 452.77,82.6
X$43312 2168 2204 44 25 2205 XNOR2_X1
* cell instance $43313 m0 *1 453.91,82.6
X$43313 2204 2233 2235 44 25 2167 OAI21_X2
* cell instance $43365 r0 *1 453.34,82.6
X$43365 2282 552 2229 2205 44 2234 25 NOR4_X2
* cell instance $43366 r0 *1 455.05,82.6
X$43366 2234 2168 2283 25 2079 44 AOI21_X2
* cell instance $43605 m0 *1 350.17,91
X$43605 2370 2141 1667 25 44 2456 NAND3_X1
* cell instance $43628 r0 *1 349.79,91
X$43628 1740 2090 25 44 2455 NAND2_X1
* cell instance $43629 r0 *1 350.36,91
X$43629 2455 1759 2456 25 44 2514 MUX2_X1
* cell instance $43632 r0 *1 352.26,91
X$43632 1740 2371 25 44 2478 XNOR2_X2
* cell instance $43633 m0 *1 353.02,91
X$43633 2141 1667 25 44 2457 NAND2_X1
* cell instance $43635 m0 *1 353.59,91
X$43635 1669 2371 44 25 2439 XNOR2_X1
* cell instance $43638 m0 *1 359.29,91
X$43638 2144 2338 2337 44 25 2489 OAI21_X4
* cell instance $43639 m0 *1 361.76,91
X$43639 25 1581 1876 2144 2145 2461 44 NOR4_X4
* cell instance $43642 m0 *1 367.46,91
X$43642 2439 2443 2372 2444 2545 44 25 AOI211_X2
* cell instance $43643 m0 *1 369.17,91
X$43643 25 2416 2443 2444 2372 44 AOI21_X4
* cell instance $43647 r0 *1 358.72,91
X$43647 2183 2460 2459 44 25 2448 OAI21_X2
* cell instance $43648 r0 *1 360.05,91
X$43648 2487 2461 2264 25 44 2460 NOR3_X1
* cell instance $43652 r0 *1 361.38,91
X$43652 2222 2264 2462 25 44 NOR2_X4
* cell instance $43654 r0 *1 363.85,91
X$43654 2264 2358 44 25 2479 AND2_X1
* cell instance $43658 r0 *1 365.94,91
X$43658 2489 2479 44 25 2463 AND2_X1
* cell instance $43659 r0 *1 366.7,91
X$43659 2103 44 1842 25 BUF_X4
* cell instance $43661 r0 *1 368.41,91
X$43661 2517 2342 2265 44 25 2444 OAI21_X2
* cell instance $43663 m0 *1 372.21,91
X$43663 25 1686 2415 2463 2403 2416 44 OAI211_X4
* cell instance $43670 r0 *1 373.54,91
X$43670 2416 2463 25 44 2493 NOR2_X2
* cell instance $43673 r0 *1 377.72,91
X$43673 2464 2343 2496 2497 2483 44 25 AOI211_X2
* cell instance $43676 m0 *1 381.33,91
X$43676 25 2403 2404 2345 2346 2305 44 OAI22_X4
* cell instance $43678 m0 *1 384.56,91
X$43678 2448 2417 44 25 2305 AND2_X2
* cell instance $43679 m0 *1 385.51,91
X$43679 2329 2448 2417 25 2375 44 AOI21_X1
* cell instance $43682 m0 *1 387.22,91
X$43682 2377 2418 2329 25 44 2419 OR3_X1
* cell instance $43683 m0 *1 388.17,91
X$43683 2329 2418 2377 25 44 2465 NOR3_X1
* cell instance $43684 m0 *1 388.93,91
X$43684 2306 2465 1364 44 2449 25 OAI21_X1
* cell instance $43687 r0 *1 381.14,91
X$43687 2464 2269 25 44 2404 OR2_X2
* cell instance $43688 r0 *1 382.09,91
X$43688 2417 2448 25 44 2406 NAND2_X2
* cell instance $43690 r0 *1 383.42,91
X$43690 25 2483 2524 2048 2374 2406 44 AOI22_X4
* cell instance $43691 r0 *1 386.65,91
X$43691 25 2418 2377 2345 2064 2305 44 OAI22_X4
* cell instance $43693 m0 *1 391.59,91
X$43693 2449 2412 2421 2420 2592 44 25 AOI211_X2
* cell instance $43694 m0 *1 390.83,91
X$43694 2412 2419 2411 25 2484 44 AOI21_X1
* cell instance $43695 m0 *1 393.3,91
X$43695 2421 2420 25 44 2466 NAND2_X1
* cell instance $43699 m0 *1 397.86,91
X$43699 2422 2423 2369 44 25 2450 OAI21_X2
* cell instance $43700 m0 *1 399.19,91
X$43700 25 2501 2380 2451 2450 44 AOI21_X4
* cell instance $43702 r0 *1 392.92,91
X$43702 2484 2466 25 44 2498 NAND2_X1
* cell instance $43705 r0 *1 394.06,91
X$43705 2307 2466 2484 44 25 2499 AND3_X2
* cell instance $43709 r0 *1 398.81,91
X$43709 2423 2499 25 44 2310 XNOR2_X2
* cell instance $43712 m0 *1 402.04,91
X$43712 1626 2349 2381 44 25 2467 AND3_X1
* cell instance $43713 m0 *1 403.75,91
X$43713 2381 2349 1626 25 44 2424 NAND3_X2
* cell instance $43714 m0 *1 405.08,91
X$43714 2424 2273 2310 44 2425 25 OAI21_X1
* cell instance $43718 r0 *1 405.27,91
X$43718 2333 2500 2486 2467 25 2454 44 NAND4_X2
* cell instance $43721 m0 *1 406.98,91
X$43721 2425 2454 2382 44 25 2468 AND3_X1
* cell instance $43722 m0 *1 408.12,91
X$43722 2382 2454 2425 25 44 2427 NAND3_X2
* cell instance $43726 r0 *1 408.69,91
X$43726 2500 2486 25 44 2383 NOR2_X1
* cell instance $43729 r0 *1 410.4,91
X$43729 2087 2191 25 44 2520 OR2_X1
* cell instance $43731 m0 *1 411.54,91
X$43731 2468 2426 25 2385 44 NAND2_X4
* cell instance $43733 m0 *1 413.25,91
X$43733 2427 2384 2386 25 44 NOR2_X4
* cell instance $43734 m0 *1 414.96,91
X$43734 2426 2468 2410 639 2453 25 44 OAI211_X2
* cell instance $43736 m0 *1 420.28,91
X$43736 2452 2387 2073 2047 2379 2431 25 44 OAI221_X2
* cell instance $43737 m0 *1 417.05,91
X$43737 25 2385 2195 2351 2428 2312 44 OAI211_X4
* cell instance $43740 m0 *1 424.08,91
X$43740 2386 729 2359 44 25 2446 OAI21_X2
* cell instance $43741 m0 *1 425.41,91
X$43741 2402 2428 1932 1364 25 44 2445 NAND4_X1
* cell instance $43743 m0 *1 426.55,91
X$43743 2385 729 2379 25 44 2447 NAND3_X1
* cell instance $43745 m0 *1 427.5,91
X$43745 2385 1932 2388 25 2389 44 AOI21_X2
* cell instance $43747 m0 *1 429.02,91
X$43747 2198 1976 2447 2445 2442 44 25 AOI211_X2
* cell instance $43750 m0 *1 431.68,91
X$43750 2430 2432 2431 2399 25 44 2471 AOI22_X2
* cell instance $43752 m0 *1 433.58,91
X$43752 1416 2430 2432 25 2469 44 AOI21_X1
* cell instance $43753 m0 *1 434.34,91
X$43753 2433 2469 1893 25 2482 44 AOI21_X1
* cell instance $43755 m0 *1 435.86,91
X$43755 2433 2481 2482 25 44 2440 MUX2_X1
* cell instance $43759 r0 *1 423.32,91
X$43759 2385 1932 2379 44 2485 25 NOR3_X2
* cell instance $43760 r0 *1 424.65,91
X$43760 25 2519 2485 2083 2534 2314 44 OAI22_X4
* cell instance $43761 r0 *1 427.88,91
X$43761 2388 2385 1932 25 44 2535 NAND3_X2
* cell instance $43762 r0 *1 429.21,91
X$43762 2385 1168 25 44 2503 NOR2_X1
* cell instance $43767 r0 *1 435.29,91
X$43767 2433 25 44 2505 INV_X1
* cell instance $43769 r0 *1 435.86,91
X$43769 2505 2481 25 44 2437 XNOR2_X2
* cell instance $43772 r0 *1 438.9,91
X$43772 2507 2229 25 44 2470 NAND2_X1
* cell instance $43773 m0 *1 439.85,91
X$43773 2471 2442 25 44 2472 OR2_X1
* cell instance $43774 m0 *1 439.09,91
X$43774 2442 2471 2229 44 2480 25 OAI21_X1
* cell instance $43778 m0 *1 445.93,91
X$43778 2440 2441 2235 2474 25 44 2397 NAND4_X1
* cell instance $43780 m0 *1 447.07,91
X$43780 2434 2391 25 44 2354 NAND2_X1
* cell instance $43781 m0 *1 447.64,91
X$43781 25 2434 2391 2233 2435 2229 44 AOI22_X4
* cell instance $43782 m0 *1 450.87,91
X$43782 2229 2281 2435 44 2436 25 OAI21_X1
* cell instance $43783 m0 *1 451.63,91
X$43783 2436 1898 25 44 2438 NAND2_X1
* cell instance $43784 m0 *1 452.2,91
X$43784 2437 2235 25 44 2476 NOR2_X1
* cell instance $43786 r0 *1 439.47,91
X$43786 2470 2480 2538 44 25 2473 MUX2_X2
* cell instance $43787 r0 *1 441.18,91
X$43787 2507 2472 1893 44 25 2435 MUX2_X2
* cell instance $43791 r0 *1 446.88,91
X$43791 2392 2508 25 44 1898 NAND2_X2
* cell instance $43792 r0 *1 447.83,91
X$43792 2473 2474 2392 25 44 2475 OR3_X1
* cell instance $43793 r0 *1 448.78,91
X$43793 2437 2392 2508 2512 25 44 2393 NAND4_X1
* cell instance $43794 r0 *1 449.73,91
X$43794 2473 2512 2395 44 25 2513 AND3_X1
* cell instance $43797 r0 *1 452.58,91
X$43797 2476 2473 25 44 2477 NOR2_X1
* cell instance $43799 m0 *1 453.15,91
X$43799 2474 2438 25 44 2030 XNOR2_X2
* cell instance $43848 r0 *1 453.15,91
X$43848 1898 25 44 552 INV_X2
* cell instance $44087 m0 *1 353.97,96.6
X$44087 2090 2457 1759 25 2553 44 AOI21_X2
* cell instance $44088 m0 *1 355.3,96.6
X$44088 2090 1759 2457 44 25 2573 AND3_X1
* cell instance $44092 m0 *1 360.24,96.6
X$44092 2553 2573 2462 2458 2265 2554 25 44 OAI221_X2
* cell instance $44093 m0 *1 362.33,96.6
X$44093 2554 2414 25 44 2577 NOR2_X1
* cell instance $44096 m0 *1 365.18,96.6
X$44096 2401 2146 25 44 2613 NOR2_X1
* cell instance $44120 r0 *1 360.24,96.6
X$44120 2146 2553 2573 25 44 2584 NOR3_X1
* cell instance $44122 r0 *1 361.19,96.6
X$44122 2458 2462 2584 44 2611 25 OAI21_X1
* cell instance $44123 r0 *1 361.95,96.6
X$44123 2554 2611 2414 44 25 2464 MUX2_X2
* cell instance $44124 r0 *1 363.66,96.6
X$44124 25 2612 2613 2543 2615 2666 44 NOR4_X4
* cell instance $44125 r0 *1 367.08,96.6
X$44125 2342 2265 763 44 2612 25 NOR3_X2
* cell instance $44126 m0 *1 367.84,96.6
X$44126 25 2517 2265 2342 2521 44 NOR3_X4
* cell instance $44128 m0 *1 370.5,96.6
X$44128 2268 1512 25 44 2491 NOR2_X2
* cell instance $44131 r0 *1 369.17,96.6
X$44131 2265 2585 25 44 2586 XNOR2_X2
* cell instance $44132 r0 *1 371.07,96.6
X$44132 2342 2268 25 44 2585 NOR2_X2
* cell instance $44133 m0 *1 372.02,96.6
X$44133 2578 2545 2576 2577 2415 2418 25 44 OAI221_X2
* cell instance $44138 r0 *1 373.54,96.6
X$44138 25 2586 2415 2545 2374 2578 44 OAI22_X4
* cell instance $44139 m0 *1 375.44,96.6
X$44139 1907 2545 2578 44 25 2555 OAI21_X2
* cell instance $44143 r0 *1 376.77,96.6
X$44143 2522 2492 25 44 2682 NAND2_X1
* cell instance $44146 r0 *1 378.48,96.6
X$44146 2555 2587 2556 25 44 2670 NAND3_X2
* cell instance $44147 m0 *1 378.86,96.6
X$44147 2555 2523 2548 25 44 2045 AND3_X4
* cell instance $44149 m0 *1 380.95,96.6
X$44149 2523 2548 2374 2406 25 44 2581 AOI22_X2
* cell instance $44153 r0 *1 380.95,96.6
X$44153 2149 25 44 2589 BUF_X2
* cell instance $44155 r0 *1 382.47,96.6
X$44155 25 2017 2347 2556 2587 44 AOI21_X4
* cell instance $44156 m0 *1 383.23,96.6
X$44156 2524 2525 2581 2302 2591 44 25 AOI211_X2
* cell instance $44159 m0 *1 385.7,96.6
X$44159 2149 2374 2406 25 44 2557 NAND3_X1
* cell instance $44164 r0 *1 384.94,96.6
X$44164 2149 2587 2556 25 44 2590 NAND3_X1
* cell instance $44166 r0 *1 386.08,96.6
X$44166 2557 2590 2525 25 44 2649 NAND3_X2
* cell instance $44167 r0 *1 387.41,96.6
X$44167 2525 2590 2557 44 25 2623 AND3_X2
* cell instance $44170 m0 *1 392.35,96.6
X$44170 2559 2498 2593 2617 44 2558 25 NOR4_X2
* cell instance $44174 m0 *1 395.01,96.6
X$44174 2015 1364 25 44 2559 NAND2_X1
* cell instance $44175 m0 *1 395.58,96.6
X$44175 2559 2499 2526 25 44 2599 MUX2_X1
* cell instance $44178 m0 *1 397.86,96.6
X$44178 2089 44 2423 25 BUF_X4
* cell instance $44179 m0 *1 399.19,96.6
X$44179 2423 2379 25 44 2560 NOR2_X1
* cell instance $44180 m0 *1 399.76,96.6
X$44180 2560 2550 2499 44 25 2561 MUX2_X2
* cell instance $44183 m0 *1 402.42,96.6
X$44183 25 2561 2583 2273 2087 2424 44 OAI211_X4
* cell instance $44184 m0 *1 405.65,96.6
X$44184 25 2486 2600 2501 2308 2601 44 NOR4_X4
* cell instance $44190 r0 *1 392.92,96.6
X$44190 2422 2616 25 44 2617 NAND2_X1
* cell instance $44192 r0 *1 395.01,96.6
X$44192 2423 1907 25 44 2595 NOR2_X2
* cell instance $44195 r0 *1 397.1,96.6
X$44195 2369 2089 2348 2594 44 2596 25 NOR4_X2
* cell instance $44196 r0 *1 398.81,96.6
X$44196 2596 2625 2598 25 44 2619 NOR3_X1
* cell instance $44198 r0 *1 399.76,96.6
X$44198 2598 2625 2596 25 44 2583 OR3_X2
* cell instance $44201 r0 *1 401.47,96.6
X$44201 2619 2599 2333 2467 2626 44 25 AOI211_X2
* cell instance $44204 r0 *1 406.6,96.6
X$44204 2600 44 2068 25 BUF_X4
* cell instance $44207 m0 *1 413.25,96.6
X$44207 2558 2045 25 44 2252 NOR2_X1
* cell instance $44213 r0 *1 415.72,96.6
X$44213 2620 2379 2602 2601 2531 44 25 AOI211_X2
* cell instance $44214 r0 *1 417.43,96.6
X$44214 2601 2602 25 44 2230 NAND2_X2
* cell instance $44217 r0 *1 419.33,96.6
X$44217 2532 2603 25 44 2533 NOR2_X1
* cell instance $44218 m0 *1 419.71,96.6
X$44218 2153 2387 2532 44 25 2618 AND3_X1
* cell instance $44221 m0 *1 422.18,96.6
X$44221 2562 2230 2313 2277 44 25 2245 AND4_X1
* cell instance $44225 r0 *1 420.09,96.6
X$44225 2533 2618 2604 44 2313 25 OAI21_X1
* cell instance $44227 r0 *1 421.04,96.6
X$44227 2252 2230 2562 25 44 2716 NAND3_X1
* cell instance $44228 r0 *1 421.8,96.6
X$44228 2562 2230 2252 2313 44 25 2317 AND4_X1
* cell instance $44231 m0 *1 424.46,96.6
X$44231 2387 2563 44 25 2580 XNOR2_X1
* cell instance $44233 r0 *1 425.98,96.6
X$44233 2564 2502 2580 44 25 2605 OAI21_X2
* cell instance $44235 m0 *1 426.74,96.6
X$44235 2502 2580 25 44 2579 OR2_X1
* cell instance $44236 m0 *1 428.26,96.6
X$44236 2429 2433 2534 2565 2575 25 44 OAI211_X2
* cell instance $44238 m0 *1 431.49,96.6
X$44238 25 2606 2504 2537 2536 2564 2579 44 AOI221_X4
* cell instance $44242 r0 *1 427.31,96.6
X$44242 25 2605 2429 2534 2631 2565 44 OAI211_X4
* cell instance $44245 r0 *1 437.38,96.6
X$44245 2606 2568 44 25 2614 AND2_X1
* cell instance $44246 r0 *1 438.14,96.6
X$44246 2614 2610 2566 2353 2170 2607 25 44 2434 OAI33_X1
* cell instance $44247 m0 *1 438.9,96.6
X$44247 2547 2567 25 44 2568 NOR2_X1
* cell instance $44248 m0 *1 438.14,96.6
X$44248 2567 2547 44 25 2566 AND2_X1
* cell instance $44251 r0 *1 439.47,96.6
X$44251 2606 2568 2575 2608 25 44 2609 AOI22_X1
* cell instance $44252 r0 *1 440.42,96.6
X$44252 2575 2608 44 25 2610 AND2_X1
* cell instance $44253 m0 *1 441.18,96.6
X$44253 551 2609 2574 25 2572 44 AOI21_X1
* cell instance $44254 m0 *1 440.61,96.6
X$44254 2547 2567 25 44 2574 NAND2_X1
* cell instance $44255 m0 *1 441.94,96.6
X$44255 2547 2539 25 44 2571 NOR2_X2
* cell instance $44259 m0 *1 443.27,96.6
X$44259 2544 2567 25 44 2569 NAND2_X1
* cell instance $44261 m0 *1 445.93,96.6
X$44261 2570 1893 25 44 2541 NOR2_X1
* cell instance $44263 m0 *1 446.5,96.6
X$44263 1893 2570 25 44 2391 OR2_X2
* cell instance $44552 m0 *1 359.86,102.2
X$44552 2640 2458 2414 2487 2665 2417 25 44 OAI221_X2
* cell instance $44553 m0 *1 361.95,102.2
X$44553 2487 2268 25 44 2665 NAND2_X1
* cell instance $44556 m0 *1 363.47,102.2
X$44556 2641 2462 25 44 2680 OR2_X1
* cell instance $44584 r0 *1 363.09,102.2
X$44584 2462 2641 2679 25 44 NOR2_X4
* cell instance $44586 m0 *1 365.56,102.2
X$44586 2705 2448 25 44 2706 NAND2_X1
* cell instance $44589 m0 *1 366.32,102.2
X$44589 2622 2490 2642 2325 2643 2725 25 44 OAI221_X2
* cell instance $44590 m0 *1 368.41,102.2
X$44590 2144 1512 25 44 2707 NOR2_X1
* cell instance $44595 r0 *1 367.65,102.2
X$44595 2643 2707 2679 2708 25 44 2726 AOI22_X1
* cell instance $44597 m0 *1 369.93,102.2
X$44597 1581 2268 25 44 2728 XNOR2_X2
* cell instance $44598 m0 *1 369.36,102.2
X$44598 1842 1581 25 44 2708 NOR2_X1
* cell instance $44599 m0 *1 371.83,102.2
X$44599 1512 2268 25 44 2683 XNOR2_X2
* cell instance $44600 m0 *1 373.73,102.2
X$44600 2679 2682 2645 2709 2668 2727 25 44 OAI221_X2
* cell instance $44602 m0 *1 376.58,102.2
X$44602 2495 2343 2588 44 25 2681 OAI21_X2
* cell instance $44604 m0 *1 378.67,102.2
X$44604 25 2343 2495 2588 2683 2711 44 NOR4_X4
* cell instance $44606 r0 *1 369.36,102.2
X$44606 2517 2644 25 44 2767 XNOR2_X2
* cell instance $44607 r0 *1 371.26,102.2
X$44607 2495 2680 25 44 2709 NAND2_X1
* cell instance $44608 r0 *1 371.83,102.2
X$44608 2668 2679 25 44 2741 NOR2_X1
* cell instance $44610 r0 *1 372.59,102.2
X$44610 2706 2741 2749 2493 2750 25 44 OAI211_X2
* cell instance $44613 r0 *1 374.87,102.2
X$44613 2683 2493 2681 25 2819 44 NAND3_X4
* cell instance $44614 r0 *1 377.34,102.2
X$44614 2681 2682 25 44 2744 NAND2_X1
* cell instance $44616 r0 *1 378.1,102.2
X$44616 25 2749 2586 2415 2589 44 AOI21_X4
* cell instance $44617 r0 *1 380.57,102.2
X$44617 2589 2415 2728 2586 25 44 2684 AOI211_X4
* cell instance $44618 m0 *1 382.66,102.2
X$44618 2711 2684 2064 2063 44 25 2712 OAI22_X1
* cell instance $44620 m0 *1 383.61,102.2
X$44620 25 2714 2645 2065 2017 44 AOI21_X4
* cell instance $44621 m0 *1 386.08,102.2
X$44621 2683 2646 2647 44 25 2673 AND3_X1
* cell instance $44622 m0 *1 387.03,102.2
X$44622 2683 2647 2646 25 2718 44 AOI21_X1
* cell instance $44626 r0 *1 383.04,102.2
X$44626 2712 1884 2713 44 25 2616 OAI21_X2
* cell instance $44627 r0 *1 384.37,102.2
X$44627 2683 2586 25 44 2713 NAND2_X1
* cell instance $44628 r0 *1 384.94,102.2
X$44628 2744 2065 2017 25 2715 44 AOI21_X2
* cell instance $44630 r0 *1 386.46,102.2
X$44630 2495 2714 25 44 2692 XNOR2_X2
* cell instance $44631 r0 *1 388.36,102.2
X$44631 2683 764 2495 25 44 2717 NOR3_X1
* cell instance $44632 m0 *1 389.12,102.2
X$44632 2331 1885 2673 2718 2648 25 44 OAI211_X2
* cell instance $44634 m0 *1 390.83,102.2
X$44634 2648 2686 25 44 2653 NAND2_X2
* cell instance $44635 m0 *1 391.78,102.2
X$44635 2685 2549 2649 25 2687 44 AOI21_X1
* cell instance $44636 m0 *1 392.54,102.2
X$44636 2549 2649 25 2689 44 NAND2_X4
* cell instance $44639 r0 *1 389.31,102.2
X$44639 2717 2746 757 2685 44 25 2686 OAI22_X2
* cell instance $44641 r0 *1 391.21,102.2
X$44641 2686 2648 44 25 2639 AND2_X2
* cell instance $44643 r0 *1 392.54,102.2
X$44643 2687 2688 1885 2331 2720 44 25 AOI211_X2
* cell instance $44645 m0 *1 398.05,102.2
X$44645 25 2650 2624 2678 2722 2721 44 OAI22_X4
* cell instance $44646 m0 *1 394.63,102.2
X$44646 25 757 2423 2689 2369 2721 44 NOR4_X4
* cell instance $44650 r0 *1 395.96,102.2
X$44650 25 2624 2331 2592 2015 44 AOI21_X4
* cell instance $44652 r0 *1 399.19,102.2
X$44652 2688 2685 757 44 25 2678 OAI21_X2
* cell instance $44654 r0 *1 402.04,102.2
X$44654 2422 2561 2651 2729 2692 2655 25 44 OAI221_X2
* cell instance $44655 m0 *1 402.99,102.2
X$44655 2597 2333 2677 25 2690 44 AOI21_X2
* cell instance $44656 m0 *1 402.42,102.2
X$44656 1885 2685 25 44 2651 NOR2_X1
* cell instance $44658 m0 *1 405.84,102.2
X$44658 2151 2653 2654 44 2627 25 NOR3_X2
* cell instance $44660 m0 *1 407.36,102.2
X$44660 2693 2694 2087 2722 2674 1929 25 44 OAI221_X2
* cell instance $44661 m0 *1 409.45,102.2
X$44661 2656 25 44 2694 INV_X2
* cell instance $44662 m0 *1 410.02,102.2
X$44662 2639 2626 2654 2655 2724 2697 44 25 AOI221_X2
* cell instance $44663 m0 *1 412.11,102.2
X$44663 2626 2582 2551 2655 2656 2695 44 25 AOI221_X2
* cell instance $44665 m0 *1 414.39,102.2
X$44665 25 2530 2697 2696 2698 44 AOI21_X4
* cell instance $44667 m0 *1 419.9,102.2
X$44667 2021 2000 1999 44 25 2630 OAI21_X2
* cell instance $44671 m0 *1 425.98,102.2
X$44671 729 2379 2428 25 2659 44 AOI21_X2
* cell instance $44675 m0 *1 440.23,102.2
X$44675 2563 2659 25 44 2660 XOR2_X1
* cell instance $44676 m0 *1 441.37,102.2
X$44676 2563 2659 25 44 2635 XNOR2_X2
* cell instance $44677 m0 *1 443.27,102.2
X$44677 2635 2661 2539 25 44 2663 NAND3_X1
* cell instance $44685 r0 *1 404.13,102.2
X$44685 2652 2594 2273 44 2691 25 NOR3_X2
* cell instance $44688 r0 *1 406.6,102.2
X$44688 2674 2693 2694 44 25 2086 OAI21_X4
* cell instance $44689 r0 *1 409.07,102.2
X$44689 2087 2693 2694 44 25 2696 OAI21_X2
* cell instance $44692 r0 *1 410.97,102.2
X$44692 2639 2656 44 25 2724 AND2_X1
* cell instance $44693 r0 *1 411.73,102.2
X$44693 25 2413 2551 2655 2656 44 AOI21_X4
* cell instance $44696 r0 *1 414.77,102.2
X$44696 2696 2698 44 25 2723 AND2_X1
* cell instance $44698 r0 *1 415.72,102.2
X$44698 2723 2697 25 44 2699 OR2_X1
* cell instance $44703 r0 *1 419.33,102.2
X$44703 2000 1999 25 44 2532 NOR2_X2
* cell instance $44705 r0 *1 420.66,102.2
X$44705 2000 1999 2699 25 44 2719 NOR3_X1
* cell instance $44707 r0 *1 421.8,102.2
X$44707 2074 2428 2719 44 2700 25 OAI21_X1
* cell instance $44709 r0 *1 425.6,102.2
X$44709 2716 2700 2701 25 2704 44 AOI21_X2
* cell instance $44712 r0 *1 428.64,102.2
X$44712 2631 2658 2701 2700 25 44 2702 AOI22_X1
* cell instance $44714 r0 *1 429.78,102.2
X$44714 2503 2215 2605 2710 25 2740 44 NAND4_X2
* cell instance $44715 r0 *1 431.49,102.2
X$44715 2605 2215 2503 2710 44 25 2607 AND4_X1
* cell instance $44719 r0 *1 433.96,102.2
X$44719 1892 2539 2703 2606 2743 2506 25 44 OAI221_X2
* cell instance $44720 r0 *1 436.05,102.2
X$44720 1892 2661 2539 25 44 2743 NAND3_X1
* cell instance $45003 m0 *1 353.97,93.8
X$45003 25 2514 2260 2488 2461 2264 44 AOI22_X4
* cell instance $45028 m0 *1 360.05,93.8
X$45028 2488 44 2103 25 BUF_X4
* cell instance $45032 m0 *1 362.33,93.8
X$45032 2264 2358 2146 44 25 2516 AND3_X1
* cell instance $45037 r0 *1 361.38,93.8
X$45037 2488 25 44 2268 INV_X4
* cell instance $45040 m0 *1 363.66,93.8
X$45040 2103 2516 2489 25 2543 44 AOI21_X2
* cell instance $45043 r0 *1 364.42,93.8
X$45043 25 2479 2489 2615 2517 1581 44 AOI22_X4
* cell instance $45045 m0 *1 365.37,93.8
X$45045 2479 2489 25 44 2492 NAND2_X2
* cell instance $45046 m0 *1 366.51,93.8
X$45046 2185 2103 25 44 2490 NAND2_X1
* cell instance $45049 m0 *1 368.79,93.8
X$45049 25 2491 2478 2521 2496 2546 44 OAI211_X4
* cell instance $45052 m0 *1 375.82,93.8
X$45052 2459 2492 25 44 2497 OR2_X2
* cell instance $45053 m0 *1 376.77,93.8
X$45053 25 2495 2343 2345 2496 2497 44 AOI22_X4
* cell instance $45055 m0 *1 386.08,93.8
X$45055 2269 1907 2377 25 44 NOR2_X4
* cell instance $45061 r0 *1 367.65,93.8
X$45061 25 2546 2185 2401 2146 44 AOI21_X4
* cell instance $45063 r0 *1 370.88,93.8
X$45063 2491 2546 2521 44 25 2522 OAI21_X2
* cell instance $45066 r0 *1 372.78,93.8
X$45066 2492 2459 25 44 2578 NOR2_X2
* cell instance $45069 r0 *1 374.68,93.8
X$45069 2343 1678 2492 2522 2587 44 25 AOI211_X2
* cell instance $45070 r0 *1 376.39,93.8
X$45070 1678 2522 2492 25 2523 44 AOI21_X2
* cell instance $45073 r0 *1 378.67,93.8
X$45073 2269 2464 2343 44 2548 25 NOR3_X2
* cell instance $45074 r0 *1 380,93.8
X$45074 2269 2464 25 44 2556 NOR2_X2
* cell instance $45077 r0 *1 383.23,93.8
X$45077 1907 2269 25 44 2524 OR2_X2
* cell instance $45078 r0 *1 384.18,93.8
X$45078 2587 2556 25 44 2373 NAND2_X1
* cell instance $45079 r0 *1 384.75,93.8
X$45079 2494 25 44 2525 INV_X1
* cell instance $45083 r0 *1 387.79,93.8
X$45083 25 2494 2377 2346 2549 2347 44 OAI211_X4
* cell instance $45087 r0 *1 395.96,93.8
X$45087 2423 1364 25 44 2526 NAND2_X1
* cell instance $45091 r0 *1 399.19,93.8
X$45091 2015 2379 25 44 2550 NOR2_X1
* cell instance $45093 m0 *1 399.57,93.8
X$45093 2015 2499 25 44 2500 XNOR2_X2
* cell instance $45095 m0 *1 405.27,93.8
X$45095 1678 2500 2501 2273 44 2674 25 OR4_X2
* cell instance $45102 r0 *1 404.89,93.8
X$45102 25 1678 2500 2501 2273 2551 44 NOR4_X4
* cell instance $45103 m0 *1 410.97,93.8
X$45103 1848 2018 2552 2413 2520 2139 25 44 OAI221_X2
* cell instance $45104 m0 *1 407.74,93.8
X$45104 25 1848 2675 2413 2113 2528 44 OAI211_X4
* cell instance $45108 r0 *1 409.07,93.8
X$45108 2527 2529 1765 25 44 2528 NAND3_X2
* cell instance $45109 r0 *1 410.4,93.8
X$45109 2582 2527 2529 1886 25 2191 44 NAND4_X2
* cell instance $45110 r0 *1 412.11,93.8
X$45110 1886 2527 2529 25 44 2552 NAND3_X1
* cell instance $45114 r0 *1 417.62,93.8
X$45114 2530 2531 44 25 2154 AND2_X1
* cell instance $45115 r0 *1 418.38,93.8
X$45115 2531 2530 25 44 2084 NAND2_X1
* cell instance $45118 r0 *1 419.52,93.8
X$45118 2533 2530 25 44 2286 NAND2_X2
* cell instance $45119 m0 *1 419.71,93.8
X$45119 2532 2387 2153 25 44 2248 NAND3_X1
* cell instance $45125 m0 *1 422.37,93.8
X$45125 2379 2047 2073 44 25 2502 OAI21_X2
* cell instance $45127 m0 *1 425.03,93.8
X$45127 2502 2428 2402 25 2519 44 AOI21_X2
* cell instance $45131 m0 *1 430.16,93.8
X$45131 2328 2400 25 44 2504 OR2_X1
* cell instance $45134 m0 *1 435.48,93.8
X$45134 2446 2535 2433 44 25 2507 AND3_X1
* cell instance $45140 r0 *1 428.64,93.8
X$45140 2400 2328 25 44 2565 NOR2_X2
* cell instance $45142 r0 *1 429.97,93.8
X$45142 2400 2328 2535 2446 2536 44 25 AOI211_X2
* cell instance $45144 r0 *1 432.06,93.8
X$45144 2505 2536 2537 2504 2634 44 25 AOI211_X2
* cell instance $45148 r0 *1 435.1,93.8
X$45148 2563 2446 2535 2433 44 25 2547 AND4_X1
* cell instance $45151 r0 *1 438.14,93.8
X$45151 2539 25 44 2353 INV_X1
* cell instance $45155 m0 *1 440.04,93.8
X$45155 25 1893 2472 2278 2540 2518 44 AOI22_X4
* cell instance $45160 r0 *1 439.85,93.8
X$45160 2538 25 44 551 INV_X4
* cell instance $45161 r0 *1 440.8,93.8
X$45161 2507 2563 25 44 2544 NAND2_X1
* cell instance $45162 r0 *1 441.37,93.8
X$45162 2539 2507 44 25 2540 AND2_X1
* cell instance $45163 r0 *1 442.13,93.8
X$45163 25 551 2569 2571 2511 2567 44 OAI22_X4
* cell instance $45165 r0 *1 445.74,93.8
X$45165 2473 2572 2541 44 25 2508 OAI21_X2
* cell instance $45168 r0 *1 447.64,93.8
X$45168 2319 25 44 2509 INV_X1
* cell instance $45169 r0 *1 448.02,93.8
X$45169 2473 2511 2512 44 25 2542 AND3_X1
* cell instance $45170 m0 *1 450.87,93.8
X$45170 2513 2511 44 1941 25 XOR2_X2
* cell instance $45171 m0 *1 448.21,93.8
X$45171 25 1978 2509 2515 552 2510 2513 2511 44 OAI222_X4
* cell instance $45179 r0 *1 448.97,93.8
X$45179 2509 2542 2508 2318 44 25 2510 OAI22_X1
* cell instance $45180 r0 *1 449.92,93.8
X$45180 2508 2318 25 44 2515 OR2_X1
* cell instance $45527 r0 *1 347.89,77
X$45527 25 1752 2003 1983 2004 44 AOI21_X4
* cell instance $45528 m0 *1 351.31,77
X$45528 1639 1696 1919 1747 25 2141 44 NAND4_X2
* cell instance $45529 m0 *1 349.6,77
X$45529 1832 1670 2005 1919 2004 25 44 OAI211_X2
* cell instance $45530 m0 *1 353.02,77
X$45530 1740 2005 1782 25 44 2120 NOR3_X1
* cell instance $45531 m0 *1 353.78,77
X$45531 1696 1639 1747 1960 44 25 2050 AND4_X2
* cell instance $45534 r0 *1 350.36,77
X$45534 1670 1832 25 44 2090 NAND2_X2
* cell instance $45537 r0 *1 351.88,77
X$45537 25 1747 1960 1798 1639 2143 44 NAND4_X4
* cell instance $45539 r0 *1 356.82,77
X$45539 2051 2082 44 25 2091 AND2_X1
* cell instance $45540 r0 *1 357.58,77
X$45540 2082 2051 25 44 2123 NAND2_X1
* cell instance $45542 r0 *1 358.34,77
X$45542 1752 2007 25 44 2092 NOR2_X1
* cell instance $45544 m0 *1 358.53,77
X$45544 1752 2007 1819 25 44 2008 NOR3_X1
* cell instance $45546 m0 *1 362.52,77
X$45546 2007 1752 2039 25 44 2052 OR3_X2
* cell instance $45551 m0 *1 369.17,77
X$45551 2009 1784 25 44 2053 NOR2_X1
* cell instance $45553 m0 *1 370.5,77
X$45553 2096 1411 2042 2010 25 2011 44 NAND4_X2
* cell instance $45558 r0 *1 359.1,77
X$45558 1800 1752 25 44 2093 NAND2_X2
* cell instance $45564 r0 *1 362.14,77
X$45564 25 2007 1752 2039 2145 44 NOR3_X4
* cell instance $45568 r0 *1 367.46,77
X$45568 25 1752 1800 2009 2055 1784 44 OAI211_X4
* cell instance $45569 r0 *1 370.69,77
X$45569 2009 1784 1747 44 2126 25 OAI21_X1
* cell instance $45570 r0 *1 371.45,77
X$45570 2011 1801 2126 25 44 2129 MUX2_X1
* cell instance $45573 r0 *1 374.49,77
X$45573 1908 2055 1924 25 44 2099 MUX2_X1
* cell instance $45574 r0 *1 375.82,77
X$45574 1924 1879 25 44 2130 NOR2_X1
* cell instance $45576 r0 *1 376.58,77
X$45576 2099 2085 25 44 2100 OR2_X1
* cell instance $45579 m0 *1 380.19,77
X$45579 25 1839 2045 2057 2025 44 NOR3_X4
* cell instance $45580 m0 *1 384.37,77
X$45580 1966 1967 25 44 2012 XNOR2_X2
* cell instance $45581 m0 *1 386.27,77
X$45581 1965 763 1968 44 25 2013 OAI21_X2
* cell instance $45585 r0 *1 381.52,77
X$45585 2056 1993 25 44 2104 OR2_X1
* cell instance $45588 r0 *1 382.85,77
X$45588 1426 1760 1970 44 2105 25 OAI21_X1
* cell instance $45589 r0 *1 383.61,77
X$45589 2057 2045 2067 25 44 NOR2_X4
* cell instance $45590 r0 *1 385.32,77
X$45590 1761 1735 2103 44 25 2059 MUX2_X2
* cell instance $45592 r0 *1 387.22,77
X$45592 1760 1842 1737 25 44 2150 MUX2_X1
* cell instance $45593 m0 *1 388.17,77
X$45593 1995 1969 2060 2017 2048 2014 44 25 AOI221_X2
* cell instance $45596 m0 *1 391.02,77
X$45596 1912 2014 25 44 2015 XNOR2_X2
* cell instance $45597 m0 *1 392.92,77
X$45597 2014 1912 44 2089 25 XOR2_X2
* cell instance $45600 m0 *1 397.86,77
X$45600 1844 2063 2064 25 44 2049 NOR3_X1
* cell instance $45601 m0 *1 398.62,77
X$45601 2049 2016 1765 44 1883 25 OAI21_X1
* cell instance $45602 m0 *1 399.38,77
X$45602 1882 2065 2017 25 2016 44 AOI21_X1
* cell instance $45603 m0 *1 400.14,77
X$45603 1926 1882 2017 2065 2109 44 25 AOI211_X2
* cell instance $45608 r0 *1 388.55,77
X$45608 2059 1626 25 44 2060 NAND2_X1
* cell instance $45611 r0 *1 392.54,77
X$45611 2061 44 1884 25 BUF_X4
* cell instance $45614 r0 *1 394.82,77
X$45614 2061 25 44 764 INV_X4
* cell instance $45617 r0 *1 396.34,77
X$45617 2059 2063 2064 44 2107 25 NOR3_X2
* cell instance $45620 r0 *1 399.57,77
X$45620 1882 1831 1765 25 44 2108 NAND3_X1
* cell instance $45621 r0 *1 400.33,77
X$45621 2065 2017 1831 1882 44 25 2111 AND4_X1
* cell instance $45623 r0 *1 404.51,77
X$45623 2151 2087 2068 1274 1317 2018 25 44 2066 OAI33_X1
* cell instance $45625 r0 *1 406.6,77
X$45625 2066 1886 2086 2088 2069 44 25 AOI211_X2
* cell instance $45627 m0 *1 407.55,77
X$45627 2068 1385 25 44 2088 NOR2_X1
* cell instance $45629 m0 *1 408.69,77
X$45629 1848 2018 25 44 1928 NAND2_X1
* cell instance $45635 r0 *1 409.64,77
X$45635 1887 2069 1539 2139 2070 44 25 AOI211_X2
* cell instance $45636 m0 *1 410.59,77
X$45636 2068 25 44 1952 INV_X2
* cell instance $45645 r0 *1 416.29,77
X$45645 2114 1386 25 44 2072 NOR2_X1
* cell instance $45646 m0 *1 417.05,77
X$45646 2047 2019 2073 2071 1890 2020 44 25 AOI221_X2
* cell instance $45648 m0 *1 419.14,77
X$45648 2021 2072 1999 2000 1996 25 44 OAI211_X2
* cell instance $45651 m0 *1 424.08,77
X$45651 2070 1932 1974 25 44 2023 MUX2_X1
* cell instance $45652 m0 *1 425.41,77
X$45652 2046 1932 1974 25 2083 44 AOI21_X2
* cell instance $45656 r0 *1 417.62,77
X$45656 2047 2073 2084 2074 2136 1998 25 44 OAI221_X2
* cell instance $45657 r0 *1 419.71,77
X$45657 2137 2073 2047 2019 2046 44 25 AOI211_X2
* cell instance $45660 r0 *1 422.56,77
X$45660 25 2116 2073 2047 2070 2084 2074 44 OAI221_X4
* cell instance $45663 m0 *1 428.83,77
X$45663 2075 2076 2044 2045 2022 44 25 2024 OAI221_X1
* cell instance $45665 m0 *1 429.97,77
X$45665 2024 25 44 1994 INV_X1
* cell instance $45668 m0 *1 432.63,77
X$45668 2041 1439 2067 25 44 1975 NAND3_X1
* cell instance $45669 m0 *1 433.39,77
X$45669 25 2025 2022 2044 2035 1944 44 NAND4_X4
* cell instance $45672 m0 *1 437.76,77
X$45672 2040 2026 25 44 2041 NOR2_X1
* cell instance $45675 m0 *1 440.04,77
X$45675 1977 25 44 2028 INV_X1
* cell instance $45676 m0 *1 440.42,77
X$45676 2028 1853 25 44 2027 NAND2_X1
* cell instance $45677 m0 *1 440.99,77
X$45677 2027 2026 2028 25 44 2037 MUX2_X1
* cell instance $45678 m0 *1 442.32,77
X$45678 2028 2036 2037 1529 44 25 2038 OAI22_X2
* cell instance $45679 m0 *1 444.03,77
X$45679 1979 2026 1977 25 44 1936 MUX2_X1
* cell instance $45680 m0 *1 445.36,77
X$45680 1978 25 44 1853 INV_X1
* cell instance $45682 m0 *1 451.82,77
X$45682 2079 25 44 1894 INV_X1
* cell instance $45686 r0 *1 428.83,77
X$45686 2076 2131 2075 25 44 1933 OR3_X1
* cell instance $45689 r0 *1 436.62,77
X$45689 2131 2077 1977 25 44 NOR2_X4
* cell instance $45693 r0 *1 443.27,77
X$45693 1978 1529 1482 25 2036 44 AOI21_X1
* cell instance $45696 r0 *1 445.93,77
X$45696 25 1978 2077 2078 1855 44 NOR3_X4
* cell instance $45697 r0 *1 448.59,77
X$45697 1978 2077 2078 25 44 1980 OR3_X2
* cell instance $45699 r0 *1 452.77,77
X$45699 1858 44 1482 25 BUF_X4
* cell instance $45703 r0 *1 455.43,77
X$45703 2080 25 44 1618 BUF_X2
* cell instance $45705 r0 *1 456.38,77
X$45705 1566 2080 1777 25 2029 44 AOI21_X2
* cell instance $45706 m0 *1 457.33,77
X$45706 2034 2030 2029 44 25 1657 OAI21_X2
* cell instance $45712 m0 *1 459.99,77
X$45712 2029 2030 25 44 2033 NOR2_X1
* cell instance $45714 m0 *1 460.56,77
X$45714 2030 2029 44 25 2031 AND2_X1
* cell instance $45715 m0 *1 461.32,77
X$45715 2031 2032 25 44 2034 NAND2_X1
* cell instance $45718 r0 *1 460.37,77
X$45718 2081 44 1529 25 BUF_X4
* cell instance $45720 r0 *1 462.08,77
X$45720 2081 1858 25 1439 44 NAND2_X4
* cell instance $45722 m0 *1 462.27,77
X$45722 25 1716 2033 2032 2031 44 AOI21_X4
* cell instance $46014 m0 *1 326.42,26.6
X$46014 467 158 44 25 536 AND2_X1
* cell instance $46016 m0 *1 327.94,26.6
X$46016 554 25 44 518 INV_X1
* cell instance $46036 r0 *1 326.42,26.6
X$46036 536 555 554 44 25 683 HA_X1
* cell instance $46038 m0 *1 331.74,26.6
X$46038 520 25 44 538 INV_X1
* cell instance $46039 m0 *1 328.7,26.6
X$46039 25 430 502 556 518 503 44 FA_X1
* cell instance $46041 m0 *1 332.31,26.6
X$46041 504 522 405 44 25 521 HA_X1
* cell instance $46042 m0 *1 334.21,26.6
X$46042 521 25 44 557 INV_X1
* cell instance $46045 r0 *1 329.84,26.6
X$46045 406 60 44 25 555 AND2_X1
* cell instance $46047 r0 *1 331.36,26.6
X$46047 25 538 537 539 557 556 44 FA_X1
* cell instance $46050 m0 *1 336.49,26.6
X$46050 406 34 44 25 522 AND2_X1
* cell instance $46052 m0 *1 338.2,26.6
X$46052 523 25 44 603 INV_X1
* cell instance $46055 m0 *1 340.29,26.6
X$46055 25 449 606 505 524 525 44 FA_X1
* cell instance $46064 r0 *1 341.43,26.6
X$46064 34 323 25 44 559 NAND2_X1
* cell instance $46068 r0 *1 343.33,26.6
X$46068 505 25 44 560 INV_X1
* cell instance $46069 r0 *1 343.71,26.6
X$46069 560 506 604 44 25 540 HA_X1
* cell instance $46072 m0 *1 345.99,26.6
X$46072 526 25 44 527 CLKBUF_X3
* cell instance $46073 m0 *1 353.02,26.6
X$46073 507 44 508 25 BUF_X4
* cell instance $46079 r0 *1 347.51,26.6
X$46079 513 25 44 323 CLKBUF_X3
* cell instance $46083 r0 *1 352.07,26.6
X$46083 527 528 436 44 25 577 OAI21_X2
* cell instance $46084 r0 *1 353.4,26.6
X$46084 541 527 436 25 563 44 AOI21_X2
* cell instance $46085 r0 *1 354.73,26.6
X$46085 436 528 509 25 574 44 AOI21_X2
* cell instance $46088 r0 *1 356.63,26.6
X$46088 564 44 579 25 BUF_X4
* cell instance $46091 m0 *1 360.05,26.6
X$46091 530 25 44 565 INV_X1
* cell instance $46093 m0 *1 362.14,26.6
X$46093 471 25 44 511 INV_X1
* cell instance $46098 r0 *1 361.38,26.6
X$46098 565 511 612 44 25 580 HA_X1
* cell instance $46101 m0 *1 365.94,26.6
X$46101 512 25 44 614 INV_X1
* cell instance $46105 r0 *1 367.27,26.6
X$46105 25 297 543 616 566 544 44 FA_X1
* cell instance $46107 m0 *1 368.22,26.6
X$46107 513 47 44 25 566 AND2_X1
* cell instance $46109 m0 *1 372.21,26.6
X$46109 25 219 567 546 533 532 44 FA_X1
* cell instance $46114 r0 *1 373.73,26.6
X$46114 568 25 44 569 INV_X1
* cell instance $46116 r0 *1 374.49,26.6
X$46116 546 25 44 545 INV_X1
* cell instance $46120 r0 *1 376.2,26.6
X$46120 514 25 44 547 INV_X1
* cell instance $46122 m0 *1 379.62,26.6
X$46122 27 25 44 213 BUF_X2
* cell instance $46132 r0 *1 386.65,26.6
X$46132 27 47 44 25 549 AND2_X1
* cell instance $46137 m0 *1 392.92,26.6
X$46137 516 535 761 44 25 562 HA_X1
* cell instance $46143 r0 *1 392.54,26.6
X$46143 213 291 44 25 762 AND2_X1
* cell instance $46145 r0 *1 393.68,26.6
X$46145 562 25 44 561 INV_X1
* cell instance $46150 r0 *1 395.58,26.6
X$46150 406 513 42 27 25 44 609 OR4_X1
* cell instance $46154 r0 *1 399.38,26.6
X$46154 159 877 588 44 25 558 HA_X1
* cell instance $46156 m0 *1 400.52,26.6
X$46156 301 291 186 25 44 534 NOR3_X1
* cell instance $46158 m0 *1 402.8,26.6
X$46158 201 25 44 301 CLKBUF_X3
* cell instance $46161 m0 *1 415.91,26.6
X$46161 531 195 25 44 553 NOR2_X1
* cell instance $46162 m0 *1 416.48,26.6
X$46162 479 529 25 44 531 XOR2_X1
* cell instance $46163 m0 *1 417.62,26.6
X$46163 303 481 25 44 529 NAND2_X1
* cell instance $46170 r0 *1 412.68,26.6
X$46170 25 30 553 43 2895 478 44 DFFR_X2
* cell instance $46172 m0 *1 420.28,26.6
X$46172 303 481 479 480 25 44 550 NAND4_X1
* cell instance $46175 m0 *1 421.42,26.6
X$46175 517 195 25 44 519 NOR2_X1
* cell instance $46176 m0 *1 421.99,26.6
X$46176 25 30 519 43 482 480 44 DFFR_X2
* cell instance $46462 m0 *1 334.4,57.4
X$46462 25 1373 1400 1370 1452 1341 44 OR4_X4
* cell instance $46464 r0 *1 335.54,57.4
X$46464 1268 1134 1141 25 44 1418 NAND3_X1
* cell instance $46465 r0 *1 336.3,57.4
X$46465 1420 1418 25 44 1419 OR2_X1
* cell instance $46468 m0 *1 338.96,57.4
X$46468 1146 1371 1134 1141 1136 1452 44 25 AOI221_X2
* cell instance $46472 r0 *1 339.34,57.4
X$46472 1058 1264 1144 1266 1585 44 25 AOI211_X2
* cell instance $46474 r0 *1 341.24,57.4
X$46474 1264 1146 25 44 1420 NAND2_X1
* cell instance $46475 r0 *1 341.81,57.4
X$46475 1144 1268 1266 25 44 1505 NAND3_X2
* cell instance $46477 m0 *1 342.95,57.4
X$46477 1291 1304 1267 25 44 1403 NAND3_X2
* cell instance $46478 m0 *1 345.04,57.4
X$46478 1142 1372 25 44 1454 NOR2_X1
* cell instance $46483 r0 *1 343.71,57.4
X$46483 1267 1304 1291 44 25 1464 AND3_X2
* cell instance $46486 r0 *1 345.42,57.4
X$46486 25 1454 1403 1349 1421 1455 44 OAI211_X4
* cell instance $46487 m0 *1 347.7,57.4
X$46487 1046 1061 1107 44 25 1544 OAI21_X4
* cell instance $46492 r0 *1 349.41,57.4
X$46492 1266 1422 44 25 1455 AND2_X2
* cell instance $46495 r0 *1 351.31,57.4
X$46495 1422 1266 25 44 1493 NAND2_X2
* cell instance $46496 m0 *1 352.83,57.4
X$46496 1374 1406 1407 44 25 1465 OAI21_X2
* cell instance $46497 m0 *1 352.07,57.4
X$46497 1146 1268 44 25 1374 AND2_X1
* cell instance $46501 m0 *1 366.51,57.4
X$46501 1376 1270 1375 25 44 1511 NAND3_X2
* cell instance $46504 r0 *1 352.26,57.4
X$46504 25 1374 1147 1587 1422 1266 44 AOI22_X4
* cell instance $46514 r0 *1 366.7,57.4
X$46514 1375 1270 1376 44 25 1467 AND3_X1
* cell instance $46515 r0 *1 367.65,57.4
X$46515 1376 1270 1375 25 44 1547 NAND3_X2
* cell instance $46519 m0 *1 371.45,57.4
X$46519 1377 1381 1375 25 1423 44 AOI21_X1
* cell instance $46522 r0 *1 371.64,57.4
X$46522 1378 1457 1423 1456 1424 1878 44 25 AOI221_X2
* cell instance $46523 m0 *1 372.78,57.4
X$46523 1375 1381 25 44 1456 NAND2_X1
* cell instance $46528 m0 *1 375.82,57.4
X$46528 1063 1379 25 44 1380 XNOR2_X2
* cell instance $46532 r0 *1 373.73,57.4
X$46532 1145 978 25 44 1469 NOR2_X1
* cell instance $46534 r0 *1 374.49,57.4
X$46534 1470 1421 1241 44 1457 25 OAI21_X1
* cell instance $46535 r0 *1 375.25,57.4
X$46535 1152 978 25 44 1471 NAND2_X1
* cell instance $46538 r0 *1 376.96,57.4
X$46538 25 1379 1145 1375 1472 44 AOI21_X4
* cell instance $46539 r0 *1 379.43,57.4
X$46539 1152 1241 25 44 1473 XNOR2_X2
* cell instance $46541 r0 *1 384.37,57.4
X$46541 1425 25 44 1497 INV_X1
* cell instance $46542 r0 *1 384.75,57.4
X$46542 1428 1425 1472 25 44 1538 NAND3_X2
* cell instance $46543 m0 *1 386.46,57.4
X$46543 1382 1426 25 44 1428 NOR2_X1
* cell instance $46544 m0 *1 385.7,57.4
X$46544 1426 1382 25 44 1427 OR2_X1
* cell instance $46546 m0 *1 387.22,57.4
X$46546 25 1272 1430 1425 1382 1375 44 NOR4_X4
* cell instance $46549 r0 *1 386.08,57.4
X$46549 1498 1425 1382 25 44 1470 OR3_X2
* cell instance $46550 r0 *1 387.22,57.4
X$46550 1425 1381 1428 25 1429 44 AOI21_X2
* cell instance $46553 r0 *1 389.12,57.4
X$46553 1430 44 1426 25 BUF_X4
* cell instance $46557 m0 *1 391.97,57.4
X$46557 1383 1361 25 44 1460 OR2_X1
* cell instance $46559 m0 *1 392.73,57.4
X$46559 1460 44 1554 25 BUF_X4
* cell instance $46561 m0 *1 394.25,57.4
X$46561 1119 1384 25 1430 44 NAND2_X4
* cell instance $46563 r0 *1 391.78,57.4
X$46563 1361 1383 1644 25 44 NOR2_X4
* cell instance $46564 r0 *1 393.49,57.4
X$46564 1430 1272 1461 25 44 NOR2_X4
* cell instance $46566 m0 *1 396.53,57.4
X$46566 1384 44 1431 25 BUF_X4
* cell instance $46574 r0 *1 400.33,57.4
X$46574 1416 1272 1501 25 44 NOR2_X4
* cell instance $46577 m0 *1 402.04,57.4
X$46577 1385 44 1386 25 BUF_X4
* cell instance $46580 m0 *1 408.12,57.4
X$46580 737 633 25 44 1433 NAND2_X2
* cell instance $46582 m0 *1 409.26,57.4
X$46582 1434 737 25 44 1280 XNOR2_X2
* cell instance $46586 m0 *1 415.91,57.4
X$46586 1434 1431 25 44 1258 NAND2_X2
* cell instance $46587 m0 *1 416.86,57.4
X$46587 1387 1388 1258 1162 25 44 1390 AOI22_X2
* cell instance $46589 m0 *1 420.09,57.4
X$46589 1323 1390 25 44 1459 OR2_X1
* cell instance $46590 m0 *1 420.85,57.4
X$46590 25 1323 1435 1095 1459 1119 44 AOI22_X4
* cell instance $46595 m0 *1 434.15,57.4
X$46595 1082 1032 1326 1438 25 44 1458 OR4_X1
* cell instance $46597 m0 *1 438.33,57.4
X$46597 1480 1442 1391 25 1402 44 AOI21_X2
* cell instance $46601 r0 *1 403.18,57.4
X$46601 25 1502 1462 915 1433 1436 44 AOI22_X4
* cell instance $46602 r0 *1 406.41,57.4
X$46602 1432 1554 1433 44 25 1218 MUX2_X2
* cell instance $46606 r0 *1 410.21,57.4
X$46606 633 25 44 1323 INV_X2
* cell instance $46610 r0 *1 417.81,57.4
X$46610 1478 1477 1281 1431 1434 1408 44 25 AOI221_X2
* cell instance $46614 r0 *1 421.23,57.4
X$46614 1164 1390 25 44 1435 XNOR2_X2
* cell instance $46618 r0 *1 428.45,57.4
X$46618 1326 1438 25 44 1122 OR2_X2
* cell instance $46620 r0 *1 430.16,57.4
X$46620 1458 1293 1437 25 1499 44 AOI21_X2
* cell instance $46623 r0 *1 434.72,57.4
X$46623 1441 1439 1440 25 44 1225 MUX2_X1
* cell instance $46625 r0 *1 437.57,57.4
X$46625 1436 1391 1442 25 1169 44 AOI21_X1
* cell instance $46626 r0 *1 438.33,57.4
X$46626 1443 1495 1479 25 1082 44 NAND3_X4
* cell instance $46627 r0 *1 440.8,57.4
X$46627 1495 1443 1479 44 25 1444 AND3_X1
* cell instance $46629 m0 *1 441.56,57.4
X$46629 1171 1391 1442 25 1035 44 AOI21_X1
* cell instance $46630 m0 *1 443.84,57.4
X$46630 680 1392 1441 25 44 1401 NOR3_X1
* cell instance $46632 r0 *1 441.75,57.4
X$46632 1481 1083 25 44 1480 NAND2_X2
* cell instance $46633 r0 *1 442.7,57.4
X$46633 1441 1451 1447 44 25 1442 OAI21_X2
* cell instance $46635 m0 *1 446.69,57.4
X$46635 1392 1441 1081 680 44 1453 25 NOR4_X2
* cell instance $46636 m0 *1 444.98,57.4
X$46636 1453 1399 44 999 25 XOR2_X2
* cell instance $46643 r0 *1 451.44,57.4
X$46643 1449 1446 44 25 1397 XNOR2_X1
* cell instance $46645 m0 *1 453.91,57.4
X$46645 1395 1394 25 44 1173 XNOR2_X2
* cell instance $46646 m0 *1 453.34,57.4
X$46646 680 1393 25 44 1394 NOR2_X1
* cell instance $46697 r0 *1 455.81,57.4
X$46697 1448 1451 1447 25 44 1450 NOR3_X1
* cell instance $46698 r0 *1 456.57,57.4
X$46698 1450 1439 1532 25 1179 44 AOI21_X2
* cell instance $46932 m0 *1 340.1,63
X$46932 1141 1504 25 44 1578 XNOR2_X2
* cell instance $46933 m0 *1 342,63
X$46933 1505 1420 25 44 1542 NOR2_X2
* cell instance $46953 r0 *1 340.86,63
X$46953 1236 1586 25 44 1628 NAND2_X1
* cell instance $46955 r0 *1 341.62,63
X$46955 1092 1585 25 1586 44 OR2_X4
* cell instance $46959 m0 *1 344.09,63
X$46959 1047 1570 1543 25 1622 44 AOI21_X2
* cell instance $46960 m0 *1 346.94,63
X$46960 1349 1455 25 44 1588 NOR2_X2
* cell instance $46963 m0 *1 348.84,63
X$46963 1544 1545 44 25 1630 AND2_X2
* cell instance $46967 r0 *1 344.66,63
X$46967 1587 1630 25 44 1631 NOR2_X1
* cell instance $46968 r0 *1 345.23,63
X$46968 25 1631 1632 1667 1622 1589 44 AOI22_X4
* cell instance $46972 r0 *1 349.79,63
X$46972 25 1693 1405 1590 1587 44 AOI21_X4
* cell instance $46974 m0 *1 350.93,63
X$46974 1545 1544 25 1590 44 NAND2_X4
* cell instance $46978 r0 *1 352.83,63
X$46978 1590 1047 1591 44 25 1668 OAI21_X2
* cell instance $46980 m0 *1 353.78,63
X$46980 1546 44 1381 25 BUF_X4
* cell instance $46984 r0 *1 354.35,63
X$46984 1668 1346 1472 25 44 1670 NAND3_X2
* cell instance $46987 m0 *1 357.96,63
X$46987 25 1579 1535 1507 1534 1592 44 NAND4_X4
* cell instance $46989 m0 *1 361.38,63
X$46989 1547 1313 1545 1544 1595 44 25 AOI211_X2
* cell instance $46990 m0 *1 363.09,63
X$46990 1547 1313 25 44 1593 NOR2_X2
* cell instance $46993 r0 *1 358.15,63
X$46993 1047 1421 1591 44 25 1633 OAI21_X2
* cell instance $46998 r0 *1 362.14,63
X$46998 1634 1593 44 25 1594 AND2_X1
* cell instance $46999 r0 *1 362.9,63
X$46999 1310 1581 25 44 1634 NOR2_X1
* cell instance $47001 r0 *1 363.66,63
X$47001 1509 1581 25 44 1675 NOR2_X1
* cell instance $47003 m0 *1 366.89,63
X$47003 1310 1472 1548 25 1635 44 AOI21_X2
* cell instance $47004 m0 *1 364.42,63
X$47004 25 1838 1535 1381 1467 44 AOI21_X4
* cell instance $47005 m0 *1 368.22,63
X$47005 1548 25 44 1597 INV_X1
* cell instance $47010 r0 *1 364.61,63
X$47010 1595 1596 25 44 1676 NOR2_X1
* cell instance $47013 r0 *1 366.32,63
X$47013 1509 1512 25 1596 44 NAND2_X4
* cell instance $47014 r0 *1 368.03,63
X$47014 1597 1509 1510 44 1636 25 NOR3_X2
* cell instance $47015 r0 *1 369.36,63
X$47015 1509 1510 1597 44 25 1638 OAI21_X2
* cell instance $47019 m0 *1 378.86,63
X$47019 1549 1550 1626 44 1701 25 OAI21_X1
* cell instance $47022 m0 *1 383.61,63
X$47022 1515 1516 25 44 1599 NAND2_X1
* cell instance $47025 m0 *1 385.13,63
X$47025 1538 1517 25 44 1700 NAND2_X1
* cell instance $47031 r0 *1 384.94,63
X$47031 1601 1600 25 44 1704 NOR2_X1
* cell instance $47032 r0 *1 385.51,63
X$47032 25 1601 1600 1518 1756 1429 44 OAI22_X4
* cell instance $47034 m0 *1 386.84,63
X$47034 1518 1429 25 44 1641 NOR2_X1
* cell instance $47037 m0 *1 389.88,63
X$47037 1065 1381 1552 1414 44 25 1601 AND4_X1
* cell instance $47042 r0 *1 389.69,63
X$47042 1519 1381 1552 25 1600 44 AOI21_X2
* cell instance $47045 r0 *1 392.92,63
X$47045 1519 1552 25 44 1736 NOR2_X2
* cell instance $47048 m0 *1 394.44,63
X$47048 1627 877 1553 44 25 1643 OAI21_X2
* cell instance $47051 r0 *1 394.82,63
X$47051 1602 1554 1472 25 44 1627 NAND3_X1
* cell instance $47054 r0 *1 396.15,63
X$47054 1472 1644 44 25 1645 XNOR2_X1
* cell instance $47055 m0 *1 397.1,63
X$47055 1065 1421 1474 25 44 1647 OR3_X2
* cell instance $47058 m0 *1 398.43,63
X$47058 1317 1274 1552 25 44 NOR2_X4
* cell instance $47061 m0 *1 406.98,63
X$47061 1555 44 633 25 BUF_X4
* cell instance $47062 m0 *1 408.31,63
X$47062 1556 1584 25 44 1475 XNOR2_X2
* cell instance $47063 m0 *1 410.21,63
X$47063 1556 25 44 1432 INV_X1
* cell instance $47064 m0 *1 410.59,63
X$47064 1560 1432 1323 1539 25 44 1688 NAND4_X1
* cell instance $47065 m0 *1 411.54,63
X$47065 1560 1539 25 44 1584 NAND2_X1
* cell instance $47069 r0 *1 397.48,63
X$47069 1414 1647 25 44 1602 XNOR2_X2
* cell instance $47073 r0 *1 403.37,63
X$47073 1416 1498 1626 25 44 NOR2_X4
* cell instance $47074 r0 *1 405.08,63
X$47074 1364 1254 1501 44 25 1686 AND3_X2
* cell instance $47077 r0 *1 407.93,63
X$47077 1644 1555 1556 25 44 1687 MUX2_X1
* cell instance $47078 r0 *1 409.26,63
X$47078 1687 982 25 44 1624 NOR2_X1
* cell instance $47080 r0 *1 410.02,63
X$47080 1386 1432 1560 25 44 1649 OR3_X1
* cell instance $47081 r0 *1 410.97,63
X$47081 1689 1688 1691 25 44 1692 NAND3_X1
* cell instance $47082 r0 *1 411.73,63
X$47082 1560 1556 633 1539 25 44 1691 NAND4_X1
* cell instance $47084 m0 *1 414.2,63
X$47084 25 1388 1523 1522 1583 1319 44 NAND4_X4
* cell instance $47090 r0 *1 414.77,63
X$47090 25 1388 1650 1603 1298 1692 1624 44 OAI221_X4
* cell instance $47091 r0 *1 417.24,63
X$47091 1476 1650 1603 44 25 1583 OAI21_X2
* cell instance $47094 m0 *1 418.76,63
X$47094 1171 1474 1604 44 25 1478 OAI21_X2
* cell instance $47096 r0 *1 418.95,63
X$47096 1604 1171 1474 44 1603 25 NOR3_X2
* cell instance $47098 m0 *1 421.42,63
X$47098 731 1556 44 25 1605 XNOR2_X1
* cell instance $47100 m0 *1 422.56,63
X$47100 25 1499 1556 1555 1651 731 44 OAI22_X4
* cell instance $47106 r0 *1 422.37,63
X$47106 1474 1605 1652 25 44 1164 OR3_X2
* cell instance $47110 r0 *1 428.26,63
X$47110 1607 1608 1606 969 44 25 991 AND4_X2
* cell instance $47111 m0 *1 428.64,63
X$47111 1326 1610 1555 1330 25 44 1607 OR4_X1
* cell instance $47113 m0 *1 429.78,63
X$47113 1165 1285 1540 1580 25 44 1609 NAND4_X1
* cell instance $47114 m0 *1 430.73,63
X$47114 1540 1326 1610 44 1608 25 OAI21_X1
* cell instance $47118 r0 *1 429.59,63
X$47118 1606 1608 25 44 1655 NAND2_X1
* cell instance $47119 r0 *1 430.16,63
X$47119 1609 1726 1607 25 44 1654 NAND3_X1
* cell instance $47122 m0 *1 434.34,63
X$47122 1558 1557 25 44 1611 OR2_X1
* cell instance $47124 m0 *1 435.1,63
X$47124 1557 1558 25 44 1612 NOR2_X1
* cell instance $47125 m0 *1 435.67,63
X$47125 1559 1343 25 44 1558 NOR2_X1
* cell instance $47126 m0 *1 436.24,63
X$47126 1343 1559 1557 25 44 1560 OR3_X2
* cell instance $47127 m0 *1 437.38,63
X$47127 1443 1495 25 44 1559 NAND2_X1
* cell instance $47128 m0 *1 437.95,63
X$47128 1577 1615 1561 25 1613 44 AOI21_X2
* cell instance $47129 m0 *1 439.28,63
X$47129 1615 1443 1495 25 44 1576 NAND3_X1
* cell instance $47131 m0 *1 440.23,63
X$47131 1576 1343 25 44 1577 NOR2_X1
* cell instance $47136 r0 *1 434.91,63
X$47136 1613 25 44 1684 INV_X1
* cell instance $47137 r0 *1 435.29,63
X$47137 1681 1613 1611 25 44 1438 NAND3_X2
* cell instance $47138 r0 *1 436.62,63
X$47138 1614 1709 1610 25 44 1681 NOR3_X1
* cell instance $47141 r0 *1 444.22,63
X$47141 1657 1617 25 44 1616 NOR2_X1
* cell instance $47142 r0 *1 444.79,63
X$47142 1658 1657 1617 44 1614 25 NOR3_X2
* cell instance $47145 r0 *1 447.07,63
X$47145 1672 1659 25 44 1658 NOR2_X1
* cell instance $47318 m0 *1 335.16,54.6
X$47318 1195 1057 1302 1268 1141 1341 44 25 AOI221_X2
* cell instance $47320 m0 *1 340.48,54.6
X$47320 1059 1144 1106 25 44 1303 MUX2_X1
* cell instance $47322 r0 *1 335.54,54.6
X$47322 1268 1134 1141 25 44 1370 NOR3_X1
* cell instance $47324 r0 *1 336.68,54.6
X$47324 1419 1292 1302 25 1400 44 AOI21_X1
* cell instance $47327 r0 *1 338.39,54.6
X$47327 1140 1107 1292 44 1371 25 OAI21_X1
* cell instance $47330 r0 *1 340.1,54.6
X$47330 1136 1146 1264 25 1372 44 AOI21_X2
* cell instance $47331 r0 *1 341.43,54.6
X$47331 1372 1267 1303 25 1302 44 AOI21_X2
* cell instance $47332 m0 *1 342.38,54.6
X$47332 1110 1106 44 25 1304 AND2_X1
* cell instance $47338 r0 *1 345.99,54.6
X$47338 25 1061 1107 1292 1291 1405 44 NOR4_X4
* cell instance $47340 m0 *1 349.79,54.6
X$47340 25 1349 1202 1350 1352 44 AOI21_X4
* cell instance $47342 m0 *1 352.26,54.6
X$47342 1134 1351 1292 25 44 1352 OR3_X1
* cell instance $47343 m0 *1 353.21,54.6
X$47343 1112 1140 25 44 1351 NOR2_X1
* cell instance $47345 m0 *1 355.3,54.6
X$47345 1150 959 958 44 1308 25 NOR3_X2
* cell instance $47348 m0 *1 358.34,54.6
X$47348 1269 1145 25 44 1409 NAND2_X1
* cell instance $47350 m0 *1 359.67,54.6
X$47350 1150 959 958 1357 44 1307 25 NOR4_X2
* cell instance $47352 m0 *1 361.57,54.6
X$47352 1149 1355 25 44 1310 XNOR2_X2
* cell instance $47353 m0 *1 363.47,54.6
X$47353 1311 1148 1018 25 44 1355 NAND3_X2
* cell instance $47357 r0 *1 351.69,54.6
X$47357 1141 1134 1307 44 25 1406 AND3_X1
* cell instance $47358 r0 *1 352.64,54.6
X$47358 1292 1351 1134 25 44 1407 NOR3_X1
* cell instance $47360 r0 *1 353.59,54.6
X$47360 25 1308 1409 1146 1268 1422 44 NAND4_X4
* cell instance $47364 r0 *1 359.1,54.6
X$47364 958 1353 25 44 1512 XNOR2_X2
* cell instance $47367 r0 *1 361.95,54.6
X$47367 959 1355 25 44 1509 XNOR2_X2
* cell instance $47370 r0 *1 364.8,54.6
X$47370 1018 1312 25 44 1411 XNOR2_X2
* cell instance $47372 m0 *1 365.94,54.6
X$47372 1269 1150 25 44 1312 NOR2_X2
* cell instance $47374 m0 *1 371.45,54.6
X$47374 1311 1063 25 44 1377 NAND2_X1
* cell instance $47377 r0 *1 366.7,54.6
X$47377 1111 1312 25 44 1625 XNOR2_X2
* cell instance $47379 r0 *1 371.64,54.6
X$47379 1209 1063 25 44 1378 NOR2_X1
* cell instance $47382 m0 *1 375.25,54.6
X$47382 1271 1241 1209 1211 25 44 1314 NAND4_X1
* cell instance $47383 m0 *1 373.92,54.6
X$47383 1253 1020 1063 44 1424 25 NOR3_X2
* cell instance $47384 m0 *1 376.2,54.6
X$47384 1112 1063 25 44 1359 NAND2_X2
* cell instance $47385 m0 *1 377.15,54.6
X$47385 1271 1152 25 44 1315 NOR2_X2
* cell instance $47386 m0 *1 378.1,54.6
X$47386 904 1359 25 44 1360 XNOR2_X2
* cell instance $47390 r0 *1 374.3,54.6
X$47390 1271 1145 1413 1241 1314 1376 25 44 OAI221_X2
* cell instance $47391 r0 *1 376.39,54.6
X$47391 1152 1211 25 44 1413 NAND2_X1
* cell instance $47392 r0 *1 376.96,54.6
X$47392 1020 1315 25 44 1415 XNOR2_X2
* cell instance $47396 r0 *1 380.19,54.6
X$47396 1211 1315 25 44 1416 XNOR2_X2
* cell instance $47398 m0 *1 381.14,54.6
X$47398 870 1359 25 44 1364 XNOR2_X2
* cell instance $47403 r0 *1 389.69,54.6
X$47403 1414 1114 1383 44 25 1382 OAI21_X2
* cell instance $47405 m0 *1 391.21,54.6
X$47405 1214 1316 25 44 1414 XNOR2_X2
* cell instance $47411 r0 *1 391.21,54.6
X$47411 1065 1274 1383 25 44 NOR2_X4
* cell instance $47416 r0 *1 395.77,54.6
X$47416 1275 1385 25 44 1384 NOR2_X2
* cell instance $47418 r0 *1 396.91,54.6
X$47418 1272 44 1333 25 BUF_X4
* cell instance $47421 r0 *1 399.38,54.6
X$47421 1274 1317 25 44 1417 OR2_X1
* cell instance $47422 r0 *1 400.14,54.6
X$47422 1417 44 1385 25 BUF_X4
* cell instance $47424 r0 *1 401.85,54.6
X$47424 1260 44 1100 25 BUF_X4
* cell instance $47426 m0 *1 404.32,54.6
X$47426 25 1278 1318 1218 944 982 44 OAI22_X4
* cell instance $47434 r0 *1 410.97,54.6
X$47434 1319 25 44 737 INV_X2
* cell instance $47437 r0 *1 412.11,54.6
X$47437 1410 1412 1320 44 25 1025 MUX2_X2
* cell instance $47438 m0 *1 413.44,54.6
X$47438 1162 25 44 1320 INV_X1
* cell instance $47442 m0 *1 414.77,54.6
X$47442 1258 25 44 1321 INV_X1
* cell instance $47444 m0 *1 415.91,54.6
X$47444 1074 1367 1162 1322 25 44 1368 NOR4_X1
* cell instance $47445 m0 *1 416.86,54.6
X$47445 1191 1258 44 25 1476 AND2_X1
* cell instance $47448 m0 *1 422.18,54.6
X$47448 25 1365 1281 1363 1322 1324 44 OAI22_X4
* cell instance $47450 m0 *1 426.93,54.6
X$47450 1327 1325 25 44 1363 NOR2_X2
* cell instance $47451 m0 *1 427.88,54.6
X$47451 1285 1326 1329 25 1327 44 AOI21_X1
* cell instance $47452 m0 *1 428.64,54.6
X$47452 1165 1328 1123 25 44 1330 NOR3_X1
* cell instance $47453 m0 *1 429.4,54.6
X$47453 1356 1329 1325 25 44 1354 MUX2_X1
* cell instance $47454 m0 *1 430.73,54.6
X$47454 1331 1293 25 44 1329 NAND2_X1
* cell instance $47458 m0 *1 433.77,54.6
X$47458 1173 1348 25 44 1123 XNOR2_X2
* cell instance $47460 m0 *1 435.86,54.6
X$47460 1333 1345 725 25 1347 44 AOI21_X2
* cell instance $47461 m0 *1 437.19,54.6
X$47461 25 1348 1347 1084 1332 44 AOI21_X4
* cell instance $47463 m0 *1 439.85,54.6
X$47463 1334 1336 1082 25 44 1335 NAND3_X2
* cell instance $47465 m0 *1 441.37,54.6
X$47465 1337 1336 44 1325 25 XOR2_X2
* cell instance $47469 r0 *1 414.58,54.6
X$47469 1321 1387 1388 25 1412 44 AOI21_X1
* cell instance $47471 r0 *1 415.72,54.6
X$47471 1367 1322 25 44 1387 NOR2_X2
* cell instance $47472 r0 *1 416.67,54.6
X$47472 1387 1388 25 44 1389 NAND2_X1
* cell instance $47474 r0 *1 417.62,54.6
X$47474 1389 1408 1258 44 1410 25 OAI21_X1
* cell instance $47477 r0 *1 427.5,54.6
X$47477 1404 1329 1328 44 1324 25 NOR3_X2
* cell instance $47478 r0 *1 428.83,54.6
X$47478 1165 1326 44 1404 25 XOR2_X2
* cell instance $47479 r0 *1 430.54,54.6
X$47479 1331 1325 44 25 1437 AND2_X1
* cell instance $47482 r0 *1 437.57,54.6
X$47482 1345 1402 25 44 1332 XNOR2_X2
* cell instance $47483 r0 *1 439.47,54.6
X$47483 25 1326 1287 1335 1396 44 AOI21_X4
* cell instance $47487 r0 *1 444.03,54.6
X$47487 1035 1401 1083 44 1398 25 OAI21_X1
* cell instance $47491 r0 *1 446.12,54.6
X$47491 1398 1399 44 1340 25 XOR2_X2
* cell instance $47493 m0 *1 449.73,54.6
X$47493 1397 1333 25 44 1174 NAND2_X2
* cell instance $47495 m0 *1 450.68,54.6
X$47495 1130 1339 25 44 1336 XNOR2_X2
* cell instance $47496 m0 *1 452.58,54.6
X$47496 1176 725 25 44 1339 NOR2_X1
* cell instance $47497 m0 *1 453.15,54.6
X$47497 1231 1338 25 44 1396 XNOR2_X2
* cell instance $47799 m0 *1 340.67,60.2
X$47799 1110 1268 1146 25 44 1504 NAND3_X2
* cell instance $47802 m0 *1 343.52,60.2
X$47802 1420 1042 25 44 1570 NAND2_X1
* cell instance $47805 r0 *1 340.86,60.2
X$47805 1140 1504 44 25 1629 XNOR2_X1
* cell instance $47807 r0 *1 343.52,60.2
X$47807 1267 1505 44 25 1571 AND2_X1
* cell instance $47808 r0 *1 344.28,60.2
X$47808 1505 1267 25 44 1543 NAND2_X1
* cell instance $47809 r0 *1 344.85,60.2
X$47809 1109 1506 1571 44 25 1572 OAI21_X2
* cell instance $47810 m0 *1 345.99,60.2
X$47810 1372 1142 25 44 1463 OR2_X2
* cell instance $47811 m0 *1 345.23,60.2
X$47811 1046 1146 1264 25 1506 44 AOI21_X1
* cell instance $47813 m0 *1 347.13,60.2
X$47813 1042 1146 1264 25 1545 44 NAND3_X4
* cell instance $47816 m0 *1 350.17,60.2
X$47816 1464 1463 1534 25 44 NOR2_X4
* cell instance $47818 m0 *1 351.88,60.2
X$47818 1464 1463 1465 1493 1546 44 25 AOI211_X2
* cell instance $47819 m0 *1 353.59,60.2
X$47819 1465 1493 25 1507 44 NAND2_X4
* cell instance $47823 m0 *1 360.05,60.2
X$47823 25 1309 1310 1313 1511 1508 44 NOR4_X4
* cell instance $47829 r0 *1 359.29,60.2
X$47829 1507 1534 1579 1535 44 25 1623 AND4_X2
* cell instance $47832 r0 *1 361.19,60.2
X$47832 1547 25 44 1579 INV_X1
* cell instance $47835 r0 *1 362.71,60.2
X$47835 1309 44 1581 25 BUF_X4
* cell instance $47836 r0 *1 364.04,60.2
X$47836 1466 1510 1511 44 25 1750 OAI21_X2
* cell instance $47837 m0 *1 364.8,60.2
X$47837 1466 25 44 1535 INV_X2
* cell instance $47842 r0 *1 365.37,60.2
X$47842 1207 1509 1512 1467 25 1591 44 NAND4_X2
* cell instance $47843 r0 *1 367.08,60.2
X$47843 1511 1313 25 44 1548 NOR2_X1
* cell instance $47847 r0 *1 372.97,60.2
X$47847 1468 1513 1471 44 25 1639 OAI21_X4
* cell instance $47848 m0 *1 375.06,60.2
X$47848 1248 1375 1472 25 1513 44 AOI21_X2
* cell instance $47849 m0 *1 373.35,60.2
X$47849 1424 1469 1470 1510 44 25 1468 OAI22_X2
* cell instance $47850 m0 *1 376.39,60.2
X$47850 978 1379 25 44 1702 XNOR2_X2
* cell instance $47854 r0 *1 378.48,60.2
X$47854 1473 1472 1375 25 1549 44 AOI21_X1
* cell instance $47855 r0 *1 379.24,60.2
X$47855 1514 1470 1510 25 44 1550 NOR3_X1
* cell instance $47856 r0 *1 380,60.2
X$47856 1473 1375 1472 25 44 1598 NAND3_X2
* cell instance $47857 m0 *1 380.38,60.2
X$47857 1473 25 44 1514 INV_X1
* cell instance $47861 m0 *1 384.56,60.2
X$47861 1497 1421 1427 44 25 1517 OAI21_X2
* cell instance $47863 m0 *1 386.08,60.2
X$47863 1427 1497 1421 44 1518 25 NOR3_X2
* cell instance $47865 r0 *1 381.33,60.2
X$47865 1514 1510 1470 44 25 1551 OAI21_X2
* cell instance $47867 r0 *1 383.04,60.2
X$47867 25 1515 1516 1696 1538 1517 44 AOI22_X4
* cell instance $47870 m0 *1 389.12,60.2
X$47870 1421 1385 1361 1383 1414 1516 25 44 OAI221_X2
* cell instance $47871 m0 *1 387.79,60.2
X$47871 1381 44 1472 25 BUF_X4
* cell instance $47873 r0 *1 388.55,60.2
X$47873 1421 44 1510 25 BUF_X4
* cell instance $47874 r0 *1 389.88,60.2
X$47874 1552 1381 1065 1414 25 1515 44 NAND4_X2
* cell instance $47876 m0 *1 391.59,60.2
X$47876 1414 1383 1361 44 25 1519 OAI21_X2
* cell instance $47882 r0 *1 394.06,60.2
X$47882 1472 1260 1519 25 44 1553 OR3_X1
* cell instance $47884 m0 *1 395.77,60.2
X$47884 1520 1190 25 1498 44 NAND2_X4
* cell instance $47888 r0 *1 396.91,60.2
X$47888 1260 1552 25 1474 44 NAND2_X4
* cell instance $47889 m0 *1 399.57,60.2
X$47889 1520 44 1083 25 BUF_X4
* cell instance $47890 m0 *1 397.86,60.2
X$47890 1222 1474 1520 25 44 NOR2_X4
* cell instance $47892 m0 *1 403.94,60.2
X$47892 1323 1386 1503 44 25 1502 OAI21_X2
* cell instance $47893 m0 *1 405.27,60.2
X$47893 1475 1319 44 25 1503 XNOR2_X1
* cell instance $47894 m0 *1 406.41,60.2
X$47894 1475 982 25 44 1541 NAND2_X1
* cell instance $47897 m0 *1 408.69,60.2
X$47897 1475 1555 44 1434 25 XOR2_X2
* cell instance $47898 m0 *1 410.4,60.2
X$47898 1539 44 982 25 BUF_X4
* cell instance $47906 r0 *1 406.03,60.2
X$47906 1475 1319 1541 25 44 1521 MUX2_X1
* cell instance $47907 r0 *1 407.36,60.2
X$47907 1521 633 25 44 1462 NAND2_X1
* cell instance $47910 m0 *1 414.58,60.2
X$47910 1322 25 44 1522 INV_X1
* cell instance $47913 m0 *1 418,60.2
X$47913 1477 1478 25 44 1162 NAND2_X2
* cell instance $47914 m0 *1 418.95,60.2
X$47914 1408 1322 25 44 1500 NOR2_X1
* cell instance $47919 r0 *1 417.05,60.2
X$47919 1367 25 44 1523 INV_X1
* cell instance $47920 r0 *1 417.43,60.2
X$47920 1523 1388 25 44 1524 NAND2_X1
* cell instance $47925 r0 *1 426.55,60.2
X$47925 1500 1524 1582 1438 25 44 969 AOI22_X2
* cell instance $47926 r0 *1 428.26,60.2
X$47926 1438 1326 25 44 1285 NOR2_X2
* cell instance $47927 m0 *1 430.73,60.2
X$47927 1293 1437 44 25 1540 AND2_X1
* cell instance $47928 m0 *1 428.26,60.2
X$47928 25 1555 1122 1293 1437 44 AOI21_X4
* cell instance $47931 r0 *1 429.21,60.2
X$47931 1326 1540 25 44 1582 NOR2_X1
* cell instance $47933 m0 *1 435.1,60.2
X$47933 1436 1539 1441 25 1440 44 AOI21_X1
* cell instance $47936 m0 *1 438.9,60.2
X$47936 1479 25 44 1496 INV_X1
* cell instance $47937 m0 *1 439.28,60.2
X$47937 1496 1287 25 44 1557 OR2_X1
* cell instance $47942 r0 *1 438.9,60.2
X$47942 1445 1479 1562 25 44 1561 NAND3_X1
* cell instance $47945 m0 *1 444.03,60.2
X$47945 1481 1483 1083 25 44 1492 NAND3_X1
* cell instance $47946 m0 *1 442.7,60.2
X$47946 1529 1482 1483 25 44 1391 NAND3_X2
* cell instance $47950 m0 *1 447.26,60.2
X$47950 1485 1484 25 44 1525 OR2_X1
* cell instance $47951 m0 *1 448.02,60.2
X$47951 1484 1485 25 44 1536 NAND2_X1
* cell instance $47952 m0 *1 448.59,60.2
X$47952 1485 1484 25 44 1526 XNOR2_X2
* cell instance $47954 r0 *1 444.22,60.2
X$47954 1537 25 44 1495 BUF_X2
* cell instance $47955 r0 *1 444.98,60.2
X$47955 1575 1445 1479 1537 25 44 1610 AOI22_X2
* cell instance $47958 r0 *1 447.64,60.2
X$47958 1658 1525 1536 44 1575 25 OAI21_X1
* cell instance $47960 r0 *1 448.59,60.2
X$47960 25 1574 1526 1485 1479 1084 44 OAI22_X4
* cell instance $47962 m0 *1 451.06,60.2
X$47962 1451 1494 1483 1480 44 25 1446 OAI22_X1
* cell instance $47963 m0 *1 452.01,60.2
X$47963 1480 1482 25 44 1494 NAND2_X1
* cell instance $47964 m0 *1 452.58,60.2
X$47964 1483 1480 1393 1333 44 25 1531 OAI22_X2
* cell instance $47965 m0 *1 454.29,60.2
X$47965 1448 1451 1447 1491 44 1533 25 NOR4_X2
* cell instance $47966 m0 *1 456,60.2
X$47966 1486 1333 1492 25 1448 44 AOI21_X2
* cell instance $47968 m0 *1 457.52,60.2
X$47968 1490 1449 25 44 1486 NAND2_X1
* cell instance $47971 m0 *1 459.04,60.2
X$47971 1486 1333 25 44 1487 NOR2_X1
* cell instance $47972 m0 *1 459.61,60.2
X$47972 1487 1451 1447 25 44 1489 NOR3_X1
* cell instance $47973 m0 *1 460.37,60.2
X$47973 1231 1488 1489 44 25 1484 OAI21_X2
* cell instance $47980 r0 *1 453.34,60.2
X$47980 1783 1441 25 44 1393 NOR2_X1
* cell instance $47981 r0 *1 453.91,60.2
X$47981 25 1573 1533 1439 1563 44 AOI21_X4
* cell instance $47982 r0 *1 456.38,60.2
X$47982 1491 1448 25 44 1569 NOR2_X1
* cell instance $47983 r0 *1 456.95,60.2
X$47983 1564 1568 1531 25 1532 44 AOI21_X1
* cell instance $47984 r0 *1 457.71,60.2
X$47984 1527 1528 25 44 1491 NAND2_X1
* cell instance $47985 r0 *1 458.28,60.2
X$47985 1486 1528 25 44 1565 NOR2_X1
* cell instance $47987 r0 *1 459.23,60.2
X$47987 1566 25 44 1527 INV_X1
* cell instance $47990 r0 *1 460.18,60.2
X$47990 1530 1482 1529 25 1488 44 AOI21_X1
* cell instance $48284 r0 *1 340.29,65.8
X$48284 1542 1586 25 44 1738 NOR2_X2
* cell instance $48286 m0 *1 340.48,65.8
X$48286 25 1588 1628 1542 1669 1586 44 OAI22_X4
* cell instance $48287 r0 *1 341.24,65.8
X$48287 1586 1236 44 25 1739 AND2_X1
* cell instance $48289 r0 *1 342.38,65.8
X$48289 1092 1585 25 44 1741 NOR2_X2
* cell instance $48291 m0 *1 344.28,65.8
X$48291 1047 1508 25 44 1632 XNOR2_X2
* cell instance $48294 m0 *1 346.94,65.8
X$48294 25 1455 1242 1201 1589 1586 44 OAI22_X4
* cell instance $48295 m0 *1 350.17,65.8
X$48295 1590 1109 1508 25 1796 44 NAND3_X4
* cell instance $48296 m0 *1 352.64,65.8
X$48296 25 1694 1346 1546 1668 44 AOI21_X4
* cell instance $48298 m0 *1 355.87,65.8
X$48298 25 1109 1594 1507 1534 1674 44 NAND4_X4
* cell instance $48299 m0 *1 359.29,65.8
X$48299 25 1310 1593 1507 1534 1637 44 NAND4_X4
* cell instance $48300 m0 *1 362.71,65.8
X$48300 1634 1675 1595 44 25 1734 MUX2_X2
* cell instance $48301 m0 *1 364.42,65.8
X$48301 1676 1595 1675 25 1698 44 AOI21_X1
* cell instance $48305 m0 *1 367.65,65.8
X$48305 1635 1636 1697 44 1823 25 OAI21_X1
* cell instance $48306 m0 *1 368.41,65.8
X$48306 1678 1313 1581 25 44 1697 NOR3_X1
* cell instance $48307 m0 *1 369.17,65.8
X$48307 1680 1638 1637 25 1732 44 AOI21_X2
* cell instance $48308 m0 *1 370.5,65.8
X$48308 1686 1207 1512 25 44 1680 NAND3_X1
* cell instance $48310 m0 *1 372.02,65.8
X$48310 1696 1639 1682 1732 44 25 1699 AND4_X1
* cell instance $48311 m0 *1 373.16,65.8
X$48311 1700 1734 1682 25 1733 44 AOI21_X2
* cell instance $48312 m0 *1 374.49,65.8
X$48312 1698 1640 1641 44 1683 25 OAI21_X1
* cell instance $48315 m0 *1 376.2,65.8
X$48315 1700 1520 1599 25 1786 44 AOI21_X2
* cell instance $48321 r0 *1 347.51,65.8
X$48321 1201 1586 1242 1455 1630 1744 25 44 OAI221_X2
* cell instance $48325 r0 *1 350.93,65.8
X$48325 1734 1693 1744 25 44 1782 NAND3_X2
* cell instance $48326 r0 *1 352.26,65.8
X$48326 1693 1744 25 1695 44 NAND2_X4
* cell instance $48328 r0 *1 354.16,65.8
X$48328 25 1109 1695 1669 1745 1682 44 NOR4_X4
* cell instance $48330 r0 *1 358.34,65.8
X$48330 1507 1534 1109 1594 44 25 1746 AND4_X1
* cell instance $48336 r0 *1 365.94,65.8
X$48336 25 1752 1635 1636 1757 1728 44 NOR4_X4
* cell instance $48337 r0 *1 369.36,65.8
X$48337 25 1682 1732 1696 1639 1800 44 NAND4_X4
* cell instance $48340 r0 *1 373.73,65.8
X$48340 25 1755 1786 1752 1733 44 AOI21_X4
* cell instance $48342 r0 *1 377.72,65.8
X$48342 1701 1380 1756 25 44 1787 NOR3_X1
* cell instance $48343 r0 *1 378.48,65.8
X$48343 1787 1788 1758 44 1924 25 OAI21_X1
* cell instance $48346 r0 *1 379.81,65.8
X$48346 1702 1696 1790 25 1788 44 AOI21_X1
* cell instance $48349 r0 *1 381.14,65.8
X$48349 1703 1790 1683 1754 1829 25 44 OAI211_X2
* cell instance $48350 m0 *1 382.66,65.8
X$48350 1426 1704 1641 44 1703 25 OAI21_X1
* cell instance $48355 m0 *1 391.21,65.8
X$48355 25 1642 1736 1643 1685 1737 44 NOR4_X4
* cell instance $48356 m0 *1 394.63,65.8
X$48356 1642 1736 1643 1685 25 44 1735 OR4_X1
* cell instance $48358 m0 *1 396.53,65.8
X$48358 1431 1645 44 25 1793 AND2_X1
* cell instance $48359 m0 *1 397.29,65.8
X$48359 1705 1645 1646 25 1729 44 AOI21_X1
* cell instance $48360 m0 *1 398.05,65.8
X$48360 763 877 25 44 1705 NOR2_X1
* cell instance $48361 m0 *1 398.62,65.8
X$48361 1731 1647 25 44 1648 XNOR2_X2
* cell instance $48363 m0 *1 400.71,65.8
X$48363 1385 1729 1100 44 1730 25 OAI21_X1
* cell instance $48367 r0 *1 382.85,65.8
X$48367 1754 1683 1703 44 1804 25 OAI21_X1
* cell instance $48371 r0 *1 390.83,65.8
X$48371 1552 1510 25 44 1762 NAND2_X2
* cell instance $48372 r0 *1 391.78,65.8
X$48372 1644 1762 44 25 1763 XNOR2_X1
* cell instance $48373 r0 *1 392.92,65.8
X$48373 1763 1648 25 44 1758 NOR2_X2
* cell instance $48374 r0 *1 393.87,65.8
X$48374 1759 1648 1793 44 25 1685 AND3_X1
* cell instance $48377 r0 *1 397.1,65.8
X$48377 1793 1646 1705 1431 25 44 1764 AOI22_X2
* cell instance $48380 r0 *1 399.38,65.8
X$48380 1414 25 44 1731 INV_X1
* cell instance $48382 r0 *1 399.95,65.8
X$48382 1648 1730 44 25 1926 XNOR2_X1
* cell instance $48385 m0 *1 404.13,65.8
X$48385 1254 1364 1501 25 1678 44 NAND3_X4
* cell instance $48387 m0 *1 409.83,65.8
X$48387 1649 633 1690 25 44 1689 MUX2_X1
* cell instance $48388 m0 *1 411.16,65.8
X$48388 1556 1560 25 44 1690 OR2_X1
* cell instance $48397 r0 *1 417.43,65.8
X$48397 1706 1431 1766 25 1650 44 AOI21_X2
* cell instance $48398 r0 *1 418.76,65.8
X$48398 1766 1706 1431 25 44 1477 NAND3_X2
* cell instance $48400 r0 *1 420.28,65.8
X$48400 1767 1651 25 44 1766 XNOR2_X2
* cell instance $48402 m0 *1 420.66,65.8
X$48402 1651 1767 44 1604 25 XOR2_X2
* cell instance $48405 r0 *1 422.56,65.8
X$48405 1171 25 44 1706 INV_X2
* cell instance $48408 m0 *1 423.51,65.8
X$48408 1653 1708 1556 25 44 NOR2_X4
* cell instance $48410 m0 *1 429.02,65.8
X$48410 1654 25 44 1769 INV_X1
* cell instance $48411 m0 *1 429.4,65.8
X$48411 1654 1655 1824 25 44 1367 OR3_X2
* cell instance $48413 m0 *1 432.06,65.8
X$48413 1483 1439 1084 44 1727 25 OAI21_X1
* cell instance $48415 m0 *1 433.58,65.8
X$48415 1725 1656 1684 25 44 1726 NOR3_X1
* cell instance $48417 r0 *1 423.89,65.8
X$48417 1808 1707 25 44 1767 NOR2_X2
* cell instance $48418 r0 *1 424.84,65.8
X$48418 725 680 25 44 1707 NOR2_X1
* cell instance $48422 r0 *1 428.07,65.8
X$48422 1706 1794 44 25 1652 XNOR2_X1
* cell instance $48426 r0 *1 430.54,65.8
X$48426 1441 680 1727 44 1794 25 OAI21_X1
* cell instance $48429 r0 *1 432.44,65.8
X$48429 1084 1439 25 44 1768 NOR2_X2
* cell instance $48432 m0 *1 434.72,65.8
X$48432 1791 1614 1612 1900 44 1606 25 NOR4_X2
* cell instance $48433 m0 *1 437.95,65.8
X$48433 1710 1612 25 44 1679 NAND2_X1
* cell instance $48434 m0 *1 436.81,65.8
X$48434 1709 1679 44 25 1725 XNOR2_X1
* cell instance $48437 m0 *1 438.9,65.8
X$48437 1710 1562 25 44 1615 NAND2_X1
* cell instance $48440 m0 *1 443.46,65.8
X$48440 1712 1616 1677 25 44 1710 MUX2_X1
* cell instance $48441 m0 *1 444.79,65.8
X$48441 1659 1714 1712 44 1677 25 OAI21_X1
* cell instance $48442 m0 *1 445.55,65.8
X$48442 1714 1671 1723 1617 1722 1715 25 44 1537 OAI33_X1
* cell instance $48443 m0 *1 446.88,65.8
X$48443 1716 1712 1673 25 44 1672 NAND3_X1
* cell instance $48447 m0 *1 456.95,65.8
X$48447 1721 1717 1568 25 1660 44 AOI21_X1
* cell instance $48450 m0 *1 458.66,65.8
X$48450 1449 1618 44 25 1665 AND2_X1
* cell instance $48452 m0 *1 460.18,65.8
X$48452 1566 1665 44 25 1662 XNOR2_X1
* cell instance $48453 m0 *1 461.32,65.8
X$48453 1780 25 44 1661 INV_X1
* cell instance $48461 r0 *1 440.61,65.8
X$48461 1724 1711 25 44 1771 NOR2_X1
* cell instance $48462 r0 *1 441.18,65.8
X$48462 1772 1711 1785 44 1709 25 OAI21_X1
* cell instance $48463 r0 *1 441.94,65.8
X$48463 1785 1617 25 44 1724 NAND2_X1
* cell instance $48465 r0 *1 443.27,65.8
X$48465 1774 1714 25 44 1785 NOR2_X1
* cell instance $48466 r0 *1 443.84,65.8
X$48466 1573 1716 1712 25 44 1711 NAND3_X1
* cell instance $48467 r0 *1 444.6,65.8
X$48467 1713 1482 25 44 1774 NOR2_X1
* cell instance $48468 r0 *1 445.17,65.8
X$48468 1673 25 44 1714 INV_X1
* cell instance $48469 r0 *1 445.55,65.8
X$48469 1482 1713 1712 25 1723 44 AOI21_X1
* cell instance $48470 r0 *1 446.31,65.8
X$48470 1482 1713 1673 44 1715 25 OAI21_X1
* cell instance $48474 r0 *1 450.68,65.8
X$48474 1776 44 1441 25 BUF_X4
* cell instance $48478 r0 *1 454.48,65.8
X$48478 1490 1783 1776 1395 25 44 1721 NOR4_X1
* cell instance $48479 r0 *1 455.43,65.8
X$48479 1718 1817 25 44 1130 XNOR2_X2
* cell instance $48480 r0 *1 457.33,65.8
X$48480 1718 1449 25 44 1568 NOR2_X2
* cell instance $48482 r0 *1 458.66,65.8
X$48482 1781 1719 1566 44 1620 25 OAI21_X1
* cell instance $48483 r0 *1 459.42,65.8
X$48483 1718 1528 25 44 1720 NAND2_X1
* cell instance $48484 r0 *1 459.99,65.8
X$48484 1720 1665 1779 1777 44 25 1781 OAI22_X1
* cell instance $48761 m0 *1 340.29,68.6
X$48761 25 1740 1738 1507 1739 44 AOI21_X4
* cell instance $48782 r0 *1 341.05,68.6
X$48782 1629 1738 1507 1739 1873 44 25 AOI211_X2
* cell instance $48785 r0 *1 344.47,68.6
X$48785 1630 1587 25 44 1864 OR2_X2
* cell instance $48786 r0 *1 345.42,68.6
X$48786 25 1833 1630 1109 1508 44 AOI21_X4
* cell instance $48788 m0 *1 346.18,68.6
X$48788 1587 1741 1346 25 1742 44 AOI21_X2
* cell instance $48790 m0 *1 348.46,68.6
X$48790 1346 1741 25 44 1743 NAND2_X2
* cell instance $48793 r0 *1 347.89,68.6
X$48793 25 1421 1743 1796 1818 44 NOR3_X4
* cell instance $48796 m0 *1 351.31,68.6
X$48796 1744 1693 1734 44 25 1919 AND3_X1
* cell instance $48798 m0 *1 353.4,68.6
X$48798 1346 1421 1578 25 1745 44 NAND3_X4
* cell instance $48799 m0 *1 352.64,68.6
X$48799 1744 1693 44 25 1819 AND2_X1
* cell instance $48801 m0 *1 356.06,68.6
X$48801 1109 1695 1669 1745 44 1640 25 OR4_X2
* cell instance $48804 m0 *1 359.1,68.6
X$48804 1750 1592 1748 1633 1674 1749 44 25 AOI221_X2
* cell instance $48805 m0 *1 361.19,68.6
X$48805 25 1747 1748 1592 1750 44 AOI21_X4
* cell instance $48806 m0 *1 363.66,68.6
X$48806 1639 1798 1634 1749 25 1751 44 NAND4_X2
* cell instance $48811 r0 *1 353.4,68.6
X$48811 25 1782 1669 1745 1797 44 NOR3_X4
* cell instance $48812 r0 *1 356.06,68.6
X$48812 1594 1109 25 44 1866 NAND2_X1
* cell instance $48814 r0 *1 357.39,68.6
X$48814 1823 1640 1834 1835 1820 1753 25 44 OAI221_X2
* cell instance $48818 r0 *1 361.57,68.6
X$48818 1836 1797 25 44 1821 OR2_X1
* cell instance $48819 r0 *1 362.33,68.6
X$48819 25 1867 1821 1876 1751 1754 44 AOI22_X4
* cell instance $48822 m0 *1 367.46,68.6
X$48822 25 1753 1784 1799 1637 1638 44 AOI22_X4
* cell instance $48827 r0 *1 368.22,68.6
X$48827 1797 1798 1047 25 44 1826 NAND3_X1
* cell instance $48828 r0 *1 368.98,68.6
X$48828 1047 1797 44 25 1922 AND2_X1
* cell instance $48829 r0 *1 369.74,68.6
X$48829 1752 1756 1784 1826 1800 1803 25 44 OAI221_X2
* cell instance $48831 m0 *1 374.3,68.6
X$48831 1696 44 1798 25 BUF_X4
* cell instance $48832 m0 *1 372.59,68.6
X$48832 1699 1754 1801 25 44 NOR2_X4
* cell instance $48834 m0 *1 376.58,68.6
X$48834 1380 1879 1756 1701 44 1828 25 NOR4_X2
* cell instance $48835 m0 *1 376.01,68.6
X$48835 1380 1599 25 44 1908 NAND2_X1
* cell instance $48836 m0 *1 378.29,68.6
X$48836 1704 1922 1757 25 1789 44 AOI21_X2
* cell instance $48837 m0 *1 379.62,68.6
X$48837 25 1759 1758 1760 1789 1801 44 AOI22_X4
* cell instance $48840 m0 *1 383.8,68.6
X$48840 1599 1758 1759 44 25 1761 MUX2_X2
* cell instance $48846 r0 *1 380,68.6
X$48846 1802 1551 1598 25 1790 44 AOI21_X2
* cell instance $48847 r0 *1 381.33,68.6
X$48847 1702 1760 1803 1829 44 2056 25 NOR4_X2
* cell instance $48848 r0 *1 383.04,68.6
X$48848 1702 1803 1790 25 1805 44 AOI21_X1
* cell instance $48849 r0 *1 383.8,68.6
X$48849 1829 1803 25 44 1830 NOR2_X1
* cell instance $48850 r0 *1 384.37,68.6
X$48850 1828 1805 1761 1830 1993 44 25 AOI211_X2
* cell instance $48851 r0 *1 386.08,68.6
X$48851 1805 1828 25 44 1840 OR2_X1
* cell instance $48855 m0 *1 392.16,68.6
X$48855 25 1554 1759 1648 1762 1642 44 NOR4_X4
* cell instance $48860 r0 *1 392.35,68.6
X$48860 1552 1554 1414 25 1806 44 AOI21_X1
* cell instance $48864 m0 *1 397.48,68.6
X$48864 1602 1764 25 44 1831 XNOR2_X2
* cell instance $48868 r0 *1 398.24,68.6
X$48868 1552 44 1765 25 BUF_X4
* cell instance $48870 m0 *1 401.47,68.6
X$48870 1436 1602 25 44 1927 NAND2_X2
* cell instance $48874 m0 *1 405.65,68.6
X$48874 1644 1765 1436 25 44 NOR2_X4
* cell instance $48877 m0 *1 409.64,68.6
X$48877 1765 44 1539 25 BUF_X4
* cell instance $48881 m0 *1 416.29,68.6
X$48881 1426 44 1081 25 BUF_X4
* cell instance $48887 r0 *1 403.37,68.6
X$48887 1415 1461 25 1802 44 NAND2_X4
* cell instance $48891 r0 *1 406.41,68.6
X$48891 1554 1385 25 1807 44 NAND2_X4
* cell instance $48892 r0 *1 408.12,68.6
X$48892 1554 1765 25 44 1891 NOR2_X2
* cell instance $48897 m0 *1 424.08,68.6
X$48897 1795 1441 25 44 1708 NOR2_X2
* cell instance $48898 m0 *1 423.32,68.6
X$48898 1768 1539 1707 25 1795 44 AOI21_X1
* cell instance $48900 m0 *1 425.22,68.6
X$48900 680 725 25 44 1809 XNOR2_X2
* cell instance $48905 r0 *1 424.08,68.6
X$48905 1768 1441 25 44 1808 NOR2_X1
* cell instance $48907 r0 *1 425.41,68.6
X$48907 1441 1539 25 44 1827 NAND2_X1
* cell instance $48908 r0 *1 425.98,68.6
X$48908 25 1827 1809 1768 1653 1807 44 OAI22_X4
* cell instance $48910 m0 *1 428.26,68.6
X$48910 1933 991 1769 1825 25 846 44 NAND4_X2
* cell instance $48912 m0 *1 431.68,68.6
X$48912 1483 1431 25 44 1770 NAND2_X1
* cell instance $48913 m0 *1 432.25,68.6
X$48913 1171 1770 25 44 1792 OR2_X1
* cell instance $48914 m0 *1 433.01,68.6
X$48914 680 1792 1822 44 1226 25 OAI21_X1
* cell instance $48915 m0 *1 433.77,68.6
X$48915 1706 1447 25 44 1810 NOR2_X1
* cell instance $48917 m0 *1 435.1,68.6
X$48917 1439 25 44 680 INV_X4
* cell instance $48923 r0 *1 432.63,68.6
X$48923 1770 1171 1891 1529 1810 25 44 1822 AOI221_X1
* cell instance $48927 m0 *1 440.23,68.6
X$48927 1771 1773 1711 25 44 1791 MUX2_X1
* cell instance $48928 m0 *1 441.75,68.6
X$48928 1773 1617 25 44 1772 NOR2_X1
* cell instance $48931 m0 *1 444.6,68.6
X$48931 1657 1712 1773 25 44 1722 MUX2_X1
* cell instance $48935 r0 *1 440.61,68.6
X$48935 1392 1775 25 44 1852 NOR2_X1
* cell instance $48936 r0 *1 441.18,68.6
X$48936 1392 1811 25 44 1171 XNOR2_X2
* cell instance $48940 r0 *1 445.55,68.6
X$48940 1775 1862 25 44 1399 XNOR2_X2
* cell instance $48942 r0 *1 448.97,68.6
X$48942 1861 1812 44 1776 25 XOR2_X2
* cell instance $48943 r0 *1 450.68,68.6
X$48943 25 1498 1775 1392 1854 44 NOR3_X4
* cell instance $48945 m0 *1 450.87,68.6
X$48945 1498 1775 1392 25 44 1783 OR3_X2
* cell instance $48947 m0 *1 454.29,68.6
X$48947 1395 1783 1776 44 25 1777 OAI21_X2
* cell instance $48951 m0 *1 458.09,68.6
X$48951 1395 1618 25 44 1814 OR2_X1
* cell instance $48953 m0 *1 459.04,68.6
X$48953 1490 1779 25 44 1816 NAND2_X1
* cell instance $48959 r0 *1 455.43,68.6
X$48959 1395 1529 1855 25 1817 44 AOI21_X2
* cell instance $48961 r0 *1 457.52,68.6
X$48961 1854 1483 1395 25 44 1813 NAND3_X1
* cell instance $48963 r0 *1 458.66,68.6
X$48963 1816 1813 1814 25 1719 44 AOI21_X1
* cell instance $48966 r0 *1 460.37,68.6
X$48966 1856 1815 25 44 1663 NOR2_X1
* cell instance $48967 m0 *1 461.32,68.6
X$48967 1780 1815 25 44 1231 OR2_X2
* cell instance $48968 m0 *1 460.75,68.6
X$48968 1778 1779 25 44 1780 NOR2_X1
* cell instance $49250 m0 *1 345.42,71.4
X$49250 25 1421 1201 1833 1874 44 NOR3_X4
* cell instance $49251 m0 *1 348.08,71.4
X$49251 1201 1510 1833 44 25 1832 OAI21_X2
* cell instance $49252 m0 *1 349.41,71.4
X$49252 1510 1743 1796 25 44 1860 OR3_X2
* cell instance $49272 r0 *1 344.66,71.4
X$49272 1109 1508 25 44 1918 XNOR2_X2
* cell instance $49276 r0 *1 347.89,71.4
X$49276 1381 1833 1743 44 25 1897 OAI21_X4
* cell instance $49277 r0 *1 350.36,71.4
X$49277 1873 1897 25 44 1835 NAND2_X2
* cell instance $49278 m0 *1 351.12,71.4
X$49278 25 1796 1587 1306 1839 44 NOR3_X4
* cell instance $49280 m0 *1 353.78,71.4
X$49280 1306 1864 1866 44 1899 25 NOR3_X2
* cell instance $49285 r0 *1 352.26,71.4
X$49285 1874 1694 1667 1782 1834 44 25 AOI211_X2
* cell instance $49287 m0 *1 356.44,71.4
X$49287 1373 1818 25 44 1820 NOR2_X2
* cell instance $49292 m0 *1 357.77,71.4
X$49292 1820 1835 1834 44 25 1754 OAI21_X4
* cell instance $49295 r0 *1 357.96,71.4
X$49295 1109 1381 1508 25 1875 44 AOI21_X2
* cell instance $49300 m0 *1 361.57,71.4
X$49300 1797 1836 25 44 1837 NOR2_X2
* cell instance $49302 m0 *1 362.52,71.4
X$49302 1749 1639 1798 25 44 1867 NAND3_X2
* cell instance $49303 m0 *1 363.85,71.4
X$49303 1901 1623 1838 44 25 1921 OAI21_X4
* cell instance $49306 m0 *1 368.6,71.4
X$49306 1797 1047 25 44 2009 NAND2_X2
* cell instance $49307 m0 *1 369.55,71.4
X$49307 1639 1798 1747 25 1757 44 NAND3_X4
* cell instance $49311 r0 *1 361.57,71.4
X$49311 1746 1875 25 44 1836 NOR2_X1
* cell instance $49312 r0 *1 362.14,71.4
X$49312 1875 1746 1838 1623 1901 1903 25 44 OAI221_X2
* cell instance $49315 r0 *1 364.8,71.4
X$49315 1903 1877 1756 44 1902 25 NOR3_X2
* cell instance $49319 r0 *1 367.46,71.4
X$49319 1907 1625 25 44 1901 NOR2_X2
* cell instance $49322 r0 *1 370.12,71.4
X$49322 1878 44 1877 25 BUF_X4
* cell instance $49327 r0 *1 376.58,71.4
X$49327 1798 1520 25 44 1923 NAND2_X2
* cell instance $49329 m0 *1 380.19,71.4
X$49329 1598 1551 25 44 1925 NAND2_X1
* cell instance $49331 m0 *1 380.76,71.4
X$49331 1598 1551 1804 1803 1520 1970 44 25 AOI221_X2
* cell instance $49333 m0 *1 383.04,71.4
X$49333 1804 1520 1803 25 1910 44 AOI21_X1
* cell instance $49335 m0 *1 384.56,71.4
X$49335 1842 1761 1830 44 25 1872 AND3_X1
* cell instance $49337 m0 *1 386.27,71.4
X$49337 1840 1872 25 44 1912 XNOR2_X2
* cell instance $49343 m0 *1 390.07,71.4
X$49343 1818 1510 877 25 1841 44 AOI21_X2
* cell instance $49344 m0 *1 391.59,71.4
X$49344 1841 1842 1554 1552 25 44 1913 NAND4_X1
* cell instance $49345 m0 *1 392.54,71.4
X$49345 1385 1644 1842 1841 25 44 1914 OR4_X1
* cell instance $49346 m0 *1 393.68,71.4
X$49346 1841 763 1644 25 44 1881 NAND3_X1
* cell instance $49348 m0 *1 394.63,71.4
X$49348 1554 763 1841 25 44 1915 OR3_X1
* cell instance $49349 m0 *1 395.58,71.4
X$49349 1842 1841 44 25 1843 XNOR2_X1
* cell instance $49350 m0 *1 396.72,71.4
X$49350 1843 1385 25 44 1871 NOR2_X2
* cell instance $49353 r0 *1 393.11,71.4
X$49353 1806 1880 25 44 2062 NOR2_X1
* cell instance $49354 r0 *1 393.68,71.4
X$49354 1881 1913 1914 1915 25 44 1880 NAND4_X1
* cell instance $49357 m0 *1 398.24,71.4
X$49357 1644 1871 25 44 1844 XNOR2_X2
* cell instance $49360 m0 *1 400.33,71.4
X$49360 1844 1884 1885 44 25 1870 OAI21_X2
* cell instance $49361 m0 *1 401.66,71.4
X$49361 25 1845 1474 1917 1870 44 AOI21_X4
* cell instance $49366 r0 *1 399,71.4
X$49366 1554 1871 25 44 1882 XNOR2_X2
* cell instance $49367 r0 *1 400.9,71.4
X$49367 1882 1765 25 44 1958 NAND2_X1
* cell instance $49368 r0 *1 401.47,71.4
X$49368 1883 757 1957 25 44 1847 MUX2_X1
* cell instance $49369 r0 *1 402.8,71.4
X$49369 1885 1884 25 44 1917 NAND2_X1
* cell instance $49372 r0 *1 405.08,71.4
X$49372 1831 1845 25 44 1887 XNOR2_X2
* cell instance $49374 m0 *1 406.03,71.4
X$49374 1845 1831 44 1846 25 XOR2_X2
* cell instance $49376 m0 *1 408.69,71.4
X$49376 1847 1807 25 44 1886 NAND2_X2
* cell instance $49378 m0 *1 409.83,71.4
X$49378 1807 1847 44 25 1869 AND2_X1
* cell instance $49379 m0 *1 410.59,71.4
X$49379 1869 25 44 1848 CLKBUF_X3
* cell instance $49381 m0 *1 411.73,71.4
X$49381 1886 1386 25 44 1916 NOR2_X1
* cell instance $49383 r0 *1 406.98,71.4
X$49383 1887 1474 25 44 1954 NOR2_X1
* cell instance $49385 r0 *1 407.93,71.4
X$49385 1954 1928 1891 1474 1731 25 44 1953 AOI221_X1
* cell instance $49389 r0 *1 411.73,71.4
X$49389 1916 639 1888 25 44 2136 MUX2_X1
* cell instance $49390 m0 *1 412.87,71.4
X$49390 1847 1386 25 44 1888 NOR2_X1
* cell instance $49394 m0 *1 418,71.4
X$49394 1846 1848 25 44 1890 NAND2_X1
* cell instance $49400 m0 *1 433.2,71.4
X$49400 1868 1849 25 44 1824 NAND2_X1
* cell instance $49403 r0 *1 413.25,71.4
X$49403 1887 1886 25 44 1889 NAND2_X1
* cell instance $49404 r0 *1 413.82,71.4
X$49404 1889 1911 1887 25 44 1905 MUX2_X1
* cell instance $49405 r0 *1 415.15,71.4
X$49405 1932 1951 25 44 1911 NOR2_X1
* cell instance $49407 r0 *1 415.91,71.4
X$49407 1887 1431 25 44 1930 NOR2_X1
* cell instance $49409 r0 *1 416.67,71.4
X$49409 1846 1848 1474 44 1931 25 NOR3_X2
* cell instance $49411 r0 *1 418.19,71.4
X$49411 1890 1909 1846 25 44 1906 MUX2_X1
* cell instance $49412 r0 *1 419.52,71.4
X$49412 1846 1474 25 44 1950 NOR2_X1
* cell instance $49413 r0 *1 420.09,71.4
X$49413 1081 1905 1906 25 1947 44 AOI21_X2
* cell instance $49415 r0 *1 422.18,71.4
X$49415 1891 25 44 1973 INV_X1
* cell instance $49417 r0 *1 425.6,71.4
X$49417 1386 1892 1807 44 1904 25 OAI21_X1
* cell instance $49421 r0 *1 433.39,71.4
X$49421 1892 1904 1893 44 25 1812 MUX2_X2
* cell instance $49422 m0 *1 434.34,71.4
X$49422 1975 1580 25 44 1900 NAND2_X1
* cell instance $49424 m0 *1 434.91,71.4
X$49424 1946 1849 1580 1868 44 25 1443 AND4_X2
* cell instance $49431 r0 *1 436.43,71.4
X$49431 1893 1892 1431 25 44 1934 NAND3_X1
* cell instance $49433 m0 *1 440.04,71.4
X$49433 1392 1850 44 25 1851 AND2_X1
* cell instance $49434 m0 *1 438.9,71.4
X$49434 1863 1775 25 44 1850 XOR2_X1
* cell instance $49435 m0 *1 440.8,71.4
X$49435 1851 1811 1852 25 44 1481 MUX2_X1
* cell instance $49436 m0 *1 442.13,71.4
X$49436 1865 2038 1617 1573 25 1849 44 NAND4_X2
* cell instance $49439 r0 *1 440.61,71.4
X$49439 1812 1898 1431 25 44 1811 NAND3_X2
* cell instance $49442 r0 *1 443.65,71.4
X$49442 1451 1447 1853 44 1935 25 OAI21_X1
* cell instance $49443 m0 *1 444.41,71.4
X$49443 1529 1853 25 44 1713 NAND2_X1
* cell instance $49447 m0 *1 446.31,71.4
X$49447 1863 552 25 44 1862 NOR2_X1
* cell instance $49448 m0 *1 445.36,71.4
X$49448 1673 1712 1716 44 25 1865 AND3_X1
* cell instance $49451 m0 *1 450.68,71.4
X$49451 1859 44 1483 25 BUF_X4
* cell instance $49452 m0 *1 448.78,71.4
X$49452 1812 1861 25 44 1859 XNOR2_X2
* cell instance $49458 r0 *1 452.39,71.4
X$49458 1894 1857 25 44 1943 NOR2_X1
* cell instance $49461 m0 *1 455.62,71.4
X$49461 1857 1855 1718 1717 1395 1778 44 25 AOI221_X2
* cell instance $49462 m0 *1 454.67,71.4
X$49462 1854 1859 25 44 1717 NAND2_X2
* cell instance $49463 m0 *1 457.71,71.4
X$49463 1449 1854 1483 25 1895 44 AOI21_X2
* cell instance $49464 m0 *1 459.04,71.4
X$49464 1718 1528 1858 1895 44 1815 25 NOR4_X2
* cell instance $49465 m0 *1 460.75,71.4
X$49465 1778 1779 1858 1857 1856 44 25 AOI211_X2
* cell instance $49470 r0 *1 454.86,71.4
X$49470 1190 2117 1896 44 25 1176 OAI21_X2
* cell instance $49471 r0 *1 456.19,71.4
X$49471 1395 1940 1717 25 1896 44 AOI21_X1
* cell instance $49474 r0 *1 457.52,71.4
X$49474 1618 1483 1395 25 44 1939 NAND3_X2
* cell instance $49771 m0 *1 344.47,74.2
X$49771 25 1864 1918 1572 2005 1742 44 OAI22_X4
* cell instance $49777 r0 *1 348.46,74.2
X$49777 1818 1373 25 44 2003 OR2_X2
* cell instance $49778 m0 *1 349.03,74.2
X$49778 1373 1818 1873 1897 1984 44 25 AOI211_X2
* cell instance $49780 m0 *1 350.74,74.2
X$49780 1874 1694 2006 25 44 NOR2_X4
* cell instance $49781 m0 *1 352.45,74.2
X$49781 25 1596 1694 1874 1695 1960 44 NOR4_X4
* cell instance $49784 r0 *1 349.41,74.2
X$49784 1897 1873 44 25 1983 AND2_X1
* cell instance $49786 r0 *1 350.93,74.2
X$49786 1578 1897 25 1959 44 NAND2_X4
* cell instance $49790 r0 *1 354.73,74.2
X$49790 1819 1984 1983 1920 25 44 2051 AOI22_X1
* cell instance $49791 r0 *1 355.68,74.2
X$49791 1695 1373 1818 25 44 1986 NOR3_X1
* cell instance $49792 r0 *1 356.44,74.2
X$49792 1986 1834 1961 1920 2003 2082 44 25 AOI221_X2
* cell instance $49793 m0 *1 357.2,74.2
X$49793 1695 1674 1633 25 1961 44 AOI21_X1
* cell instance $49795 m0 *1 357.96,74.2
X$49795 1746 1875 1819 44 1920 25 NOR3_X2
* cell instance $49797 m0 *1 359.48,74.2
X$49797 1674 1633 25 44 2007 NAND2_X2
* cell instance $49802 m0 *1 364.04,74.2
X$49802 25 1596 1756 1877 1903 1945 44 NOR4_X4
* cell instance $49803 m0 *1 360.81,74.2
X$49803 25 1902 1837 1945 2094 1752 44 OAI22_X4
* cell instance $49809 r0 *1 363.47,74.2
X$49809 1623 1838 25 44 2010 NOR2_X2
* cell instance $49810 r0 *1 364.42,74.2
X$49810 25 1596 1756 1877 1921 2039 44 NOR4_X4
* cell instance $49812 m0 *1 368.79,74.2
X$49812 25 1756 1877 1921 1784 44 NOR3_X4
* cell instance $49814 m0 *1 371.45,74.2
X$49814 1921 1922 1757 25 1962 44 AOI21_X1
* cell instance $49815 m0 *1 372.21,74.2
X$49815 1922 1757 25 44 1989 NAND2_X1
* cell instance $49816 m0 *1 372.78,74.2
X$49816 1907 1878 1756 44 1990 25 NOR3_X2
* cell instance $49821 r0 *1 370.5,74.2
X$49821 1878 1756 25 44 2042 NOR2_X2
* cell instance $49822 r0 *1 371.45,74.2
X$49822 25 1989 2011 1990 2054 1921 44 OAI22_X4
* cell instance $49824 m0 *1 377.72,74.2
X$49824 1461 1925 1798 44 25 1963 AND3_X1
* cell instance $49825 m0 *1 375.25,74.2
X$49825 1755 877 1923 44 25 1965 OAI21_X4
* cell instance $49826 m0 *1 378.67,74.2
X$49826 1925 1922 1757 25 1991 44 AOI21_X1
* cell instance $49828 m0 *1 385.51,74.2
X$49828 1956 1910 1842 25 44 2058 NAND3_X2
* cell instance $49829 m0 *1 386.84,74.2
X$49829 1761 1520 25 44 1968 NAND2_X1
* cell instance $49830 m0 *1 387.41,74.2
X$49830 1760 1426 25 44 1956 NOR2_X1
* cell instance $49835 r0 *1 375.63,74.2
X$49835 1925 1755 1879 1923 2085 25 44 OAI211_X2
* cell instance $49837 r0 *1 378.1,74.2
X$49837 1925 1461 1798 25 1964 44 AOI21_X1
* cell instance $49838 r0 *1 378.86,74.2
X$49838 1963 1759 1964 1801 1991 1966 44 25 AOI221_X2
* cell instance $49842 r0 *1 383.61,74.2
X$49842 1761 1966 1520 1965 25 2106 44 NAND4_X2
* cell instance $49843 r0 *1 385.32,74.2
X$49843 1760 763 1498 1965 44 1967 25 NOR4_X2
* cell instance $49845 r0 *1 387.22,74.2
X$49845 1956 1965 1842 1966 25 44 1995 NAND4_X1
* cell instance $49846 r0 *1 388.17,74.2
X$49846 763 1968 1970 44 1969 25 OAI21_X1
* cell instance $49849 r0 *1 392.35,74.2
X$49849 1626 1364 25 1907 44 NAND2_X4
* cell instance $49852 m0 *1 400.71,74.2
X$49852 1882 1884 1958 25 44 1957 MUX2_X1
* cell instance $49858 m0 *1 407.17,74.2
X$49858 1953 1955 25 44 2001 NAND2_X1
* cell instance $49860 m0 *1 407.74,74.2
X$49860 1954 1929 1952 25 44 1955 NAND3_X1
* cell instance $49861 m0 *1 408.5,74.2
X$49861 25 1971 1928 1952 1929 44 AOI21_X4
* cell instance $49867 r0 *1 409.45,74.2
X$49867 2001 2070 1807 2002 1974 44 25 AOI211_X2
* cell instance $49868 r0 *1 411.16,74.2
X$49868 2139 1971 1846 25 2002 44 AOI21_X1
* cell instance $49870 m0 *1 416.86,74.2
X$49870 1971 1846 1930 1931 1951 1948 44 25 AOI221_X2
* cell instance $49872 m0 *1 418.95,74.2
X$49872 1950 1909 2020 1931 1932 1949 44 25 AOI221_X2
* cell instance $49876 m0 *1 434.72,74.2
X$49876 1944 25 44 1946 INV_X1
* cell instance $49878 m0 *1 436.62,74.2
X$49878 1976 1934 25 44 1392 XNOR2_X2
* cell instance $49883 m0 *1 444.03,74.2
X$49883 1977 1935 1936 1451 25 44 1659 AOI22_X2
* cell instance $49884 m0 *1 445.74,74.2
X$49884 25 1392 1857 1944 1937 1987 44 NOR4_X4
* cell instance $49885 m0 *1 449.16,74.2
X$49885 1392 1857 1944 1937 44 1938 25 OR4_X2
* cell instance $49887 r0 *1 418,74.2
X$49887 2021 1971 1999 2000 1972 25 44 OAI211_X2
* cell instance $49891 r0 *1 421.04,74.2
X$49891 1973 1998 1972 1996 44 25 1997 AND4_X1
* cell instance $49892 r0 *1 422.18,74.2
X$49892 25 1972 1996 1973 1998 2043 44 NAND4_X4
* cell instance $49893 r0 *1 425.6,74.2
X$49893 1997 25 44 1892 CLKBUF_X3
* cell instance $49896 r0 *1 428.83,74.2
X$49896 1949 1948 44 25 1976 AND2_X2
* cell instance $49898 r0 *1 432.82,74.2
X$49898 1975 1994 44 25 1868 AND2_X1
* cell instance $49901 r0 *1 434.15,74.2
X$49901 1975 1992 1849 2025 25 44 1656 NAND4_X1
* cell instance $49905 r0 *1 437.57,74.2
X$49905 1992 1977 1853 25 44 2040 NAND3_X1
* cell instance $49909 r0 *1 443.65,74.2
X$49909 1977 1978 25 44 1979 NOR2_X1
* cell instance $49911 r0 *1 444.41,74.2
X$49911 1977 1988 25 44 1773 XNOR2_X2
* cell instance $49913 r0 *1 446.69,74.2
X$49913 2026 1978 1858 1529 1988 44 25 AOI211_X2
* cell instance $49917 r0 *1 449.73,74.2
X$49917 25 1858 1980 1982 1987 44 AOI21_X4
* cell instance $49918 m0 *1 451.06,74.2
X$49918 1980 1943 1941 44 25 1712 OAI21_X4
* cell instance $49920 m0 *1 453.53,74.2
X$49920 1855 1939 1938 44 25 1447 OAI21_X4
* cell instance $49921 m0 *1 456,74.2
X$49921 1939 1938 1855 1857 1942 44 25 1940 OAI221_X1
* cell instance $49922 m0 *1 457.14,74.2
X$49922 1528 1941 1718 25 1942 44 AOI21_X1
* cell instance $49927 r0 *1 453.34,74.2
X$49927 1985 1483 1618 44 25 1982 AND3_X1
* cell instance $49928 r0 *1 454.29,74.2
X$49928 1985 44 1395 25 BUF_X4
* cell instance $49931 r0 *1 458.85,74.2
X$49931 25 1451 1857 1981 1779 44 AOI21_X4
* cell instance $49932 m0 *1 459.23,74.2
X$49932 1941 1718 1895 44 25 1981 OAI21_X2
* cell instance $49982 r0 *1 461.32,74.2
X$49982 1858 1857 1981 44 25 2032 OAI21_X2
* cell instance $50234 r0 *1 334.59,51.8
X$50234 25 1266 1140 1195 1057 44 AOI21_X4
* cell instance $50236 r0 *1 337.82,51.8
X$50236 1014 44 1268 25 BUF_X4
* cell instance $50237 m0 *1 338.39,51.8
X$50237 1107 1058 44 25 1196 XNOR2_X1
* cell instance $50239 m0 *1 339.53,51.8
X$50239 1291 1199 1196 44 25 1263 AND3_X1
* cell instance $50241 m0 *1 340.67,51.8
X$50241 1200 1264 25 44 1197 NAND2_X1
* cell instance $50242 m0 *1 341.24,51.8
X$50242 1200 1110 25 44 1265 NAND2_X1
* cell instance $50243 m0 *1 341.81,51.8
X$50243 1091 1292 834 44 1199 25 NOR3_X2
* cell instance $50244 m0 *1 343.14,51.8
X$50244 834 1091 1292 44 25 1344 OAI21_X2
* cell instance $50246 m0 *1 345.23,51.8
X$50246 25 1201 1143 1199 1305 44 AOI21_X4
* cell instance $50249 m0 *1 349.41,51.8
X$50249 25 1242 1202 1203 1296 44 AOI21_X4
* cell instance $50253 r0 *1 339.15,51.8
X$50253 1014 1266 25 44 1291 NAND2_X2
* cell instance $50254 r0 *1 340.1,51.8
X$50254 25 1306 1263 1059 1265 44 AOI21_X4
* cell instance $50256 r0 *1 342.95,51.8
X$50256 1091 1107 25 44 1267 NOR2_X2
* cell instance $50257 r0 *1 343.9,51.8
X$50257 1344 1238 1295 44 25 1346 OAI21_X4
* cell instance $50258 r0 *1 346.37,51.8
X$50258 1107 1268 1266 25 44 1305 NAND3_X2
* cell instance $50260 r0 *1 348.08,51.8
X$50260 1266 1268 1107 44 25 1295 AND3_X2
* cell instance $50262 r0 *1 349.6,51.8
X$50262 1268 1146 25 44 1202 NAND2_X2
* cell instance $50263 r0 *1 350.55,51.8
X$50263 1307 1134 1141 25 44 1350 NAND3_X2
* cell instance $50266 r0 *1 355.68,51.8
X$50266 25 958 959 1150 1269 1264 44 NOR4_X4
* cell instance $50267 r0 *1 359.1,51.8
X$50267 957 1353 25 44 1309 XNOR2_X2
* cell instance $50268 m0 *1 360.62,51.8
X$50268 25 1148 1112 1018 1149 1353 44 NAND4_X4
* cell instance $50269 m0 *1 359.86,51.8
X$50269 1248 1149 957 25 44 1244 NAND3_X1
* cell instance $50271 m0 *1 364.23,51.8
X$50271 1019 1151 25 44 1466 XNOR2_X2
* cell instance $50272 m0 *1 366.13,51.8
X$50272 25 1205 1206 1313 1139 1151 44 AOI22_X4
* cell instance $50276 r0 *1 361.57,51.8
X$50276 25 1148 1311 957 1149 1292 44 NAND4_X4
* cell instance $50278 r0 *1 366.51,51.8
X$50278 1315 1111 1269 25 44 1206 MUX2_X1
* cell instance $50419 m0 *1 321.86,35
X$50419 727 25 44 467 BUF_X2
* cell instance $50440 r0 *1 322.62,35
X$50440 786 44 158 25 BUF_X4
* cell instance $50443 r0 *1 326.23,35
X$50443 25 682 768 821 791 820 44 FA_X1
* cell instance $50444 m0 *1 326.99,35
X$50444 513 158 44 25 791 AND2_X1
* cell instance $50448 m0 *1 334.59,35
X$50448 733 25 44 799 BUF_X2
* cell instance $50454 r0 *1 330.41,35
X$50454 821 621 796 44 25 822 HA_X1
* cell instance $50458 r0 *1 337.25,35
X$50458 769 799 648 25 864 44 AOI21_X2
* cell instance $50464 r0 *1 340.86,35
X$50464 650 799 25 44 739 NAND2_X2
* cell instance $50469 r0 *1 344.66,35
X$50469 740 770 829 25 44 900 NAND3_X2
* cell instance $50470 m0 *1 345.04,35
X$50470 644 738 704 25 44 740 NAND3_X1
* cell instance $50472 m0 *1 345.8,35
X$50472 704 644 25 44 770 OR2_X1
* cell instance $50473 m0 *1 346.56,35
X$50473 650 25 44 704 INV_X1
* cell instance $50477 m0 *1 350.93,35
X$50477 25 800 745 793 742 746 747 44 AOI221_X4
* cell instance $50480 r0 *1 345.99,35
X$50480 830 804 801 25 44 829 MUX2_X1
* cell instance $50481 r0 *1 347.32,35
X$50481 644 771 704 25 44 830 NAND3_X1
* cell instance $50482 r0 *1 348.08,35
X$50482 573 527 44 25 802 AND2_X1
* cell instance $50485 r0 *1 353.4,35
X$50485 527 573 650 625 25 44 805 NAND4_X1
* cell instance $50486 r0 *1 354.35,35
X$50486 805 771 774 708 793 44 25 AOI211_X2
* cell instance $50488 m0 *1 354.54,35
X$50488 578 705 794 44 25 806 MUX2_X2
* cell instance $50490 m0 *1 357.96,35
X$50490 508 579 44 25 706 AND2_X1
* cell instance $50491 m0 *1 358.72,35
X$50491 749 608 752 753 44 25 707 AND4_X2
* cell instance $50492 m0 *1 360.05,35
X$50492 706 709 625 581 25 44 752 NAND4_X1
* cell instance $50500 r0 *1 358.91,35
X$50500 772 773 25 44 794 NAND2_X1
* cell instance $50501 r0 *1 359.48,35
X$50501 772 706 773 25 44 753 NAND3_X1
* cell instance $50506 r0 *1 362.14,35
X$50506 25 1049 651 773 772 44 AOI21_X4
* cell instance $50509 r0 *1 365.56,35
X$50509 581 792 44 25 772 AND2_X2
* cell instance $50511 r0 *1 366.7,35
X$50511 708 774 44 25 775 AND2_X1
* cell instance $50512 r0 *1 367.46,35
X$50512 775 709 625 44 25 961 MUX2_X2
* cell instance $50513 m0 *1 368.22,35
X$50513 625 710 25 44 809 NAND2_X1
* cell instance $50514 m0 *1 368.79,35
X$50514 710 776 625 44 25 792 AND3_X2
* cell instance $50515 m0 *1 369.93,35
X$50515 656 25 44 709 INV_X1
* cell instance $50520 m0 *1 375.82,35
X$50520 656 828 777 789 745 25 44 OAI211_X2
* cell instance $50521 m0 *1 377.53,35
X$50521 758 25 44 778 BUF_X2
* cell instance $50525 r0 *1 369.17,35
X$50525 25 625 709 773 962 44 NOR3_X4
* cell instance $50527 r0 *1 372.02,35
X$50527 710 658 776 44 25 774 OAI21_X2
* cell instance $50531 r0 *1 375.44,35
X$50531 828 789 777 44 25 773 OAI21_X4
* cell instance $50532 r0 *1 377.91,35
X$50532 25 828 778 779 787 44 AOI21_X4
* cell instance $50534 m0 *1 381.14,35
X$50534 711 712 788 44 25 780 HA_X1
* cell instance $50538 m0 *1 384.75,35
X$50538 713 25 44 785 INV_X1
* cell instance $50540 m0 *1 388.17,35
X$50540 714 25 44 784 INV_X1
* cell instance $50543 m0 *1 390.26,35
X$50543 760 759 862 44 25 823 HA_X1
* cell instance $50547 r0 *1 381.33,35
X$50547 788 25 44 810 CLKBUF_X3
* cell instance $50549 r0 *1 382.66,35
X$50549 780 25 44 787 BUF_X2
* cell instance $50552 r0 *1 385.7,35
X$50552 785 824 811 44 25 825 HA_X1
* cell instance $50555 r0 *1 388.74,35
X$50555 784 823 781 44 25 824 HA_X1
* cell instance $50557 m0 *1 393.49,35
X$50557 715 761 783 44 25 782 HA_X1
* cell instance $50561 m0 *1 398.62,35
X$50561 57 764 718 44 25 766 HA_X1
* cell instance $50565 r0 *1 394.25,35
X$50565 783 716 876 44 25 860 HA_X1
* cell instance $50570 m0 *1 401.28,35
X$50570 766 25 44 719 INV_X1
* cell instance $50571 m0 *1 400.9,35
X$50571 718 25 44 767 INV_X1
* cell instance $50574 m0 *1 402.04,35
X$50574 755 756 720 25 664 44 AOI21_X1
* cell instance $50575 m0 *1 402.99,35
X$50575 54 757 720 44 25 755 HA_X1
* cell instance $50581 m0 *1 410.02,35
X$50581 818 25 44 635 INV_X1
* cell instance $50585 m0 *1 411.73,35
X$50585 723 25 44 743 INV_X1
* cell instance $50875 r0 *1 324.14,32.2
X$50875 406 158 44 25 730 AND2_X1
* cell instance $50876 m0 *1 324.71,32.2
X$50876 467 189 44 25 703 AND2_X1
* cell instance $50880 r0 *1 324.9,32.2
X$50880 730 703 637 44 25 790 HA_X1
* cell instance $50881 m0 *1 326.8,32.2
X$50881 25 646 682 640 683 637 44 FA_X1
* cell instance $50885 m0 *1 330.79,32.2
X$50885 25 570 621 732 571 640 44 FA_X1
* cell instance $50890 r0 *1 334.4,32.2
X$50890 732 734 733 44 25 769 HA_X1
* cell instance $50892 m0 *1 334.97,32.2
X$50892 684 25 44 734 INV_X1
* cell instance $50897 m0 *1 339.91,32.2
X$50897 689 641 647 44 25 648 HA_X1
* cell instance $50898 m0 *1 339.53,32.2
X$50898 686 25 44 689 INV_X1
* cell instance $50901 m0 *1 345.04,32.2
X$50901 648 650 540 25 692 44 AOI21_X1
* cell instance $50903 m0 *1 346.56,32.2
X$50903 691 645 622 44 25 643 OAI21_X2
* cell instance $50907 m0 *1 351.88,32.2
X$50907 577 623 25 44 748 NAND2_X1
* cell instance $50908 m0 *1 352.45,32.2
X$50908 649 623 577 25 747 44 AOI21_X1
* cell instance $50909 m0 *1 353.21,32.2
X$50909 573 650 25 44 649 NAND2_X1
* cell instance $50910 m0 *1 353.78,32.2
X$50910 573 695 578 651 25 44 694 AOI22_X2
* cell instance $50911 m0 *1 355.49,32.2
X$50911 563 608 25 44 696 NAND2_X1
* cell instance $50916 r0 *1 340.29,32.2
X$50916 647 25 44 650 BUF_X2
* cell instance $50920 r0 *1 345.23,32.2
X$50920 739 738 644 25 691 44 AOI21_X1
* cell instance $50921 r0 *1 345.99,32.2
X$50921 527 573 25 44 738 NAND2_X1
* cell instance $50924 r0 *1 348.46,32.2
X$50924 692 25 44 742 INV_X1
* cell instance $50929 r0 *1 351.69,32.2
X$50929 573 748 693 696 694 955 25 44 OAI221_X2
* cell instance $50930 r0 *1 353.78,32.2
X$50930 573 706 25 44 693 OR2_X1
* cell instance $50932 r0 *1 354.73,32.2
X$50932 651 696 573 25 44 705 NOR3_X1
* cell instance $50934 r0 *1 356.25,32.2
X$50934 608 563 653 652 746 25 44 OAI211_X2
* cell instance $50935 r0 *1 357.96,32.2
X$50935 579 508 25 44 652 NAND2_X1
* cell instance $50936 r0 *1 358.53,32.2
X$50936 652 653 25 44 749 OR2_X1
* cell instance $50939 m0 *1 360.24,32.2
X$50939 579 610 25 44 654 NAND2_X1
* cell instance $50941 m0 *1 364.61,32.2
X$50941 625 581 25 44 655 NAND2_X1
* cell instance $50947 r0 *1 363.47,32.2
X$50947 653 656 655 44 25 651 OAI21_X4
* cell instance $50948 m0 *1 365.75,32.2
X$50948 25 808 626 625 657 44 AOI21_X4
* cell instance $50954 r0 *1 367.08,32.2
X$50954 657 25 44 708 INV_X1
* cell instance $50956 m0 *1 369.55,32.2
X$50956 627 25 44 710 CLKBUF_X3
* cell instance $50959 m0 *1 373.54,32.2
X$50959 700 25 44 776 CLKBUF_X3
* cell instance $50963 r0 *1 371.45,32.2
X$50963 25 656 657 710 658 44 AOI21_X4
* cell instance $50966 m0 *1 374.87,32.2
X$50966 583 44 658 25 BUF_X4
* cell instance $50968 m0 *1 376.58,32.2
X$50968 584 44 779 25 BUF_X4
* cell instance $50972 r0 *1 380.95,32.2
X$50972 659 25 44 711 INV_X1
* cell instance $50973 m0 *1 381.52,32.2
X$50973 25 701 660 713 702 476 44 FA_X1
* cell instance $50975 m0 *1 384.56,32.2
X$50975 25 661 701 714 628 441 44 FA_X1
* cell instance $50979 r0 *1 381.33,32.2
X$50979 660 25 44 712 INV_X1
* cell instance $50982 m0 *1 390.45,32.2
X$50982 629 25 44 760 INV_X1
* cell instance $50989 r0 *1 392.73,32.2
X$50989 762 352 840 44 25 716 HA_X1
* cell instance $50991 m0 *1 393.49,32.2
X$50991 27 186 44 25 715 AND2_X1
* cell instance $50993 m0 *1 394.63,32.2
X$50993 587 25 44 662 INV_X1
* cell instance $50997 m0 *1 405.08,32.2
X$50997 699 630 25 44 631 NOR2_X1
* cell instance $50998 m0 *1 405.65,32.2
X$50998 592 25 44 665 INV_X1
* cell instance $50999 m0 *1 406.03,32.2
X$50999 132 639 592 44 25 754 HA_X1
* cell instance $51000 m0 *1 407.93,32.2
X$51000 632 25 44 698 INV_X1
* cell instance $51005 r0 *1 398.43,32.2
X$51005 160 763 663 44 25 717 HA_X1
* cell instance $51006 r0 *1 400.33,32.2
X$51006 717 663 765 25 589 44 AOI21_X1
* cell instance $51007 r0 *1 401.09,32.2
X$51007 767 664 719 44 765 25 OAI21_X1
* cell instance $51009 r0 *1 402.23,32.2
X$51009 722 720 718 663 25 44 699 NAND4_X1
* cell instance $51013 r0 *1 405.27,32.2
X$51013 665 666 721 44 756 25 OAI21_X1
* cell instance $51014 r0 *1 406.03,32.2
X$51014 754 25 44 721 INV_X1
* cell instance $51015 r0 *1 406.41,32.2
X$51015 697 722 698 25 666 44 AOI21_X1
* cell instance $51016 r0 *1 407.17,32.2
X$51016 168 729 722 44 25 697 HA_X1
* cell instance $51018 r0 *1 409.83,32.2
X$51018 397 751 667 44 25 723 HA_X1
* cell instance $51019 m0 *1 412.68,32.2
X$51019 376 635 668 44 25 690 HA_X1
* cell instance $51020 m0 *1 411.73,32.2
X$51020 593 631 685 44 25 636 AND3_X1
* cell instance $51021 m0 *1 414.58,32.2
X$51021 690 335 668 25 669 44 AOI21_X1
* cell instance $51022 m0 *1 415.34,32.2
X$51022 688 634 25 44 687 NAND2_X1
* cell instance $51024 m0 *1 421.99,32.2
X$51024 480 633 681 44 25 672 HA_X1
* cell instance $51025 m0 *1 423.89,32.2
X$51025 334 680 674 44 25 677 HA_X1
* cell instance $51026 m0 *1 425.79,32.2
X$51026 677 674 678 25 634 44 AOI21_X1
* cell instance $51027 m0 *1 426.55,32.2
X$51027 675 25 44 676 INV_X1
* cell instance $51083 r0 *1 411.73,32.2
X$51083 667 668 670 636 25 744 44 NAND4_X2
* cell instance $51084 r0 *1 413.44,32.2
X$51084 667 25 44 741 INV_X1
* cell instance $51086 r0 *1 414.01,32.2
X$51086 741 669 743 44 736 25 OAI21_X1
* cell instance $51088 r0 *1 414.96,32.2
X$51088 735 670 736 25 688 44 AOI21_X1
* cell instance $51089 r0 *1 415.72,32.2
X$51089 478 737 670 44 25 735 HA_X1
* cell instance $51092 r0 *1 419.9,32.2
X$51092 671 634 25 44 685 NAND2_X1
* cell instance $51094 r0 *1 421.99,32.2
X$51094 418 731 673 44 25 728 HA_X1
* cell instance $51095 r0 *1 423.89,32.2
X$51095 728 672 673 25 679 44 AOI21_X1
* cell instance $51097 r0 *1 424.84,32.2
X$51097 681 673 675 674 25 44 671 NAND4_X1
* cell instance $51099 r0 *1 425.98,32.2
X$51099 676 679 726 44 678 25 OAI21_X1
* cell instance $51100 r0 *1 426.74,32.2
X$51100 396 725 675 44 25 724 HA_X1
* cell instance $51101 r0 *1 428.64,32.2
X$51101 724 25 44 726 INV_X1
* cell instance $51372 m0 *1 328.51,29.4
X$51372 502 25 44 646 INV_X1
* cell instance $51379 m0 *1 331.74,29.4
X$51379 537 25 44 570 INV_X1
* cell instance $51383 m0 *1 335.35,29.4
X$51383 539 25 44 572 INV_X1
* cell instance $51388 r0 *1 331.55,29.4
X$51388 513 60 44 25 571 AND2_X1
* cell instance $51393 r0 *1 336.68,29.4
X$51393 25 603 684 686 559 572 44 FA_X1
* cell instance $51399 r0 *1 340.29,29.4
X$51399 606 25 44 641 INV_X1
* cell instance $51402 m0 *1 344.66,29.4
X$51402 604 44 573 25 BUF_X4
* cell instance $51407 r0 *1 345.61,29.4
X$51407 25 644 540 573 541 44 AOI21_X4
* cell instance $51408 r0 *1 348.08,29.4
X$51408 574 644 25 44 622 NAND2_X1
* cell instance $51410 r0 *1 349.03,29.4
X$51410 574 576 575 44 25 804 OAI21_X4
* cell instance $51411 r0 *1 351.5,29.4
X$51411 575 576 25 44 645 NOR2_X1
* cell instance $51414 m0 *1 352.45,29.4
X$51414 528 508 25 44 576 NAND2_X2
* cell instance $51415 r0 *1 352.83,29.4
X$51415 541 25 44 623 INV_X1
* cell instance $51416 r0 *1 353.21,29.4
X$51416 542 623 577 25 578 44 AOI21_X2
* cell instance $51418 m0 *1 353.78,29.4
X$51418 573 579 508 25 44 542 NAND3_X1
* cell instance $51420 r0 *1 354.54,29.4
X$51420 623 577 608 563 25 44 695 AOI22_X1
* cell instance $51423 m0 *1 355.68,29.4
X$51423 25 608 509 508 510 44 AOI21_X4
* cell instance $51425 m0 *1 359.1,29.4
X$51425 25 575 510 579 580 44 AOI21_X4
* cell instance $51426 m0 *1 361.57,29.4
X$51426 612 25 44 581 CLKBUF_X3
* cell instance $51431 r0 *1 357.39,29.4
X$51431 508 25 44 610 INV_X1
* cell instance $51432 r0 *1 357.77,29.4
X$51432 610 579 510 25 44 611 OR3_X1
* cell instance $51433 r0 *1 358.72,29.4
X$51433 611 508 575 44 25 750 OAI21_X2
* cell instance $51435 r0 *1 360.24,29.4
X$51435 580 510 610 25 44 624 NOR3_X1
* cell instance $51440 r0 *1 362.52,29.4
X$51440 25 653 580 581 626 44 AOI21_X4
* cell instance $51443 m0 *1 366.89,29.4
X$51443 614 543 615 44 25 626 HA_X1
* cell instance $51448 r0 *1 367.65,29.4
X$51448 615 44 625 25 BUF_X4
* cell instance $51450 r0 *1 369.74,29.4
X$51450 582 567 627 44 25 657 HA_X1
* cell instance $51451 m0 *1 370.12,29.4
X$51451 616 25 44 582 INV_X1
* cell instance $51457 m0 *1 373.35,29.4
X$51457 545 569 700 44 25 583 HA_X1
* cell instance $51460 m0 *1 378.29,29.4
X$51460 513 291 44 25 617 AND2_X1
* cell instance $51462 m0 *1 382.09,29.4
X$51462 301 323 25 44 702 NAND2_X1
* cell instance $51465 m0 *1 385.89,29.4
X$51465 467 301 44 25 548 AND2_X1
* cell instance $51466 m0 *1 386.65,29.4
X$51466 549 548 619 44 25 585 HA_X1
* cell instance $51468 m0 *1 388.74,29.4
X$51468 619 25 44 620 INV_X1
* cell instance $51473 r0 *1 375.82,29.4
X$51473 547 642 584 44 25 758 HA_X1
* cell instance $51474 r0 *1 377.72,29.4
X$51474 25 475 642 659 617 369 44 FA_X1
* cell instance $51476 r0 *1 386.84,29.4
X$51476 585 25 44 628 INV_X1
* cell instance $51477 r0 *1 387.22,29.4
X$51477 25 354 661 629 620 515 44 FA_X1
* cell instance $51479 r0 *1 390.64,29.4
X$51479 586 25 44 759 INV_X1
* cell instance $51481 m0 *1 391.21,29.4
X$51481 25 561 586 587 618 353 44 FA_X1
* cell instance $51488 m0 *1 395.58,29.4
X$51488 406 513 44 25 613 AND2_X1
* cell instance $51494 r0 *1 400.14,29.4
X$51494 590 589 443 609 591 638 25 44 OAI221_X2
* cell instance $51495 m0 *1 400.9,29.4
X$51495 244 613 443 25 593 44 AOI21_X1
* cell instance $51496 m0 *1 400.52,29.4
X$51496 588 25 44 590 INV_X1
* cell instance $51497 m0 *1 401.66,29.4
X$51497 558 25 44 591 INV_X1
* cell instance $51505 r0 *1 405.08,29.4
X$51505 607 595 592 588 25 44 630 NAND4_X1
* cell instance $51507 m0 *1 406.41,29.4
X$51507 196 552 607 44 25 594 HA_X1
* cell instance $51511 m0 *1 409.26,29.4
X$51511 229 551 595 44 25 605 HA_X1
* cell instance $51516 m0 *1 419.71,29.4
X$51516 601 195 25 44 600 NOR2_X1
* cell instance $51517 m0 *1 420.28,29.4
X$51517 597 550 44 25 601 XNOR2_X1
* cell instance $51531 r0 *1 408.31,29.4
X$51531 605 594 595 25 632 44 AOI21_X1
* cell instance $51535 r0 *1 411.54,29.4
X$51535 687 636 228 593 638 25 44 602 AOI221_X1
* cell instance $51538 r0 *1 413.63,29.4
X$51538 602 596 44 25 599 AND2_X1
* cell instance $51541 r0 *1 418.19,29.4
X$51541 25 30 600 43 597 418 44 DFFR_X2
* cell instance $51544 r0 *1 423.32,29.4
X$51544 25 30 599 43 2894 598 44 DFFR_X2
* cell instance $51799 m0 *1 318.06,37.8
X$51799 819 25 44 406 BUF_X2
* cell instance $51816 m0 *1 325.47,37.8
X$51816 406 189 44 25 795 AND2_X1
* cell instance $51818 m0 *1 326.23,37.8
X$51818 790 795 820 44 25 831 HA_X1
* cell instance $51820 m0 *1 331.17,37.8
X$51820 796 25 44 797 BUF_X2
* cell instance $51822 m0 *1 332.12,37.8
X$51822 822 25 44 798 CLKBUF_X2
* cell instance $51826 m0 *1 333.26,37.8
X$51826 798 797 769 25 853 44 AOI21_X1
* cell instance $51827 m0 *1 334.21,37.8
X$51827 798 797 827 25 832 44 AOI21_X1
* cell instance $51829 m0 *1 335.16,37.8
X$51829 799 769 25 44 827 OR2_X1
* cell instance $51831 m0 *1 337.44,37.8
X$51831 800 799 44 834 25 XOR2_X2
* cell instance $51834 r0 *1 334.4,37.8
X$51834 832 853 800 44 25 833 MUX2_X2
* cell instance $51839 r0 *1 338.96,37.8
X$51839 643 864 25 44 934 NAND2_X1
* cell instance $51841 m0 *1 339.72,37.8
X$51841 799 800 25 44 835 XNOR2_X2
* cell instance $51845 m0 *1 346.37,37.8
X$51845 802 803 25 44 836 NAND2_X1
* cell instance $51846 m0 *1 346.94,37.8
X$51846 802 650 25 44 801 NAND2_X1
* cell instance $51847 m0 *1 347.51,37.8
X$51847 644 704 25 44 857 NAND2_X1
* cell instance $51848 m0 *1 348.08,37.8
X$51848 802 803 650 25 44 856 NAND3_X2
* cell instance $51851 m0 *1 353.21,37.8
X$51851 508 581 528 579 44 25 803 AND4_X2
* cell instance $51852 m0 *1 354.54,37.8
X$51852 528 581 508 579 25 771 44 NAND4_X2
* cell instance $51860 r0 *1 346.18,37.8
X$51860 25 807 866 804 857 954 44 NOR4_X4
* cell instance $51867 r0 *1 361.38,37.8
X$51867 807 581 25 44 868 NAND2_X2
* cell instance $51871 r0 *1 363.66,37.8
X$51871 808 837 44 25 889 AND2_X2
* cell instance $51872 r0 *1 364.61,37.8
X$51872 837 808 838 25 44 869 NAND3_X2
* cell instance $51873 m0 *1 365.18,37.8
X$51873 581 25 44 838 INV_X1
* cell instance $51876 m0 *1 365.75,37.8
X$51876 808 839 809 44 25 807 OAI21_X4
* cell instance $51877 m0 *1 368.22,37.8
X$51877 809 839 25 44 837 OR2_X1
* cell instance $51880 r0 *1 365.94,37.8
X$51880 838 808 837 44 25 888 AND3_X1
* cell instance $51883 m0 *1 372.4,37.8
X$51883 658 776 778 25 839 44 AOI21_X2
* cell instance $51885 m0 *1 381.33,37.8
X$51885 25 810 779 863 777 826 44 OAI211_X4
* cell instance $51887 r0 *1 372.97,37.8
X$51887 710 776 25 44 872 OR2_X1
* cell instance $51888 r0 *1 373.73,37.8
X$51888 778 658 710 44 906 25 NOR3_X2
* cell instance $51891 m0 *1 385.13,37.8
X$51891 811 44 826 25 BUF_X4
* cell instance $51895 m0 *1 387.41,37.8
X$51895 825 44 863 25 BUF_X4
* cell instance $51904 r0 *1 392.35,37.8
X$51904 862 859 950 44 25 874 HA_X1
* cell instance $51905 r0 *1 394.25,37.8
X$51905 861 860 875 44 25 887 HA_X1
* cell instance $51907 m0 *1 394.44,37.8
X$51907 662 782 861 44 25 859 HA_X1
* cell instance $51913 m0 *1 401.47,37.8
X$51913 25 947 858 27 201 44 AOI21_X4
* cell instance $51919 r0 *1 401.66,37.8
X$51919 840 914 25 44 858 NAND2_X1
* cell instance $51924 r0 *1 407.36,37.8
X$51924 878 25 44 751 INV_X4
* cell instance $51925 m0 *1 408.88,37.8
X$51925 814 815 813 812 816 25 44 OAI211_X2
* cell instance $51926 m0 *1 408.12,37.8
X$51926 812 813 814 44 818 25 OAI21_X1
* cell instance $51928 r0 *1 408.31,37.8
X$51928 841 842 814 25 44 855 NOR3_X1
* cell instance $51929 r0 *1 409.07,37.8
X$51929 855 842 841 25 886 44 AOI21_X1
* cell instance $51930 r0 *1 409.83,37.8
X$51930 818 817 843 854 844 816 25 44 849 OAI33_X1
* cell instance $51931 m0 *1 411.16,37.8
X$51931 815 817 25 44 852 NAND2_X1
* cell instance $51933 m0 *1 411.73,37.8
X$51933 817 815 25 44 851 OR2_X1
* cell instance $51990 r0 *1 411.16,37.8
X$51990 844 854 852 851 850 44 25 AOI211_X2
* cell instance $51991 r0 *1 412.87,37.8
X$51991 847 886 849 850 596 25 44 OAI211_X2
* cell instance $51996 r0 *1 422.75,37.8
X$51996 848 885 846 25 44 847 NOR3_X1
* cell instance $51998 r0 *1 424.27,37.8
X$51998 882 992 25 44 845 NAND2_X1
* cell instance $52000 r0 *1 425.03,37.8
X$52000 884 883 845 25 885 44 AOI21_X1
* cell instance $52257 m0 *1 334.4,46.2
X$52257 25 1005 898 1013 1057 44 NOR3_X4
* cell instance $52259 m0 *1 338.77,46.2
X$52259 1015 1016 25 44 1058 NAND2_X1
* cell instance $52260 m0 *1 339.34,46.2
X$52260 835 1016 1015 25 1059 44 AOI21_X2
* cell instance $52264 m0 *1 343.14,46.2
X$52264 896 1017 835 44 1090 25 OAI21_X1
* cell instance $52270 r0 *1 335.35,46.2
X$52270 1040 1088 1134 25 44 NOR2_X4
* cell instance $52273 r0 *1 338.01,46.2
X$52273 1042 834 896 1017 1136 25 44 OAI211_X2
* cell instance $52275 r0 *1 341.24,46.2
X$52275 1017 834 896 25 44 1106 NOR3_X1
* cell instance $52277 r0 *1 342.38,46.2
X$52277 1107 1091 1090 896 1017 1093 25 44 1092 OAI33_X1
* cell instance $52279 r0 *1 345.23,46.2
X$52279 834 1042 1060 1111 25 44 1093 NOR4_X1
* cell instance $52281 m0 *1 348.84,46.2
X$52281 977 1018 1046 25 1091 44 NAND3_X4
* cell instance $52282 m0 *1 351.31,46.2
X$52282 977 1018 25 1061 44 NAND2_X4
* cell instance $52285 m0 *1 362.14,46.2
X$52285 579 1049 25 44 1062 XNOR2_X2
* cell instance $52290 r0 *1 350.74,46.2
X$52290 1060 1137 25 44 1109 XNOR2_X2
* cell instance $52291 r0 *1 352.64,46.2
X$52291 1110 1018 25 44 1137 NAND2_X2
* cell instance $52300 r0 *1 365.37,46.2
X$52300 1062 1018 25 44 1139 NOR2_X2
* cell instance $52301 r0 *1 366.32,46.2
X$52301 1063 1062 904 25 1150 44 NAND3_X4
* cell instance $52303 m0 *1 371.45,46.2
X$52303 773 776 44 1209 25 XOR2_X2
* cell instance $52307 m0 *1 374.87,46.2
X$52307 776 773 25 44 1152 XNOR2_X2
* cell instance $52309 m0 *1 377.53,46.2
X$52309 909 908 25 44 942 NOR2_X2
* cell instance $52315 m0 *1 394.63,46.2
X$52315 840 876 2897 44 25 1066 HA_X1
* cell instance $52321 r0 *1 378.29,46.2
X$52321 1064 942 25 44 1158 NOR2_X2
* cell instance $52322 r0 *1 379.24,46.2
X$52322 810 1098 25 44 1153 XNOR2_X2
* cell instance $52323 r0 *1 381.14,46.2
X$52323 1098 810 44 1155 25 XOR2_X2
* cell instance $52329 r0 *1 394.44,46.2
X$52329 1065 840 876 25 1159 44 NAND3_X4
* cell instance $52330 r0 *1 396.91,46.2
X$52330 840 876 1067 44 25 1358 HA_X1
* cell instance $52334 r0 *1 401.28,46.2
X$52334 915 981 1100 25 44 1068 NOR3_X1
* cell instance $52335 m0 *1 401.66,46.2
X$52335 1067 25 44 914 INV_X1
* cell instance $52339 r0 *1 402.04,46.2
X$52339 1116 1068 982 44 1102 25 OAI21_X1
* cell instance $52340 r0 *1 402.8,46.2
X$52340 1067 1069 1102 25 1071 44 AOI21_X1
* cell instance $52342 m0 *1 404.7,46.2
X$52342 1022 25 44 1070 INV_X1
* cell instance $52343 m0 *1 403.94,46.2
X$52343 1025 1022 981 25 44 1024 NAND3_X1
* cell instance $52345 m0 *1 405.27,46.2
X$52345 1025 1023 983 25 1104 44 AOI21_X1
* cell instance $52347 m0 *1 406.79,46.2
X$52347 1104 879 916 25 44 1072 NAND3_X1
* cell instance $52351 r0 *1 404.7,46.2
X$52351 751 1070 1105 44 985 25 OAI21_X1
* cell instance $52354 r0 *1 406.41,46.2
X$52354 1025 25 44 1105 INV_X1
* cell instance $52355 r0 *1 406.79,46.2
X$52355 1071 1117 1072 25 854 44 AOI21_X2
* cell instance $52358 r0 *1 408.69,46.2
X$52358 1097 1103 1118 44 1117 25 OAI21_X1
* cell instance $52360 m0 *1 409.64,46.2
X$52360 1074 1073 1101 44 25 916 OAI21_X2
* cell instance $52363 m0 *1 411.16,46.2
X$52363 1100 1026 1075 44 25 1101 AND3_X1
* cell instance $52364 m0 *1 412.11,46.2
X$52364 1075 1026 1100 25 44 1096 NAND3_X1
* cell instance $52365 m0 *1 412.87,46.2
X$52365 967 1006 1077 44 1076 25 OAI21_X1
* cell instance $52368 m0 *1 416.86,46.2
X$52368 923 920 25 44 1052 NAND2_X1
* cell instance $52371 r0 *1 410.4,46.2
X$52371 1073 1101 1074 25 44 1103 NOR3_X1
* cell instance $52374 r0 *1 411.73,46.2
X$52374 1076 1096 1099 25 44 879 NAND3_X2
* cell instance $52375 r0 *1 413.06,46.2
X$52375 1099 1076 1096 25 1097 44 AOI21_X1
* cell instance $52379 r0 *1 417.43,46.2
X$52379 737 1163 25 44 1027 OR2_X1
* cell instance $52380 m0 *1 418,46.2
X$52380 1078 1027 44 25 989 XNOR2_X1
* cell instance $52382 m0 *1 419.14,46.2
X$52382 1027 1078 44 923 25 XOR2_X2
* cell instance $52383 m0 *1 420.85,46.2
X$52383 1095 1028 44 988 25 XOR2_X2
* cell instance $52384 m0 *1 422.56,46.2
X$52384 1029 1120 25 44 1078 XNOR2_X2
* cell instance $52386 m0 *1 430.54,46.2
X$52386 995 1030 25 44 1029 XNOR2_X2
* cell instance $52388 m0 *1 433.96,46.2
X$52388 1031 1032 1082 44 25 1030 OAI21_X2
* cell instance $52393 r0 *1 421.99,46.2
X$52393 1078 1079 25 44 1094 OR2_X1
* cell instance $52394 r0 *1 422.75,46.2
X$52394 1079 1121 1078 737 25 44 1080 NOR4_X1
* cell instance $52396 r0 *1 423.89,46.2
X$52396 1080 1121 1094 25 992 44 AOI21_X2
* cell instance $52399 r0 *1 431.68,46.2
X$52399 1030 1119 1002 25 44 1135 MUX2_X1
* cell instance $52402 r0 *1 434.72,46.2
X$52402 1125 1083 25 44 996 NAND2_X1
* cell instance $52404 m0 *1 437.38,46.2
X$52404 1081 1033 1082 1089 994 1000 25 44 OAI221_X2
* cell instance $52406 m0 *1 439.47,46.2
X$52406 25 1034 997 1081 1227 1033 44 OAI211_X4
* cell instance $52408 m0 *1 444.22,46.2
X$52408 1035 1083 25 44 1036 NAND2_X1
* cell instance $52411 m0 *1 451.63,46.2
X$52411 998 44 725 25 BUF_X4
* cell instance $52462 r0 *1 438.71,46.2
X$52462 1082 1126 1089 25 1041 44 AOI21_X2
* cell instance $52464 r0 *1 443.08,46.2
X$52464 999 1133 1127 25 1087 44 AOI21_X1
* cell instance $52466 r0 *1 444.6,46.2
X$52466 1086 1084 1174 25 44 1126 MUX2_X1
* cell instance $52467 r0 *1 445.93,46.2
X$52467 998 1087 1086 44 25 1128 OAI21_X2
* cell instance $52470 r0 *1 448.4,46.2
X$52470 1085 25 44 998 INV_X2
* cell instance $52471 r0 *1 448.97,46.2
X$52471 1085 44 1084 25 BUF_X4
* cell instance $52474 r0 *1 452.2,46.2
X$52474 1132 725 1129 44 25 1089 OAI21_X2
* cell instance $52723 m0 *1 336.3,12.6
X$52723 25 235 211 238 183 237 44 FA_X1
* cell instance $52724 m0 *1 339.34,12.6
X$52724 33 158 44 25 237 AND2_X1
* cell instance $52729 m0 *1 351.5,12.6
X$52729 213 60 44 25 278 AND2_X1
* cell instance $52730 m0 *1 352.26,12.6
X$52730 123 41 44 25 281 AND2_X1
* cell instance $52755 r0 *1 337.44,12.6
X$52755 211 25 44 271 INV_X1
* cell instance $52762 r0 *1 341.43,12.6
X$52762 25 238 386 273 92 256 44 FA_X1
* cell instance $52763 r0 *1 344.47,12.6
X$52763 212 25 44 257 INV_X1
* cell instance $52765 r0 *1 350.93,12.6
X$52765 25 214 275 241 281 278 44 FA_X1
* cell instance $52769 r0 *1 357.96,12.6
X$52769 25 215 282 246 283 284 44 FA_X1
* cell instance $52770 m0 *1 359.48,12.6
X$52770 167 39 44 25 215 AND2_X1
* cell instance $52771 m0 *1 358.72,12.6
X$52771 213 26 44 25 284 AND2_X1
* cell instance $52773 m0 *1 361,12.6
X$52773 25 184 245 216 246 126 44 FA_X1
* cell instance $52777 m0 *1 366.51,12.6
X$52777 33 41 44 25 217 AND2_X1
* cell instance $52778 m0 *1 367.27,12.6
X$52778 35 39 44 25 248 AND2_X1
* cell instance $52787 r0 *1 363.28,12.6
X$52787 216 25 44 260 INV_X1
* cell instance $52791 r0 *1 366.32,12.6
X$52791 25 248 327 285 217 261 44 FA_X1
* cell instance $52792 r0 *1 369.36,12.6
X$52792 285 25 44 288 INV_X1
* cell instance $52795 m0 *1 373.73,12.6
X$52795 25 252 219 220 251 128 44 FA_X1
* cell instance $52796 m0 *1 376.96,12.6
X$52796 25 154 252 221 253 129 44 FA_X1
* cell instance $52799 m0 *1 383.23,12.6
X$52799 38 186 44 25 290 AND2_X1
* cell instance $52800 m0 *1 384.75,12.6
X$52800 42 47 44 25 255 AND2_X1
* cell instance $52805 r0 *1 379.24,12.6
X$52805 221 25 44 329 INV_X1
* cell instance $52810 r0 *1 382.47,12.6
X$52810 25 222 263 264 255 290 44 FA_X1
* cell instance $52812 m0 *1 387.41,12.6
X$52812 176 41 25 44 254 NOR2_X1
* cell instance $52815 m0 *1 390.83,12.6
X$52815 188 223 224 25 187 44 AOI21_X1
* cell instance $52816 m0 *1 391.59,12.6
X$52816 249 25 44 224 INV_X1
* cell instance $52817 m0 *1 391.97,12.6
X$52817 229 250 226 44 25 249 HA_X1
* cell instance $52821 r0 *1 391.78,12.6
X$52821 225 315 226 44 223 25 OAI21_X1
* cell instance $52823 m0 *1 395.2,12.6
X$52823 247 158 44 177 25 XOR2_X2
* cell instance $52825 m0 *1 396.91,12.6
X$52825 76 190 25 44 247 NAND2_X1
* cell instance $52828 m0 *1 400.71,12.6
X$52828 76 192 244 193 202 236 44 25 AOI221_X2
* cell instance $52832 m0 *1 405.27,12.6
X$52832 194 227 25 44 242 NOR2_X1
* cell instance $52842 r0 *1 399.95,12.6
X$52842 266 267 268 25 44 176 NAND3_X2
* cell instance $52843 r0 *1 401.28,12.6
X$52843 28 25 44 268 INV_X1
* cell instance $52844 r0 *1 401.66,12.6
X$52844 192 266 242 44 25 244 AND3_X1
* cell instance $52846 r0 *1 404.13,12.6
X$52846 267 28 2898 44 25 227 HA_X1
* cell instance $52850 r0 *1 408.12,12.6
X$52850 25 30 287 43 239 160 44 DFFR_X2
* cell instance $52851 m0 *1 410.21,12.6
X$52851 240 82 25 44 287 NOR2_X1
* cell instance $52854 m0 *1 410.97,12.6
X$52854 239 200 25 44 240 XOR2_X1
* cell instance $52857 m0 *1 413.82,12.6
X$52857 196 229 168 25 44 136 NAND3_X1
* cell instance $52861 r0 *1 412.3,12.6
X$52861 236 228 25 44 286 NOR2_X1
* cell instance $52864 r0 *1 415.15,12.6
X$52864 25 30 230 43 269 168 44 DFFR_X2
* cell instance $52865 r0 *1 419.33,12.6
X$52865 80 25 44 272 INV_X1
* cell instance $52866 r0 *1 419.71,12.6
X$52866 25 30 233 43 231 229 44 DFFR_X2
* cell instance $52868 m0 *1 422.56,12.6
X$52868 231 234 44 25 232 XNOR2_X1
* cell instance $52881 r0 *1 424.08,12.6
X$52881 232 195 25 44 233 NOR2_X1
* cell instance $53142 m0 *1 333.26,18.2
X$53142 25 293 380 383 317 340 44 FA_X1
* cell instance $53161 r0 *1 331.74,18.2
X$53161 36 158 44 25 360 AND2_X1
* cell instance $53164 r0 *1 336.3,18.2
X$53164 25 271 382 384 361 383 44 FA_X1
* cell instance $53166 m0 *1 336.68,18.2
X$53166 38 60 44 25 340 AND2_X1
* cell instance $53170 r0 *1 339.72,18.2
X$53170 25 386 425 387 342 384 44 FA_X1
* cell instance $53172 m0 *1 344.09,18.2
X$53172 25 295 342 256 345 344 44 FA_X1
* cell instance $53174 m0 *1 347.13,18.2
X$53174 213 189 44 25 344 AND2_X1
* cell instance $53175 m0 *1 347.89,18.2
X$53175 123 32 44 25 345 AND2_X1
* cell instance $53178 r0 *1 344.28,18.2
X$53178 32 323 25 44 385 NAND2_X1
* cell instance $53180 r0 *1 350.93,18.2
X$53180 25 310 362 363 389 388 44 FA_X1
* cell instance $53181 m0 *1 352.26,18.2
X$53181 41 323 25 44 389 NAND2_X1
* cell instance $53185 m0 *1 355.11,18.2
X$53185 39 323 25 44 390 NAND2_X1
* cell instance $53186 m0 *1 355.68,18.2
X$53186 258 25 44 324 INV_X1
* cell instance $53188 m0 *1 362.14,18.2
X$53188 167 40 44 25 311 AND2_X1
* cell instance $53189 m0 *1 362.9,18.2
X$53189 123 48 44 25 314 AND2_X1
* cell instance $53190 m0 *1 363.66,18.2
X$53190 25 327 325 366 350 326 44 FA_X1
* cell instance $53193 m0 *1 368.98,18.2
X$53193 167 48 44 25 395 AND2_X1
* cell instance $53195 m0 *1 371.26,18.2
X$53195 42 189 44 25 317 AND2_X1
* cell instance $53199 r0 *1 353.97,18.2
X$53199 25 324 364 452 390 259 44 FA_X1
* cell instance $53205 r0 *1 361.57,18.2
X$53205 25 325 392 472 296 260 44 FA_X1
* cell instance $53208 r0 *1 366.89,18.2
X$53208 366 25 44 394 INV_X1
* cell instance $53211 r0 *1 367.84,18.2
X$53211 25 395 393 351 367 368 44 FA_X1
* cell instance $53214 m0 *1 377.15,18.2
X$53214 25 299 358 330 328 329 44 FA_X1
* cell instance $53216 m0 *1 380.19,18.2
X$53216 27 40 44 25 320 AND2_X1
* cell instance $53220 r0 *1 377.15,18.2
X$53220 467 25 44 167 BUF_X2
* cell instance $53221 r0 *1 377.91,18.2
X$53221 123 291 44 25 359 AND2_X1
* cell instance $53224 r0 *1 379.81,18.2
X$53224 330 25 44 369 INV_X1
* cell instance $53226 m0 *1 385.32,18.2
X$53226 301 36 25 44 357 NAND2_X1
* cell instance $53230 m0 *1 386.27,18.2
X$53230 25 355 354 353 356 357 44 FA_X1
* cell instance $53233 m0 *1 391.4,18.2
X$53233 33 301 44 25 352 AND2_X1
* cell instance $53237 m0 *1 393.11,18.2
X$53237 300 346 331 25 315 44 AOI21_X1
* cell instance $53238 m0 *1 393.87,18.2
X$53238 349 25 44 331 INV_X1
* cell instance $53242 m0 *1 396.72,18.2
X$53242 334 348 347 44 25 349 HA_X1
* cell instance $53245 m0 *1 401.66,18.2
X$53245 267 268 400 44 25 343 HA_X1
* cell instance $53251 r0 *1 396.91,18.2
X$53251 412 370 347 44 346 25 OAI21_X1
* cell instance $53256 r0 *1 400.52,18.2
X$53256 343 25 44 308 INV_X1
* cell instance $53258 r0 *1 402.42,18.2
X$53258 186 343 44 25 371 XNOR2_X1
* cell instance $53261 m0 *1 407.36,18.2
X$53261 341 25 44 333 INV_X1
* cell instance $53262 m0 *1 405.46,18.2
X$53262 339 267 332 44 25 341 HA_X1
* cell instance $53267 r0 *1 406.41,18.2
X$53267 398 25 44 372 INV_X1
* cell instance $53268 r0 *1 406.79,18.2
X$53268 332 333 402 44 399 25 OAI21_X1
* cell instance $53269 r0 *1 407.55,18.2
X$53269 376 400 402 44 25 398 HA_X1
* cell instance $53270 m0 *1 409.07,18.2
X$53270 25 30 338 43 339 335 44 DFFR_X2
* cell instance $53272 m0 *1 413.25,18.2
X$53272 82 335 25 44 338 NOR2_X1
* cell instance $53275 r0 *1 412.49,18.2
X$53275 25 30 337 43 375 376 44 DFFR_X2
* cell instance $53277 m0 *1 414.2,18.2
X$53277 82 374 25 44 337 NOR2_X1
* cell instance $53279 m0 *1 422.37,18.2
X$53279 25 30 304 43 2892 334 44 DFFR_X2
* cell instance $53295 r0 *1 419.33,18.2
X$53295 302 336 270 25 44 80 NAND3_X2
* cell instance $53298 r0 *1 422.37,18.2
X$53298 336 378 25 44 379 XOR2_X1
* cell instance $53299 r0 *1 423.51,18.2
X$53299 379 195 25 44 377 NOR2_X1
* cell instance $53582 m0 *1 346.37,9.8
X$53582 32 167 25 44 198 NAND2_X1
* cell instance $53604 r0 *1 337.25,9.8
X$53604 36 34 44 25 235 AND2_X1
* cell instance $53609 r0 *1 345.04,9.8
X$53609 25 198 212 122 199 155 44 FA_X1
* cell instance $53610 r0 *1 348.08,9.8
X$53610 158 213 25 44 155 NAND2_X1
* cell instance $53611 m0 *1 348.27,9.8
X$53611 142 25 44 169 INV_X1
* cell instance $53617 m0 *1 353.02,9.8
X$53617 25 172 243 259 145 171 44 FA_X1
* cell instance $53620 m0 *1 356.82,9.8
X$53620 167 41 44 25 124 AND2_X1
* cell instance $53621 m0 *1 357.58,9.8
X$53621 213 34 44 25 147 AND2_X1
* cell instance $53633 m0 *1 364.04,9.8
X$53633 25 127 184 185 178 175 44 FA_X1
* cell instance $53638 r0 *1 365.37,9.8
X$53638 185 25 44 326 INV_X1
* cell instance $53640 m0 *1 369.93,9.8
X$53640 213 41 44 25 179 AND2_X1
* cell instance $53642 m0 *1 370.69,9.8
X$53642 25 207 218 152 180 179 44 FA_X1
* cell instance $53646 r0 *1 371.83,9.8
X$53646 167 47 44 25 207 AND2_X1
* cell instance $53648 r0 *1 375.63,9.8
X$53648 25 182 251 253 208 181 44 FA_X1
* cell instance $53650 m0 *1 376.39,9.8
X$53650 123 186 44 25 208 AND2_X1
* cell instance $53652 m0 *1 378.48,9.8
X$53652 27 39 44 25 181 AND2_X1
* cell instance $53658 m0 *1 390.64,9.8
X$53658 187 156 157 44 131 25 OAI21_X1
* cell instance $53662 m0 *1 396.72,9.8
X$53662 160 177 78 44 25 191 HA_X1
* cell instance $53671 r0 *1 389.12,9.8
X$53671 168 149 210 44 25 156 HA_X1
* cell instance $53672 r0 *1 391.02,9.8
X$53672 210 25 44 188 INV_X1
* cell instance $53675 r0 *1 393.3,9.8
X$53675 189 209 44 25 204 XNOR2_X1
* cell instance $53676 r0 *1 394.44,9.8
X$53676 176 107 158 60 25 44 209 NOR4_X1
* cell instance $53678 r0 *1 395.39,9.8
X$53678 189 158 31 107 44 192 25 NOR4_X2
* cell instance $53680 r0 *1 397.29,9.8
X$53680 107 60 25 44 190 NOR2_X1
* cell instance $53682 r0 *1 398.24,9.8
X$53682 206 191 205 44 202 25 OAI21_X1
* cell instance $53684 r0 *1 399.38,9.8
X$53684 159 204 205 44 25 203 HA_X1
* cell instance $53686 r0 *1 401.66,9.8
X$53686 203 25 44 193 INV_X1
* cell instance $53690 r0 *1 404.13,9.8
X$53690 201 28 2899 44 25 194 HA_X1
* cell instance $53692 m0 *1 407.55,9.8
X$53692 25 30 174 43 173 159 44 DFFR_X2
* cell instance $53694 m0 *1 411.73,9.8
X$53694 160 25 44 170 INV_X1
* cell instance $53695 m0 *1 412.11,9.8
X$53695 166 54 57 25 44 161 NAND3_X1
* cell instance $53696 m0 *1 412.87,9.8
X$53696 161 81 170 25 44 137 NOR3_X1
* cell instance $53699 r0 *1 412.49,9.8
X$53699 161 80 25 44 200 NOR2_X1
* cell instance $53701 m0 *1 414.2,9.8
X$53701 136 81 25 44 165 NOR2_X1
* cell instance $53703 m0 *1 414.77,9.8
X$53703 132 165 44 25 162 XNOR2_X1
* cell instance $53704 m0 *1 415.91,9.8
X$53704 162 195 25 44 134 NOR2_X1
* cell instance $53705 m0 *1 416.48,9.8
X$53705 25 30 134 43 2893 132 44 DFFR_X2
* cell instance $53706 m0 *1 420.66,9.8
X$53706 163 80 44 25 164 XNOR2_X1
* cell instance $53762 r0 *1 414.96,9.8
X$53762 82 25 44 195 CLKBUF_X3
* cell instance $53765 r0 *1 417.62,9.8
X$53765 25 30 197 43 163 196 44 DFFR_X2
* cell instance $53766 r0 *1 421.8,9.8
X$53766 164 195 25 44 197 NOR2_X1
* cell instance $54013 m0 *1 340.1,7
X$54013 25 67 92 138 91 66 44 FA_X1
* cell instance $54014 m0 *1 343.14,7
X$54014 38 25 44 36 BUF_X2
* cell instance $54017 m0 *1 347.13,7
X$54017 35 34 44 25 67 AND2_X1
* cell instance $54046 r0 *1 342.95,7
X$54046 138 25 44 141 INV_X1
* cell instance $54048 r0 *1 344.09,7
X$54048 25 68 274 142 140 141 44 FA_X1
* cell instance $54049 r0 *1 347.13,7
X$54049 122 25 44 140 INV_X1
* cell instance $54053 m0 *1 349.03,7
X$54053 97 25 44 143 INV_X1
* cell instance $54058 r0 *1 349.6,7
X$54058 25 69 277 144 241 143 44 FA_X1
* cell instance $54059 r0 *1 352.64,7
X$54059 144 25 44 171 INV_X1
* cell instance $54062 m0 *1 355.3,7
X$54062 25 62 172 104 102 101 44 FA_X1
* cell instance $54064 m0 *1 358.34,7
X$54064 104 25 44 125 INV_X1
* cell instance $54068 m0 *1 369.36,7
X$54068 35 40 44 25 110 AND2_X1
* cell instance $54071 m0 *1 371.83,7
X$54071 25 71 70 72 152 115 44 FA_X1
* cell instance $54075 r0 *1 355.49,7
X$54075 123 39 44 25 146 AND2_X1
* cell instance $54076 r0 *1 356.25,7
X$54076 25 124 145 102 146 147 44 FA_X1
* cell instance $54084 r0 *1 364.04,7
X$54084 36 39 44 25 175 AND2_X1
* cell instance $54085 r0 *1 365.56,7
X$54085 35 41 44 25 127 AND2_X1
* cell instance $54090 r0 *1 374.87,7
X$54090 72 25 44 128 INV_X1
* cell instance $54093 m0 *1 378.29,7
X$54093 73 25 44 129 INV_X1
* cell instance $54098 m0 *1 381.33,7
X$54098 25 74 154 153 120 121 44 FA_X1
* cell instance $54101 r0 *1 382.28,7
X$54101 153 25 44 130 INV_X1
* cell instance $54106 m0 *1 389.12,7
X$54106 76 50 25 44 150 NAND2_X1
* cell instance $54109 m0 *1 391.97,7
X$54109 77 131 109 25 103 44 AOI21_X1
* cell instance $54110 m0 *1 392.73,7
X$54110 133 25 44 109 INV_X1
* cell instance $54115 r0 *1 385.89,7
X$54115 151 26 44 148 25 XOR2_X2
* cell instance $54119 r0 *1 388.93,7
X$54119 150 32 44 149 25 XOR2_X2
* cell instance $54120 r0 *1 390.64,7
X$54120 132 148 157 44 25 133 HA_X1
* cell instance $54126 m0 *1 395.77,7
X$54126 176 107 25 44 105 NOR2_X1
* cell instance $54128 m0 *1 397.86,7
X$54128 93 94 79 25 206 44 AOI21_X1
* cell instance $54129 m0 *1 397.48,7
X$54129 78 25 44 93 INV_X1
* cell instance $54133 m0 *1 399,7
X$54133 90 25 44 47 CLKBUF_X3
* cell instance $54136 m0 *1 412.87,7
X$54136 87 80 25 44 86 NOR2_X1
* cell instance $54137 m0 *1 413.44,7
X$54137 87 81 83 25 44 84 NOR3_X1
* cell instance $54195 r0 *1 410.02,7
X$54195 139 82 25 44 174 NOR2_X1
* cell instance $54196 r0 *1 410.59,7
X$54196 173 137 25 44 139 XOR2_X1
* cell instance $54198 r0 *1 413.25,7
X$54198 132 25 44 135 INV_X1
* cell instance $54199 r0 *1 413.63,7
X$54199 136 135 25 44 166 NOR2_X1
* cell instance $54200 r0 *1 414.2,7
X$54200 135 136 25 44 87 OR2_X1
* cell instance $54436 r0 *1 340.1,4.2
X$54436 33 60 44 25 91 AND2_X1
* cell instance $54437 r0 *1 340.86,4.2
X$54437 36 26 44 25 66 AND2_X1
* cell instance $54441 m0 *1 345.99,4.2
X$54441 36 32 44 25 95 AND2_X1
* cell instance $54443 r0 *1 346.18,4.2
X$54443 25 45 68 97 96 95 44 FA_X1
* cell instance $54444 m0 *1 347.32,4.2
X$54444 33 34 44 25 96 AND2_X1
* cell instance $54446 m0 *1 348.08,4.2
X$54446 35 26 44 25 45 AND2_X1
* cell instance $54453 m0 *1 352.45,4.2
X$54453 35 32 44 25 61 AND2_X1
* cell instance $54454 m0 *1 353.21,4.2
X$54454 33 26 44 25 100 AND2_X1
* cell instance $54459 r0 *1 351.69,4.2
X$54459 25 61 69 98 100 99 44 FA_X1
* cell instance $54460 r0 *1 354.73,4.2
X$54460 98 25 44 101 INV_X1
* cell instance $54468 m0 *1 361.19,4.2
X$54468 33 32 44 25 63 AND2_X1
* cell instance $54469 m0 *1 361.95,4.2
X$54469 25 64 62 106 63 37 44 FA_X1
* cell instance $54473 r0 *1 363.09,4.2
X$54473 106 25 44 126 INV_X1
* cell instance $54474 r0 *1 363.47,4.2
X$54474 36 41 44 25 37 AND2_X1
* cell instance $54478 r0 *1 368.41,4.2
X$54478 25 110 113 111 112 46 44 FA_X1
* cell instance $54479 m0 *1 369.93,4.2
X$54479 33 39 44 25 112 AND2_X1
* cell instance $54480 m0 *1 369.17,4.2
X$54480 38 48 44 25 46 AND2_X1
* cell instance $54484 r0 *1 371.45,4.2
X$54484 111 25 44 115 INV_X1
* cell instance $54488 r0 *1 374.49,4.2
X$54488 38 47 44 25 118 AND2_X1
* cell instance $54489 r0 *1 375.25,4.2
X$54489 25 65 71 73 119 118 44 FA_X1
* cell instance $54491 m0 *1 375.63,4.2
X$54491 42 40 44 25 119 AND2_X1
* cell instance $54492 m0 *1 376.96,4.2
X$54492 35 48 44 25 65 AND2_X1
* cell instance $54499 r0 *1 382.09,4.2
X$54499 42 48 44 25 120 AND2_X1
* cell instance $54500 r0 *1 382.85,4.2
X$54500 35 47 44 25 74 AND2_X1
* cell instance $54503 m0 *1 387.41,4.2
X$54503 49 25 44 41 CLKBUF_X3
* cell instance $54504 m0 *1 388.93,4.2
X$54504 42 25 44 33 BUF_X2
* cell instance $54507 m0 *1 396.53,4.2
X$54507 57 59 52 44 25 53 HA_X1
* cell instance $54510 r0 *1 383.61,4.2
X$54510 34 25 44 51 INV_X1
* cell instance $54513 r0 *1 387.41,4.2
X$54513 32 26 25 44 75 NOR2_X1
* cell instance $54514 r0 *1 387.98,4.2
X$54514 75 50 51 25 44 107 NAND3_X2
* cell instance $54515 r0 *1 389.31,4.2
X$54515 76 75 50 25 44 117 NAND3_X1
* cell instance $54517 r0 *1 390.26,4.2
X$54517 51 117 44 25 116 XNOR2_X1
* cell instance $54519 r0 *1 391.78,4.2
X$54519 114 25 44 77 INV_X1
* cell instance $54520 r0 *1 392.16,4.2
X$54520 54 116 114 44 25 108 HA_X1
* cell instance $54522 r0 *1 394.82,4.2
X$54522 108 103 52 44 94 25 OAI21_X1
* cell instance $54523 r0 *1 395.58,4.2
X$54523 60 105 44 25 59 XNOR2_X1
* cell instance $54524 r0 *1 396.72,4.2
X$54524 31 25 44 60 CLKBUF_X3
* cell instance $54526 r0 *1 398.43,4.2
X$54526 53 25 44 79 INV_X1
* cell instance $54534 m0 *1 407.55,4.2
X$54534 25 30 58 43 89 57 44 DFFR_X2
* cell instance $54536 m0 *1 412.49,4.2
X$54536 55 86 25 44 85 XOR2_X1
* cell instance $54537 m0 *1 413.63,4.2
X$54537 25 30 56 43 55 54 44 DFFR_X2
* cell instance $54596 r0 *1 409.64,4.2
X$54596 88 82 25 44 58 NOR2_X1
* cell instance $54598 r0 *1 410.59,4.2
X$54598 89 84 25 44 88 XOR2_X1
* cell instance $54601 r0 *1 413.63,4.2
X$54601 54 25 44 83 INV_X1
* cell instance $54602 r0 *1 414.01,4.2
X$54602 85 82 25 44 56 NOR2_X1
* cell instance $54844 m0 *1 334.21,49
X$54844 833 893 44 1140 25 XOR2_X2
* cell instance $54845 m0 *1 335.92,49
X$54845 1040 1088 1140 44 1138 25 OAI21_X1
* cell instance $54864 r0 *1 334.02,49
X$54864 893 833 25 44 1141 XNOR2_X2
* cell instance $54865 r0 *1 335.92,49
X$54865 1195 1057 1141 25 44 1183 NAND3_X1
* cell instance $54869 r0 *1 340.67,49
X$54869 1197 1198 1237 44 1236 25 OAI21_X1
* cell instance $54870 r0 *1 341.43,49
X$54870 834 1144 44 25 1198 XNOR2_X1
* cell instance $54872 r0 *1 343.33,49
X$54872 1200 1110 835 25 44 1238 NAND3_X2
* cell instance $54873 m0 *1 344.66,49
X$54873 835 1046 25 44 1108 NOR2_X1
* cell instance $54874 m0 *1 343.9,49
X$54874 1061 1107 1108 44 1237 25 OAI21_X1
* cell instance $54875 m0 *1 345.23,49
X$54875 1110 1184 1061 1045 44 1142 25 NOR4_X2
* cell instance $54879 m0 *1 349.41,49
X$54879 1184 44 1107 25 BUF_X4
* cell instance $54882 m0 *1 352.45,49
X$54882 1060 1111 1146 25 44 NOR2_X4
* cell instance $54883 m0 *1 354.16,49
X$54883 1148 1149 957 1112 25 1184 44 NAND4_X2
* cell instance $54885 m0 *1 356.06,49
X$54885 25 958 959 1150 1145 1110 44 NOR4_X4
* cell instance $54890 r0 *1 344.66,49
X$54890 835 1200 1144 25 1143 44 AOI21_X2
* cell instance $54891 r0 *1 345.99,49
X$54891 25 1111 1060 1042 1200 44 NOR3_X4
* cell instance $54894 r0 *1 349.79,49
X$54894 1241 1183 1107 25 44 1296 OR3_X1
* cell instance $54895 r0 *1 350.74,49
X$54895 1141 1134 1204 1145 44 1203 25 OR4_X2
* cell instance $54896 r0 *1 352.07,49
X$54896 1145 1204 1138 1183 1245 1244 25 44 1147 OAI33_X1
* cell instance $54898 r0 *1 353.59,49
X$54898 1112 1148 25 44 1245 NAND2_X1
* cell instance $54900 r0 *1 354.35,49
X$54900 1148 1149 957 25 44 1204 NAND3_X1
* cell instance $54903 r0 *1 356.06,49
X$54903 25 958 959 1150 1145 1144 44 NOR4_X4
* cell instance $54910 m0 *1 365.18,49
X$54910 25 1019 978 870 1148 44 NOR3_X4
* cell instance $54913 r0 *1 365.56,49
X$54913 1151 1019 25 44 1205 NOR2_X1
* cell instance $54916 r0 *1 367.27,49
X$54916 1019 1151 25 44 1246 OR2_X1
* cell instance $54919 r0 *1 368.6,49
X$54919 1151 1019 1111 25 44 1247 NAND3_X1
* cell instance $54921 m0 *1 368.98,49
X$54921 1193 1111 1112 25 44 1249 MUX2_X1
* cell instance $54922 m0 *1 370.5,49
X$54922 25 1020 1113 1063 904 1151 44 NAND4_X4
* cell instance $54925 r0 *1 369.36,49
X$54925 1247 1246 1249 44 25 1207 OAI21_X2
* cell instance $54926 r0 *1 370.69,49
X$54926 1208 1209 25 44 1193 NAND2_X1
* cell instance $54929 r0 *1 371.83,49
X$54929 870 1208 44 25 1210 XNOR2_X1
* cell instance $54930 r0 *1 372.97,49
X$54930 1113 1020 1063 25 44 1251 NAND3_X1
* cell instance $54932 m0 *1 376.01,49
X$54932 1113 1020 25 1145 44 NAND2_X4
* cell instance $54934 m0 *1 377.72,49
X$54934 25 1152 1153 1064 1154 1113 44 NOR4_X4
* cell instance $54939 r0 *1 377.15,49
X$54939 1152 1153 1064 1154 44 1253 25 OR4_X2
* cell instance $54940 r0 *1 378.48,49
X$54940 979 1155 1021 1156 44 25 1208 AND4_X2
* cell instance $54941 r0 *1 379.81,49
X$54941 25 1021 1156 979 1155 1271 44 NAND4_X4
* cell instance $54944 m0 *1 385.51,49
X$54944 908 909 1157 1114 1115 1154 25 44 OAI221_X2
* cell instance $54949 m0 *1 392.35,49
X$54949 1115 1215 25 44 1119 XNOR2_X2
* cell instance $54953 m0 *1 402.04,49
X$54953 1100 981 915 44 25 1116 AND3_X1
* cell instance $54957 m0 *1 406.98,49
X$54957 1105 967 25 44 1161 NOR2_X1
* cell instance $54961 r0 *1 385.51,49
X$54961 1156 1155 25 44 1212 NAND2_X2
* cell instance $54962 r0 *1 386.46,49
X$54962 1114 1157 1115 44 1255 25 OAI21_X1
* cell instance $54964 r0 *1 387.41,49
X$54964 1212 1158 44 1190 25 XOR2_X2
* cell instance $54966 r0 *1 390.64,49
X$54966 1115 1215 44 25 1156 AND2_X2
* cell instance $54969 r0 *1 392.54,49
X$54969 1215 1115 44 1222 25 XOR2_X2
* cell instance $54970 r0 *1 394.25,49
X$54970 1257 1159 25 44 1260 XNOR2_X2
* cell instance $54971 r0 *1 396.15,49
X$54971 1066 25 44 1274 CLKBUF_X3
* cell instance $54975 r0 *1 402.42,49
X$54975 947 1260 25 44 1220 NAND2_X2
* cell instance $54978 r0 *1 404.32,49
X$54978 1100 751 1160 25 44 1023 OR3_X1
* cell instance $54979 r0 *1 405.27,49
X$54979 751 1160 1025 44 1261 25 OAI21_X1
* cell instance $54980 r0 *1 406.03,49
X$54980 982 1218 987 44 1160 25 OAI21_X1
* cell instance $54981 r0 *1 406.79,49
X$54981 1262 1161 1219 967 1261 1118 44 25 AOI221_X2
* cell instance $54982 r0 *1 408.88,49
X$54982 1119 1100 947 25 1168 44 NAND3_X4
* cell instance $54984 m0 *1 413.06,49
X$54984 1077 25 44 1194 INV_X1
* cell instance $54985 m0 *1 411.73,49
X$54985 1194 1100 1026 25 1073 44 AOI21_X2
* cell instance $54986 m0 *1 413.44,49
X$54986 1074 25 44 1099 INV_X1
* cell instance $54991 r0 *1 413.25,49
X$54991 737 1162 25 44 1077 NOR2_X1
* cell instance $54992 r0 *1 413.82,49
X$54992 1099 1258 25 44 1300 NOR2_X1
* cell instance $54997 r0 *1 417.24,49
X$54997 1162 1221 25 44 1163 NOR2_X1
* cell instance $54998 r0 *1 417.81,49
X$54998 1221 1258 1162 25 1079 44 AOI21_X1
* cell instance $55001 m0 *1 421.99,49
X$55001 1028 1119 25 44 1282 NAND2_X2
* cell instance $55003 m0 *1 422.94,49
X$55003 1282 633 25 44 1120 NOR2_X1
* cell instance $55004 m0 *1 423.51,49
X$55004 1123 1192 25 44 1121 XNOR2_X2
* cell instance $55009 r0 *1 422.56,49
X$55009 1164 1028 44 25 1223 XNOR2_X1
* cell instance $55011 r0 *1 424.08,49
X$55011 1165 633 25 44 1192 NOR2_X1
* cell instance $55014 m0 *1 428.26,49
X$55014 1029 1122 25 44 1166 NOR2_X1
* cell instance $55016 m0 *1 428.83,49
X$55016 1122 1123 25 44 1167 NAND2_X1
* cell instance $55019 m0 *1 431.11,49
X$55019 1001 1135 44 25 1252 XNOR2_X1
* cell instance $55021 r0 *1 428.45,49
X$55021 1123 1166 1224 1165 1167 1252 25 44 1191 OAI33_X1
* cell instance $55023 r0 *1 430.16,49
X$55023 1254 1081 25 44 1133 NOR2_X1
* cell instance $55025 m0 *1 432.82,49
X$55025 1190 725 25 44 1001 XNOR2_X2
* cell instance $55030 r0 *1 435.29,49
X$55030 1225 1171 25 44 1127 NOR2_X1
* cell instance $55031 m0 *1 436.05,49
X$55031 1127 1084 1124 25 44 1125 MUX2_X1
* cell instance $55033 m0 *1 437.38,49
X$55033 1189 1170 1084 44 25 1033 MUX2_X2
* cell instance $55035 m0 *1 439.85,49
X$55035 1031 1133 1125 25 1188 44 AOI21_X1
* cell instance $55037 r0 *1 435.86,49
X$55037 1171 1225 25 44 1189 OR2_X1
* cell instance $55039 r0 *1 436.81,49
X$55039 1226 1169 25 44 1124 NOR2_X1
* cell instance $55041 r0 *1 437.76,49
X$55041 1169 1226 25 44 1170 OR2_X1
* cell instance $55044 r0 *1 439.09,49
X$55044 25 1168 1031 1228 1187 1343 44 NOR4_X4
* cell instance $55045 m0 *1 441.18,49
X$55045 1188 1126 1089 44 1172 25 OAI21_X1
* cell instance $55048 m0 *1 442.7,49
X$55048 1185 998 1186 25 1187 44 AOI21_X2
* cell instance $55049 m0 *1 444.03,49
X$55049 1174 1170 998 25 44 1185 NOR3_X1
* cell instance $55051 m0 *1 445.55,49
X$55051 998 1174 25 44 1243 OR2_X1
* cell instance $55055 m0 *1 451.63,49
X$55055 998 1177 25 44 1175 OR2_X1
* cell instance $55057 m0 *1 452.58,49
X$55057 998 1177 1178 44 1132 25 OAI21_X1
* cell instance $55058 m0 *1 453.34,49
X$55058 1179 1176 44 25 1177 AND2_X1
* cell instance $55061 m0 *1 455.05,49
X$55061 1176 1130 44 25 1235 XNOR2_X1
* cell instance $55063 m0 *1 456.95,49
X$55063 1180 1181 1131 25 1129 44 AOI21_X1
* cell instance $55071 r0 *1 442.7,49
X$55071 1190 1173 1127 44 25 1186 AND3_X1
* cell instance $55072 r0 *1 443.65,49
X$55072 1133 25 44 1239 INV_X1
* cell instance $55075 r0 *1 444.6,49
X$55075 1170 1174 25 44 1240 OR2_X1
* cell instance $55077 r0 *1 445.55,49
X$55077 1084 1086 1243 44 1229 25 OAI21_X1
* cell instance $55078 r0 *1 446.31,49
X$55078 1173 1190 25 44 1086 NAND2_X1
* cell instance $55079 r0 *1 446.88,49
X$55079 1239 1240 1174 1340 1084 1290 25 44 OAI221_X2
* cell instance $55081 r0 *1 449.35,49
X$55081 25 1084 1234 1228 1178 1175 44 AOI22_X4
* cell instance $55082 r0 *1 452.58,49
X$55082 1176 25 44 1230 INV_X1
* cell instance $55083 r0 *1 452.96,49
X$55083 1130 1182 25 44 1178 NOR2_X2
* cell instance $55084 r0 *1 453.91,49
X$55084 1231 25 44 1182 INV_X1
* cell instance $55085 r0 *1 454.29,49
X$55085 1231 1179 25 44 1233 OR2_X1
* cell instance $55086 r0 *1 455.05,49
X$55086 1232 1233 1235 44 25 1234 OAI21_X2
* cell instance $55087 r0 *1 456.38,49
X$55087 1231 1179 1230 1130 44 25 1180 AND4_X1
* cell instance $55089 r0 *1 457.9,49
X$55089 1179 1231 25 44 1181 NOR2_X1
* cell instance $55366 m0 *1 327.18,40.6
X$55366 890 768 931 44 25 933 HA_X1
* cell instance $55386 r0 *1 326.61,40.6
X$55386 513 189 44 25 932 AND2_X1
* cell instance $55388 r0 *1 327.56,40.6
X$55388 932 831 890 44 25 951 HA_X1
* cell instance $55390 r0 *1 329.65,40.6
X$55390 931 25 44 893 BUF_X2
* cell instance $55392 r0 *1 330.6,40.6
X$55392 933 25 44 1004 INV_X1
* cell instance $55394 r0 *1 331.17,40.6
X$55394 951 891 25 44 892 OR2_X1
* cell instance $55396 r0 *1 332.12,40.6
X$55396 798 797 893 44 891 25 OAI21_X1
* cell instance $55398 r0 *1 333.07,40.6
X$55398 894 798 893 44 970 25 OAI21_X1
* cell instance $55401 r0 *1 336.11,40.6
X$55401 892 643 25 44 1013 NOR2_X2
* cell instance $55402 m0 *1 337.25,40.6
X$55402 797 25 44 895 INV_X1
* cell instance $55404 m0 *1 337.63,40.6
X$55404 25 797 865 934 896 44 NOR3_X4
* cell instance $55406 m0 *1 341.05,40.6
X$55406 897 889 899 25 898 44 AOI21_X2
* cell instance $55407 m0 *1 342.38,40.6
X$55407 739 836 889 899 865 44 25 AOI211_X2
* cell instance $55409 m0 *1 345.61,40.6
X$55409 739 836 25 44 901 NOR2_X1
* cell instance $55412 m0 *1 347.13,40.6
X$55412 25 936 856 889 899 44 AOI21_X4
* cell instance $55413 m0 *1 349.6,40.6
X$55413 803 807 44 25 867 AND2_X1
* cell instance $55414 m0 *1 350.36,40.6
X$55414 867 804 866 803 956 44 25 AOI211_X2
* cell instance $55419 r0 *1 337.25,40.6
X$55419 864 895 25 44 894 NOR2_X2
* cell instance $55420 r0 *1 338.2,40.6
X$55420 934 865 797 44 1015 25 OAI21_X1
* cell instance $55421 r0 *1 338.96,40.6
X$55421 864 643 44 25 952 AND2_X2
* cell instance $55424 r0 *1 340.86,40.6
X$55424 836 739 892 25 44 897 OR3_X1
* cell instance $55427 r0 *1 345.04,40.6
X$55427 835 900 954 936 25 44 972 NOR4_X1
* cell instance $55428 r0 *1 345.99,40.6
X$55428 901 807 866 44 25 953 OAI21_X4
* cell instance $55432 r0 *1 352.64,40.6
X$55432 527 956 25 44 957 XNOR2_X2
* cell instance $55434 r0 *1 354.73,40.6
X$55434 956 527 44 958 25 XOR2_X2
* cell instance $55435 r0 *1 356.44,40.6
X$55435 707 528 44 959 25 XOR2_X2
* cell instance $55437 r0 *1 358.34,40.6
X$55437 25 903 937 750 1111 44 NOR3_X4
* cell instance $55438 m0 *1 359.48,40.6
X$55438 654 868 902 25 937 44 AOI21_X2
* cell instance $55440 m0 *1 360.81,40.6
X$55440 868 902 624 44 25 903 AND3_X1
* cell instance $55441 m0 *1 361.76,40.6
X$55441 25 868 902 866 870 869 44 OAI211_X4
* cell instance $55442 m0 *1 364.99,40.6
X$55442 581 807 44 25 871 AND2_X1
* cell instance $55444 m0 *1 365.94,40.6
X$55444 772 942 871 899 888 904 44 25 AOI221_X2
* cell instance $55448 m0 *1 372.78,40.6
X$55448 658 778 25 44 905 OR2_X1
* cell instance $55450 m0 *1 373.73,40.6
X$55450 872 658 25 44 873 NOR2_X1
* cell instance $55452 m0 *1 375.06,40.6
X$55452 774 25 44 1009 INV_X1
* cell instance $55456 r0 *1 361.19,40.6
X$55456 903 937 750 25 44 960 OR3_X1
* cell instance $55458 r0 *1 363.66,40.6
X$55458 772 941 938 25 44 902 NAND3_X2
* cell instance $55460 r0 *1 365.37,40.6
X$55460 792 938 941 25 899 44 NAND3_X4
* cell instance $55463 r0 *1 368.79,40.6
X$55463 773 792 44 25 1007 AND2_X1
* cell instance $55466 r0 *1 372.97,40.6
X$55466 905 938 941 25 974 44 AOI21_X1
* cell instance $55467 r0 *1 373.73,40.6
X$55467 974 774 872 658 907 1211 25 44 OAI221_X2
* cell instance $55468 r0 *1 375.82,40.6
X$55468 908 909 906 44 907 25 OAI21_X1
* cell instance $55469 r0 *1 376.58,40.6
X$55469 908 909 910 44 963 25 OAI21_X1
* cell instance $55471 m0 *1 376.58,40.6
X$55471 778 658 25 44 910 NOR2_X1
* cell instance $55476 r0 *1 378.48,40.6
X$55476 911 779 25 44 909 NAND2_X2
* cell instance $55477 r0 *1 379.43,40.6
X$55477 964 973 908 44 25 1021 OAI21_X2
* cell instance $55479 m0 *1 380,40.6
X$55479 810 787 25 44 911 OR2_X2
* cell instance $55484 r0 *1 381.14,40.6
X$55484 25 1098 789 912 946 44 AOI21_X4
* cell instance $55485 r0 *1 383.61,40.6
X$55485 787 863 25 44 1011 NOR2_X1
* cell instance $55486 r0 *1 384.18,40.6
X$55486 863 25 44 946 INV_X1
* cell instance $55488 r0 *1 384.75,40.6
X$55488 863 787 25 44 965 OR2_X1
* cell instance $55616 m0 *1 324.33,43.4
X$55616 1003 25 44 513 BUF_X2
* cell instance $55619 m0 *1 329.65,43.4
X$55619 933 951 25 44 1038 NOR2_X1
* cell instance $55621 m0 *1 330.41,43.4
X$55621 975 891 1004 25 1039 44 AOI21_X1
* cell instance $55622 m0 *1 331.17,43.4
X$55622 951 25 44 975 INV_X1
* cell instance $55623 m0 *1 331.55,43.4
X$55623 798 933 975 44 976 25 NOR3_X2
* cell instance $55640 r0 *1 322.43,43.4
X$55640 1037 25 44 189 CLKBUF_X3
* cell instance $55644 r0 *1 330.6,43.4
X$55644 1039 970 1038 25 1005 44 AOI21_X2
* cell instance $55646 m0 *1 333.45,43.4
X$55646 952 953 976 25 1195 44 NAND3_X4
* cell instance $55652 r0 *1 334.4,43.4
X$55652 953 952 976 44 25 1040 AND3_X1
* cell instance $55655 r0 *1 335.92,43.4
X$55655 1005 898 1013 25 44 1088 OR3_X2
* cell instance $55657 m0 *1 337.82,43.4
X$55657 25 1017 895 952 953 44 AOI21_X4
* cell instance $55658 m0 *1 337.06,43.4
X$55658 952 953 895 25 44 1016 NAND3_X1
* cell instance $55662 r0 *1 337.63,43.4
X$55662 25 894 1042 896 834 1014 44 NOR4_X4
* cell instance $55666 r0 *1 343.14,43.4
X$55666 896 1017 972 44 1045 25 OAI21_X1
* cell instance $55667 m0 *1 343.71,43.4
X$55667 25 936 954 900 1046 44 NOR3_X4
* cell instance $55668 m0 *1 346.37,43.4
X$55668 900 954 936 25 44 1042 OR3_X4
* cell instance $55671 m0 *1 350.74,43.4
X$55671 955 806 977 25 44 NOR2_X4
* cell instance $55672 m0 *1 352.45,43.4
X$55672 955 806 25 1060 44 OR2_X4
* cell instance $55677 r0 *1 350.36,43.4
X$55677 977 1137 25 44 1047 XNOR2_X2
* cell instance $55680 m0 *1 356.06,43.4
X$55680 528 707 25 44 1149 XNOR2_X2
* cell instance $55682 m0 *1 361.76,43.4
X$55682 960 44 1018 25 BUF_X4
* cell instance $55692 r0 *1 362.52,43.4
X$55692 1049 579 44 1019 25 XOR2_X2
* cell instance $55695 m0 *1 364.99,43.4
X$55695 941 792 938 25 44 866 AND3_X4
* cell instance $55696 m0 *1 368.6,43.4
X$55696 25 1007 961 962 1063 44 NOR3_X4
* cell instance $55697 m0 *1 371.26,43.4
X$55697 962 961 1007 25 44 978 OR3_X4
* cell instance $55700 m0 *1 374.3,43.4
X$55700 906 979 873 963 1009 1050 44 25 AOI221_X2
* cell instance $55701 m0 *1 376.39,43.4
X$55701 941 938 25 44 979 NAND2_X2
* cell instance $55706 r0 *1 375.25,43.4
X$55706 1050 44 1020 25 BUF_X4
* cell instance $55708 r0 *1 377.34,43.4
X$55708 25 1064 779 911 938 44 AOI21_X4
* cell instance $55709 m0 *1 377.91,43.4
X$55709 973 964 941 25 44 NOR2_X4
* cell instance $55711 m0 *1 379.62,43.4
X$55711 779 25 44 964 INV_X1
* cell instance $55714 m0 *1 381.33,43.4
X$55714 1011 912 1010 44 25 938 OAI21_X4
* cell instance $55715 m0 *1 380.38,43.4
X$55715 787 810 25 44 973 NOR2_X2
* cell instance $55716 m0 *1 383.8,43.4
X$55716 826 25 44 912 INV_X2
* cell instance $55720 m0 *1 387.22,43.4
X$55720 1010 25 44 1012 INV_X1
* cell instance $55721 m0 *1 384.75,43.4
X$55721 25 908 965 826 1012 44 AOI21_X4
* cell instance $55725 r0 *1 385.51,43.4
X$55725 826 1010 25 44 1115 XNOR2_X2
* cell instance $55729 r0 *1 388.74,43.4
X$55729 25 980 1010 1214 1054 1053 44 FA_X1
* cell instance $55730 m0 *1 389.88,43.4
X$55730 913 25 44 1054 INV_X1
* cell instance $55731 m0 *1 389.5,43.4
X$55731 781 25 44 1053 INV_X1
* cell instance $55733 m0 *1 390.45,43.4
X$55733 874 25 44 980 INV_X1
* cell instance $55742 r0 *1 394.63,43.4
X$55742 875 25 44 1065 CLKBUF_X3
* cell instance $55745 m0 *1 402.04,43.4
X$55745 981 982 25 44 971 NAND2_X1
* cell instance $55748 m0 *1 404.13,43.4
X$55748 966 981 967 25 44 984 NAND3_X1
* cell instance $55749 m0 *1 402.99,43.4
X$55749 982 915 44 25 966 XNOR2_X1
* cell instance $55754 r0 *1 403.37,43.4
X$55754 1056 914 1259 25 843 44 AOI21_X1
* cell instance $55755 r0 *1 404.13,43.4
X$55755 987 967 25 44 1022 NAND2_X1
* cell instance $55756 r0 *1 404.7,43.4
X$55756 983 984 985 1024 25 44 1055 AOI22_X1
* cell instance $55757 r0 *1 405.65,43.4
X$55757 1024 985 879 916 25 44 1056 NAND4_X1
* cell instance $55761 r0 *1 409.07,43.4
X$55761 919 1097 1103 1055 44 815 25 OR4_X2
* cell instance $55764 m0 *1 414.58,43.4
X$55764 986 25 44 1008 INV_X1
* cell instance $55766 m0 *1 414.96,43.4
X$55766 940 1008 981 25 918 44 AOI21_X1
* cell instance $55767 m0 *1 415.72,43.4
X$55767 920 967 987 25 986 44 AOI21_X1
* cell instance $55768 m0 *1 416.48,43.4
X$55768 986 922 988 25 44 968 NOR3_X1
* cell instance $55769 m0 *1 417.24,43.4
X$55769 987 920 25 44 882 NOR2_X1
* cell instance $55773 m0 *1 423.13,43.4
X$55773 990 992 25 44 925 NAND2_X1
* cell instance $55777 r0 *1 415.91,43.4
X$55777 922 940 1052 44 25 1026 OAI21_X2
* cell instance $55779 r0 *1 417.43,43.4
X$55779 920 923 44 25 1051 AND2_X1
* cell instance $55780 r0 *1 418.19,43.4
X$55780 990 988 1051 25 1006 44 AOI21_X1
* cell instance $55783 r0 *1 420.85,43.4
X$55783 1028 1095 25 44 940 XNOR2_X2
* cell instance $55786 r0 *1 423.89,43.4
X$55786 992 883 991 44 25 922 AND3_X2
* cell instance $55787 m0 *1 424.27,43.4
X$55787 991 883 992 25 44 990 NAND3_X1
* cell instance $55791 m0 *1 426.74,43.4
X$55791 991 25 44 928 INV_X1
* cell instance $55795 m0 *1 431.11,43.4
X$55795 731 993 25 44 1048 NOR2_X1
* cell instance $55801 r0 *1 430.16,43.4
X$55801 994 1048 25 44 1028 XNOR2_X2
* cell instance $55802 m0 *1 432.25,43.4
X$55802 993 731 994 25 44 1002 MUX2_X1
* cell instance $55804 m0 *1 433.58,43.4
X$55804 995 993 1031 25 44 1044 NAND3_X1
* cell instance $55806 m0 *1 434.53,43.4
X$55806 996 25 44 993 INV_X1
* cell instance $55816 r0 *1 432.06,43.4
X$55816 1001 25 44 995 INV_X1
* cell instance $55817 r0 *1 432.44,43.4
X$55817 995 1000 1044 1041 1043 1286 25 44 OAI221_X2
* cell instance $55818 r0 *1 434.53,43.4
X$55818 1041 1001 1031 25 44 1043 NAND3_X1
* cell instance $55820 r0 *1 435.48,43.4
X$55820 1032 1082 731 25 44 NOR2_X4
* cell instance $55824 r0 *1 439.85,43.4
X$55824 997 1034 25 44 1031 NAND2_X2
* cell instance $55825 r0 *1 440.8,43.4
X$55825 1034 997 44 25 994 AND2_X1
* cell instance $55828 r0 *1 443.46,43.4
X$55828 999 998 1036 44 25 1034 OAI21_X2
* cell instance $55829 r0 *1 444.79,43.4
X$55829 998 999 1036 25 44 997 OR3_X2
* cell instance $56264 m0 *1 331.17,21
X$56264 189 36 25 44 503 NAND2_X1
* cell instance $56265 m0 *1 331.74,21
X$56265 360 381 420 44 25 431 HA_X1
* cell instance $56269 m0 *1 337.44,21
X$56269 382 25 44 485 INV_X1
* cell instance $56270 m0 *1 337.82,21
X$56270 422 25 44 361 INV_X1
* cell instance $56274 m0 *1 342.95,21
X$56274 25 307 468 434 385 387 44 FA_X1
* cell instance $56299 r0 *1 331.74,21
X$56299 25 380 520 432 405 420 44 FA_X1
* cell instance $56301 r0 *1 337.82,21
X$56301 433 423 422 44 25 487 HA_X1
* cell instance $56305 r0 *1 339.72,21
X$56305 406 26 44 25 423 AND2_X1
* cell instance $56309 r0 *1 341.81,21
X$56309 425 25 44 449 INV_X1
* cell instance $56313 r0 *1 346.94,21
X$56313 25 276 469 450 427 407 44 FA_X1
* cell instance $56316 m0 *1 351.12,21
X$56316 362 25 44 408 INV_X1
* cell instance $56318 m0 *1 353.21,21
X$56318 363 25 44 409 INV_X1
* cell instance $56319 m0 *1 353.59,21
X$56319 364 25 44 453 INV_X1
* cell instance $56323 m0 *1 358.72,21
X$56323 365 25 44 437 INV_X1
* cell instance $56326 m0 *1 365.94,21
X$56326 25 262 410 494 393 394 44 FA_X1
* cell instance $56327 m0 *1 368.98,21
X$56327 123 47 44 25 367 AND2_X1
* cell instance $56333 r0 *1 353.21,21
X$56333 409 453 507 44 25 509 HA_X1
* cell instance $56335 r0 *1 358.15,21
X$56335 323 40 44 25 454 AND2_X1
* cell instance $56342 r0 *1 365.75,21
X$56342 410 25 44 493 INV_X1
* cell instance $56346 r0 *1 375.44,21
X$56346 358 25 44 474 INV_X1
* cell instance $56347 m0 *1 375.82,21
X$56347 406 25 44 123 BUF_X2
* cell instance $56352 m0 *1 381.9,21
X$56352 322 25 44 411 INV_X1
* cell instance $56361 r0 *1 381.33,21
X$56361 406 301 44 25 462 AND2_X1
* cell instance $56362 r0 *1 382.09,21
X$56362 27 48 44 25 439 AND2_X1
* cell instance $56366 r0 *1 387.79,21
X$56366 38 291 44 25 465 AND2_X1
* cell instance $56374 m0 *1 395.77,21
X$56374 396 401 429 44 25 370 HA_X1
* cell instance $56376 m0 *1 397.67,21
X$56376 40 404 44 25 401 XNOR2_X1
* cell instance $56377 m0 *1 398.81,21
X$56377 265 308 47 48 25 44 404 NOR4_X1
* cell instance $56378 m0 *1 399.76,21
X$56378 265 308 25 44 415 NOR2_X1
* cell instance $56383 r0 *1 397.1,21
X$56383 429 25 44 414 INV_X1
* cell instance $56384 r0 *1 397.48,21
X$56384 414 413 428 25 412 44 AOI21_X1
* cell instance $56386 r0 *1 398.43,21
X$56386 426 25 44 428 INV_X1
* cell instance $56387 r0 *1 398.81,21
X$56387 265 301 291 47 25 44 461 NOR4_X1
* cell instance $56388 r0 *1 399.76,21
X$56388 48 461 44 25 460 XNOR2_X1
* cell instance $56389 r0 *1 400.9,21
X$56389 418 460 416 44 25 426 HA_X1
* cell instance $56391 m0 *1 405.65,21
X$56391 373 399 372 25 424 44 AOI21_X1
* cell instance $56392 m0 *1 403.75,21
X$56392 397 371 403 44 25 444 HA_X1
* cell instance $56393 m0 *1 406.41,21
X$56393 403 25 44 373 INV_X1
* cell instance $56400 r0 *1 410.97,21
X$56400 419 244 25 44 421 NAND2_X1
* cell instance $56402 r0 *1 411.92,21
X$56402 421 29 25 44 228 NAND2_X1
* cell instance $56404 m0 *1 416.67,21
X$56404 335 376 2896 44 25 391 HA_X1
* cell instance $56405 m0 *1 414.77,21
X$56405 335 375 374 44 25 417 HA_X1
* cell instance $56406 m0 *1 418.57,21
X$56406 334 25 44 270 BUF_X2
* cell instance $56408 m0 *1 419.52,21
X$56408 391 25 44 336 CLKBUF_X2
* cell instance $56411 m0 *1 421.99,21
X$56411 25 30 377 43 378 397 44 DFFR_X2
* cell instance $56467 r0 *1 416.67,21
X$56467 417 418 396 270 25 44 488 NOR4_X1
* cell instance $56712 m0 *1 342.76,15.4
X$56712 25 273 294 276 274 257 44 FA_X1
* cell instance $56715 m0 *1 348.27,15.4
X$56715 25 277 427 388 275 169 44 FA_X1
* cell instance $56720 r0 *1 343.71,15.4
X$56720 294 25 44 307 INV_X1
* cell instance $56723 r0 *1 346.37,15.4
X$56723 167 26 44 25 295 AND2_X1
* cell instance $56730 r0 *1 352.45,15.4
X$56730 243 25 44 310 INV_X1
* cell instance $56732 m0 *1 356.06,15.4
X$56732 25 245 258 365 282 125 44 FA_X1
* cell instance $56734 m0 *1 359.1,15.4
X$56734 123 40 44 25 283 AND2_X1
* cell instance $56743 r0 *1 361.38,15.4
X$56743 213 32 44 25 313 AND2_X1
* cell instance $56744 r0 *1 362.14,15.4
X$56744 25 311 296 350 314 313 44 FA_X1
* cell instance $56746 m0 *1 367.84,15.4
X$56746 25 113 262 289 351 288 44 FA_X1
* cell instance $56747 m0 *1 367.08,15.4
X$56747 36 40 44 25 261 AND2_X1
* cell instance $56748 m0 *1 370.88,15.4
X$56748 289 25 44 298 INV_X1
* cell instance $56754 m0 *1 388.74,15.4
X$56754 41 76 44 25 292 XNOR2_X1
* cell instance $56755 m0 *1 389.88,15.4
X$56755 196 292 316 44 25 225 HA_X1
* cell instance $56760 r0 *1 369.36,15.4
X$56760 25 70 297 473 218 298 44 FA_X1
* cell instance $56764 r0 *1 376.58,15.4
X$56764 167 186 44 25 319 AND2_X1
* cell instance $56765 r0 *1 377.34,15.4
X$56765 25 319 328 321 359 320 44 FA_X1
* cell instance $56766 r0 *1 380.38,15.4
X$56766 25 263 299 322 321 130 44 FA_X1
* cell instance $56769 r0 *1 385.13,15.4
X$56769 264 25 44 318 INV_X1
* cell instance $56772 r0 *1 386.65,15.4
X$56772 291 35 25 44 355 NAND2_X1
* cell instance $56773 r0 *1 387.22,15.4
X$56773 186 33 25 44 356 NAND2_X1
* cell instance $56777 r0 *1 393.11,15.4
X$56777 316 25 44 300 INV_X1
* cell instance $56781 r0 *1 395.77,15.4
X$56781 39 312 44 25 348 XNOR2_X1
* cell instance $56782 r0 *1 396.91,15.4
X$56782 309 301 291 25 44 312 NOR3_X1
* cell instance $56783 r0 *1 397.67,15.4
X$56783 25 39 308 309 76 44 NOR3_X4
* cell instance $56785 m0 *1 398.43,15.4
X$56785 48 90 40 265 44 309 25 OR4_X2
* cell instance $56786 m0 *1 399.76,15.4
X$56786 309 39 25 44 266 NOR2_X1
* cell instance $56788 m0 *1 401.09,15.4
X$56788 28 25 44 291 CLKBUF_X3
* cell instance $56792 m0 *1 412.68,15.4
X$56792 286 25 44 82 INV_X2
* cell instance $56796 m0 *1 415.72,15.4
X$56796 280 195 25 44 230 NOR2_X1
* cell instance $56798 m0 *1 417.81,15.4
X$56798 269 279 44 25 280 XNOR2_X1
* cell instance $56799 m0 *1 418.95,15.4
X$56799 272 196 229 25 44 279 NAND3_X1
* cell instance $56813 r0 *1 400.9,15.4
X$56813 301 25 44 267 INV_X2
* cell instance $56818 r0 *1 418.19,15.4
X$56818 302 303 270 25 44 81 NAND3_X2
* cell instance $56819 r0 *1 419.52,15.4
X$56819 302 303 25 44 306 NAND2_X1
* cell instance $56820 r0 *1 420.09,15.4
X$56820 302 303 270 196 25 44 234 NAND4_X1
* cell instance $56821 r0 *1 421.04,15.4
X$56821 270 306 25 44 305 XOR2_X1
* cell instance $56822 r0 *1 422.18,15.4
X$56822 305 195 25 44 304 NOR2_X1
.ENDS parameterized_freq_divider

* cell AND4_X4
* pin PWELL,VSS
* pin A4
* pin A3
* pin A2
* pin A1
* pin ZN
* pin NWELL,VDD
.SUBCKT AND4_X4 1 2 3 4 6 7 14
* net 1 PWELL,VSS
* net 2 A4
* net 3 A3
* net 4 A2
* net 6 A1
* net 7 ZN
* net 14 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 2 14 14 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 14 3 5 14 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 5 4 14 14 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 14 6 5 14 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 1.705,0.995 PMOS_VTL
M$9 7 5 14 14 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $13 r0 *1 0.185,0.2975 NMOS_VTL
M$13 8 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $14 r0 *1 0.375,0.2975 NMOS_VTL
M$14 9 3 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.565,0.2975 NMOS_VTL
M$15 10 4 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.755,0.2975 NMOS_VTL
M$16 5 6 10 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 0.945,0.2975 NMOS_VTL
M$17 12 6 5 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.135,0.2975 NMOS_VTL
M$18 11 4 12 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.325,0.2975 NMOS_VTL
M$19 13 3 11 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.515,0.2975 NMOS_VTL
M$20 1 2 13 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.705,0.2975 NMOS_VTL
M$21 7 5 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS AND4_X4

* cell OAI222_X4
* pin PWELL,VSS
* pin ZN
* pin A1
* pin A2
* pin B2
* pin B1
* pin C1
* pin C2
* pin NWELL,VDD
.SUBCKT OAI222_X4 1 5 6 7 8 9 10 11 13
* net 1 PWELL,VSS
* net 5 ZN
* net 6 A1
* net 7 A2
* net 8 B2
* net 9 B1
* net 10 C1
* net 11 C2
* net 13 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 14 6 12 13 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 13 7 14 13 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 15 8 13 13 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 12 9 15 13 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0945P PS=0.77U PD=0.93U
* device instance $5 r0 *1 1.09,0.995 PMOS_VTL
M$5 16 10 12 13 PMOS_VTL L=0.05U W=0.63U AS=0.0945P AD=0.0441P PS=0.93U PD=0.77U
* device instance $6 r0 *1 1.28,0.995 PMOS_VTL
M$6 13 11 16 13 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.47,0.995 PMOS_VTL
M$7 4 12 13 13 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 1.85,0.995 PMOS_VTL
M$9 5 4 13 13 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 12 6 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $14 r0 *1 0.36,0.2975 NMOS_VTL
M$14 2 7 12 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.55,0.2975 NMOS_VTL
M$15 3 8 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.74,0.2975 NMOS_VTL
M$16 2 9 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $17 r0 *1 1.09,0.2975 NMOS_VTL
M$17 3 10 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $18 r0 *1 1.28,0.2975 NMOS_VTL
M$18 1 11 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.47,0.2975 NMOS_VTL
M$19 4 12 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $21 r0 *1 1.85,0.2975 NMOS_VTL
M$21 5 4 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS OAI222_X4

* cell XOR2_X1
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT XOR2_X1 1 3 4 5 6
* net 1 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 8 1 2 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.555,0.995 PMOS_VTL
M$3 7 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.745,0.995 PMOS_VTL
M$4 6 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.935,0.995 PMOS_VTL
M$5 7 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 2 1 4 4 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 4 3 2 4 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.555,0.2975 NMOS_VTL
M$8 6 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.745,0.2975 NMOS_VTL
M$9 9 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.935,0.2975 NMOS_VTL
M$10 4 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XOR2_X1

* cell OAI221_X4
* pin PWELL,VSS
* pin ZN
* pin C1
* pin C2
* pin A
* pin B1
* pin B2
* pin NWELL,VDD
.SUBCKT OAI221_X4 1 5 6 7 8 9 10 12
* net 1 PWELL,VSS
* net 5 ZN
* net 6 C1
* net 7 C2
* net 8 A
* net 9 B1
* net 10 B2
* net 12 NWELL,VDD
* device instance $1 r0 *1 0.225,0.995 PMOS_VTL
M$1 13 6 11 12 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.415,0.995 PMOS_VTL
M$2 12 7 13 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.605,0.995 PMOS_VTL
M$3 11 8 12 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.051975P PS=0.77U
+ PD=0.795U
* device instance $4 r0 *1 0.82,0.995 PMOS_VTL
M$4 14 9 11 12 PMOS_VTL L=0.05U W=0.63U AS=0.051975P AD=0.083475P PS=0.795U
+ PD=0.895U
* device instance $5 r0 *1 1.135,0.995 PMOS_VTL
M$5 12 10 14 12 PMOS_VTL L=0.05U W=0.63U AS=0.083475P AD=0.0441P PS=0.895U
+ PD=0.77U
* device instance $6 r0 *1 1.325,0.995 PMOS_VTL
M$6 4 11 12 12 PMOS_VTL L=0.05U W=1.26U AS=0.096075P AD=0.096075P PS=1.565U
+ PD=1.565U
* device instance $8 r0 *1 1.73,0.995 PMOS_VTL
M$8 5 4 12 12 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $12 r0 *1 1.135,0.2975 NMOS_VTL
M$12 1 10 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $13 r0 *1 1.325,0.2975 NMOS_VTL
M$13 4 11 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0632875P AD=0.0632875P PS=1.135U
+ PD=1.135U
* device instance $15 r0 *1 1.73,0.2975 NMOS_VTL
M$15 5 4 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $19 r0 *1 0.225,0.2975 NMOS_VTL
M$19 11 6 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $20 r0 *1 0.415,0.2975 NMOS_VTL
M$20 2 7 11 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 0.605,0.2975 NMOS_VTL
M$21 3 8 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 0.795,0.2975 NMOS_VTL
M$22 1 9 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI221_X4

* cell BUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X1 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.17,0.195 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.021875P PS=0.63U PD=0.555U
* device instance $4 r0 *1 0.36,0.2975 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X1

* cell AOI221_X4
* pin PWELL,VSS
* pin ZN
* pin C1
* pin C2
* pin A
* pin B1
* pin B2
* pin NWELL,VDD
.SUBCKT AOI221_X4 1 4 7 8 9 10 11 14
* net 1 PWELL,VSS
* net 4 ZN
* net 7 C1
* net 8 C2
* net 9 A
* net 10 B1
* net 11 B2
* net 14 NWELL,VDD
* device instance $1 r0 *1 1.16,0.995 PMOS_VTL
M$1 14 11 13 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U
+ PD=0.77U
* device instance $2 r0 *1 1.35,0.995 PMOS_VTL
M$2 3 2 14 14 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $4 r0 *1 1.73,0.995 PMOS_VTL
M$4 4 3 14 14 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $8 r0 *1 0.25,0.995 PMOS_VTL
M$8 2 7 12 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $9 r0 *1 0.44,0.995 PMOS_VTL
M$9 12 8 2 14 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 0.63,0.995 PMOS_VTL
M$10 13 9 12 14 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 0.82,0.995 PMOS_VTL
M$11 14 10 13 14 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $12 r0 *1 0.25,0.2975 NMOS_VTL
M$12 5 7 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $13 r0 *1 0.44,0.2975 NMOS_VTL
M$13 1 8 5 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0342375P PS=0.555U
+ PD=0.58U
* device instance $14 r0 *1 0.655,0.2975 NMOS_VTL
M$14 2 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.0342375P AD=0.02905P PS=0.58U
+ PD=0.555U
* device instance $15 r0 *1 0.845,0.2975 NMOS_VTL
M$15 6 10 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0549875P PS=0.555U
+ PD=0.68U
* device instance $16 r0 *1 1.16,0.2975 NMOS_VTL
M$16 1 11 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.0549875P AD=0.02905P PS=0.68U
+ PD=0.555U
* device instance $17 r0 *1 1.35,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $19 r0 *1 1.73,0.2975 NMOS_VTL
M$19 4 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS AOI221_X4

* cell OR3_X4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X4 1 2 3 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.205,0.995 PMOS_VTL
M$1 11 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.395,0.995 PMOS_VTL
M$2 10 2 11 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.585,0.995 PMOS_VTL
M$3 4 3 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.775,0.995 PMOS_VTL
M$4 9 3 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.965,0.995 PMOS_VTL
M$5 8 2 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.155,0.995 PMOS_VTL
M$6 6 1 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.345,0.995 PMOS_VTL
M$7 7 4 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.177975P AD=0.200025P PS=3.085U
+ PD=3.785U
* device instance $11 r0 *1 0.205,0.2975 NMOS_VTL
M$11 4 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $12 r0 *1 0.395,0.2975 NMOS_VTL
M$12 5 2 4 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.585,0.2975 NMOS_VTL
M$13 4 3 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.345,0.2975 NMOS_VTL
M$17 7 4 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1172375P AD=0.1317625P PS=2.225U
+ PD=2.71U
.ENDS OR3_X4

* cell CLKBUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.17,0.1875 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $5 r0 *1 0.36,0.1875 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.39U AS=0.0273P AD=0.034125P PS=0.67U PD=0.935U
.ENDS CLKBUF_X2

* cell CLKBUF_X3
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X3 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.89U AS=0.1323P AD=0.15435P PS=2.31U PD=3.01U
* device instance $5 r0 *1 0.17,0.1875 NMOS_VTL
M$5 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $6 r0 *1 0.36,0.1875 NMOS_VTL
M$6 5 2 3 3 NMOS_VTL L=0.05U W=0.585U AS=0.04095P AD=0.047775P PS=1.005U
+ PD=1.27U
.ENDS CLKBUF_X3

* cell OR2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT OR2_X4 1 2 3 5 6
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 2 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 1 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 5 4 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 4 1 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $10 r0 *1 0.36,0.2975 NMOS_VTL
M$10 3 2 4 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.93,0.2975 NMOS_VTL
M$13 5 4 3 3 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS OR2_X4

* cell OR4_X4
* pin PWELL,VSS
* pin ZN
* pin A4
* pin A3
* pin A2
* pin A1
* pin NWELL,VDD
.SUBCKT OR4_X4 1 3 4 5 6 7 8
* net 1 PWELL,VSS
* net 3 ZN
* net 4 A4
* net 5 A3
* net 6 A2
* net 7 A1
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 4 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 5 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 11 6 9 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 2 7 11 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 13 7 2 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 14 6 13 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 12 5 14 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 8 4 12 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 3 2 8 8 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 4 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $14 r0 *1 0.36,0.2975 NMOS_VTL
M$14 1 5 2 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $15 r0 *1 0.55,0.2975 NMOS_VTL
M$15 2 6 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $16 r0 *1 0.74,0.2975 NMOS_VTL
M$16 1 7 2 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $21 r0 *1 1.69,0.2975 NMOS_VTL
M$21 3 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS OR4_X4

* cell AND3_X4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AND3_X4 1 2 3 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 4 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 3 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 7 4 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 11 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 10 2 11 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 4 3 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 8 3 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 9 2 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.12,0.2975 NMOS_VTL
M$16 5 1 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 1.31,0.2975 NMOS_VTL
M$17 7 4 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS AND3_X4

* cell AOI22_X2
* pin B2
* pin B1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI22_X2 1 2 3 4 5 7 8
* net 1 B2
* net 2 B1
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 7 NWELL,VDD
* net 8 ZN
* device instance $1 r0 *1 0.175,0.995 PMOS_VTL
M$1 7 1 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.365,0.995 PMOS_VTL
M$2 6 2 7 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.935,0.995 PMOS_VTL
M$5 8 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 1.125,0.995 PMOS_VTL
M$6 6 4 8 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.175,0.2975 NMOS_VTL
M$9 12 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.365,0.2975 NMOS_VTL
M$10 8 2 12 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.555,0.2975 NMOS_VTL
M$11 10 2 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.745,0.2975 NMOS_VTL
M$12 5 1 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.935,0.2975 NMOS_VTL
M$13 11 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.125,0.2975 NMOS_VTL
M$14 8 4 11 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.315,0.2975 NMOS_VTL
M$15 9 4 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.505,0.2975 NMOS_VTL
M$16 5 3 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI22_X2

* cell INV_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X1 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.06615P PS=1.47U PD=1.47U
* device instance $2 r0 *1 0.17,0.2975 NMOS_VTL
M$2 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.043575P PS=1.04U
+ PD=1.04U
.ENDS INV_X1

* cell NOR4_X2
* pin A3
* pin A2
* pin A1
* pin A4
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT NOR4_X2 1 2 3 4 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 A4
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 12 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 11 1 12 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 10 2 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 6 3 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 9 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 13 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 8 1 13 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 4 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 6 4 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 7 1 6 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $11 r0 *1 0.59,0.2975 NMOS_VTL
M$11 6 2 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 7 3 6 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS NOR4_X2

* cell OAI22_X1
* pin B2
* pin B1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI22_X1 1 2 3 4 6 7 8
* net 1 B2
* net 2 B1
* net 3 A1
* net 4 A2
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 8 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 9 3 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 6 4 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.185,0.2975 NMOS_VTL
M$5 7 1 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.375,0.2975 NMOS_VTL
M$6 5 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.565,0.2975 NMOS_VTL
M$7 8 3 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.755,0.2975 NMOS_VTL
M$8 5 4 8 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI22_X1

* cell OR2_X2
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X2 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 3 2 4 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 4 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS OR2_X2

* cell FA_X1
* pin PWELL,VSS
* pin B
* pin CO
* pin S
* pin CI
* pin A
* pin NWELL,VDD
.SUBCKT FA_X1 1 2 3 8 11 12 14
* net 1 PWELL,VSS
* net 2 B
* net 3 CO
* net 8 S
* net 11 CI
* net 12 A
* net 14 NWELL,VDD
* device instance $1 r0 *1 0.385,1.0275 PMOS_VTL
M$1 17 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $2 r0 *1 0.575,1.0275 PMOS_VTL
M$2 4 12 17 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.765,1.0275 PMOS_VTL
M$3 15 11 4 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02265P PS=0.455U
+ PD=0.535U
* device instance $4 r0 *1 0.96,1.1025 PMOS_VTL
M$4 14 12 15 14 PMOS_VTL L=0.05U W=0.315U AS=0.02265P AD=0.02205P PS=0.535U
+ PD=0.455U
* device instance $5 r0 *1 1.15,1.1025 PMOS_VTL
M$5 15 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $6 r0 *1 0.195,0.995 PMOS_VTL
M$6 14 4 3 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.033075P PS=1.47U
+ PD=0.77U
* device instance $7 r0 *1 1.49,1.1525 PMOS_VTL
M$7 16 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $8 r0 *1 1.68,1.1525 PMOS_VTL
M$8 14 11 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $9 r0 *1 1.87,1.1525 PMOS_VTL
M$9 16 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $10 r0 *1 2.06,1.1525 PMOS_VTL
M$10 7 4 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.023625P PS=0.455U
+ PD=0.465U
* device instance $11 r0 *1 2.26,1.1525 PMOS_VTL
M$11 18 11 7 14 PMOS_VTL L=0.05U W=0.315U AS=0.023625P AD=0.02205P PS=0.465U
+ PD=0.455U
* device instance $12 r0 *1 2.45,1.1525 PMOS_VTL
M$12 19 2 18 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $13 r0 *1 2.64,1.1525 PMOS_VTL
M$13 19 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $14 r0 *1 2.83,0.995 PMOS_VTL
M$14 8 7 14 14 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $15 r0 *1 0.385,0.32 NMOS_VTL
M$15 13 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.0147P PS=0.555U
+ PD=0.35U
* device instance $16 r0 *1 0.575,0.32 NMOS_VTL
M$16 4 12 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $17 r0 *1 0.765,0.32 NMOS_VTL
M$17 5 11 4 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.015225P PS=0.35U
+ PD=0.355U
* device instance $18 r0 *1 0.96,0.32 NMOS_VTL
M$18 1 12 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.015225P AD=0.0147P PS=0.355U
+ PD=0.35U
* device instance $19 r0 *1 1.15,0.32 NMOS_VTL
M$19 5 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $20 r0 *1 0.195,0.2975 NMOS_VTL
M$20 1 4 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.021875P PS=1.04U
+ PD=0.555U
* device instance $21 r0 *1 1.49,0.195 NMOS_VTL
M$21 6 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $22 r0 *1 1.68,0.195 NMOS_VTL
M$22 1 11 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $23 r0 *1 1.87,0.195 NMOS_VTL
M$23 6 12 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $24 r0 *1 2.06,0.195 NMOS_VTL
M$24 7 4 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.01575P PS=0.35U PD=0.36U
* device instance $25 r0 *1 2.26,0.195 NMOS_VTL
M$25 9 11 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.01575P AD=0.0147P PS=0.36U PD=0.35U
* device instance $26 r0 *1 2.45,0.195 NMOS_VTL
M$26 10 2 9 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $27 r0 *1 2.64,0.195 NMOS_VTL
M$27 1 12 10 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $28 r0 *1 2.83,0.2975 NMOS_VTL
M$28 8 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS FA_X1

* cell OAI221_X1
* pin B2
* pin B1
* pin A
* pin C2
* pin C1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI221_X1 1 2 3 4 5 7 8 9
* net 1 B2
* net 2 B1
* net 3 A
* net 4 C2
* net 5 C1
* net 7 NWELL,VDD
* net 8 PWELL,VSS
* net 9 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 12 1 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 12 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 9 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 11 4 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 5 11 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 8 1 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 6 2 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 10 3 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 9 4 10 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 10 5 9 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI221_X1

* cell OAI33_X1
* pin B3
* pin B2
* pin B1
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OAI33_X1 1 2 3 4 5 6 7 8 10
* net 1 B3
* net 2 B2
* net 3 B1
* net 4 A1
* net 5 A2
* net 6 A3
* net 7 PWELL,VSS
* net 8 NWELL,VDD
* net 10 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 14 1 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 13 2 14 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 10 3 13 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 12 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 11 5 12 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 8 6 11 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.185,0.2975 NMOS_VTL
M$7 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.375,0.2975 NMOS_VTL
M$8 7 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.565,0.2975 NMOS_VTL
M$9 9 3 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.755,0.2975 NMOS_VTL
M$10 10 4 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.945,0.2975 NMOS_VTL
M$11 9 5 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.135,0.2975 NMOS_VTL
M$12 10 6 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI33_X1

* cell OR3_X1
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 9 1 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 8 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 5 1 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 4 2 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 5 3 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR3_X1

* cell NOR3_X4
* pin PWELL,VSS
* pin A1
* pin A2
* pin A3
* pin ZN
* pin NWELL,VDD
.SUBCKT NOR3_X4 1 2 3 4 5 8
* net 1 PWELL,VSS
* net 2 A1
* net 3 A2
* net 4 A3
* net 5 ZN
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 5 2 7 8 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 6 3 7 8 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 1.875,0.995 PMOS_VTL
M$9 6 4 8 8 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 5 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 5 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $21 r0 *1 1.875,0.2975 NMOS_VTL
M$21 5 4 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
.ENDS NOR3_X4

* cell AND3_X2
* pin A1
* pin A2
* pin A3
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND3_X2 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 5 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 5 3 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 9 1 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 8 2 9 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 6 3 8 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 7 4 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND3_X2

* cell INV_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X2 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 4 1 2 2 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
.ENDS INV_X2

* cell INV_X4
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X4 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 2 2 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
.ENDS INV_X4

* cell AND4_X1
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND4_X1 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 6 2 5 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 5 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 5 4 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 5 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 10 1 5 7 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 11 2 10 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $8 r0 *1 0.55,0.195 NMOS_VTL
M$8 9 3 11 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.74,0.195 NMOS_VTL
M$9 7 4 9 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 8 5 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND4_X1

* cell OAI22_X4
* pin PWELL,VSS
* pin B2
* pin B1
* pin A2
* pin ZN
* pin A1
* pin NWELL,VDD
.SUBCKT OAI22_X4 1 3 4 5 6 7 8
* net 1 PWELL,VSS
* net 3 B2
* net 4 B1
* net 5 A2
* net 6 ZN
* net 7 A1
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 9 3 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 4 9 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 11 4 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 8 3 11 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 10 3 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 6 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 12 4 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 8 3 12 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 13 5 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 6 7 13 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 14 7 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 8 5 14 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $13 r0 *1 2.45,0.995 PMOS_VTL
M$13 15 5 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $14 r0 *1 2.64,0.995 PMOS_VTL
M$14 6 7 15 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $15 r0 *1 2.83,0.995 PMOS_VTL
M$15 16 7 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $16 r0 *1 3.02,0.995 PMOS_VTL
M$16 8 5 16 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 1 3 2 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $18 r0 *1 0.36,0.2975 NMOS_VTL
M$18 2 4 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
* device instance $25 r0 *1 1.69,0.2975 NMOS_VTL
M$25 6 5 2 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $26 r0 *1 1.88,0.2975 NMOS_VTL
M$26 2 7 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI22_X4

* cell XNOR2_X1
* pin A
* pin B
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT XNOR2_X1 1 2 4 5 7
* net 1 A
* net 2 B
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.18,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.37,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 7 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 8 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 4 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.18,0.195 NMOS_VTL
M$6 9 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.37,0.195 NMOS_VTL
M$7 5 2 9 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.565,0.2975 NMOS_VTL
M$8 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.755,0.2975 NMOS_VTL
M$9 7 1 6 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.945,0.2975 NMOS_VTL
M$10 6 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X1

* cell NAND4_X4
* pin PWELL,VSS
* pin A3
* pin A4
* pin A1
* pin A2
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND4_X4 1 2 3 7 8 9 10
* net 1 PWELL,VSS
* net 2 A3
* net 3 A4
* net 7 A1
* net 8 A2
* net 9 ZN
* net 10 NWELL,VDD
* device instance $1 r0 *1 0.215,0.995 PMOS_VTL
M$1 10 7 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.975,0.995 PMOS_VTL
M$5 10 8 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.22365P PS=3.08U PD=3.23U
* device instance $9 r0 *1 1.885,0.995 PMOS_VTL
M$9 10 2 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.22365P AD=0.1764P PS=3.23U PD=3.08U
* device instance $13 r0 *1 2.645,0.995 PMOS_VTL
M$13 10 3 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $17 r0 *1 1.885,0.2975 NMOS_VTL
M$17 5 2 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 2.645,0.2975 NMOS_VTL
M$21 1 3 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $25 r0 *1 0.215,0.2975 NMOS_VTL
M$25 9 7 4 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $29 r0 *1 0.975,0.2975 NMOS_VTL
M$29 5 8 4 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND4_X4

* cell NAND2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 4 1 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 5 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND2_X4

* cell NOR4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 3 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 7 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 5 4 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR4_X1

* cell NAND4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 9 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 8 3 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X1

* cell AND3_X1
* pin A1
* pin A2
* pin A3
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 4 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 4 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 8 1 4 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 9 2 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 6 3 9 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND3_X1

* cell AND4_X2
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND4_X2 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 5 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 5 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 11 1 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.36,0.2975 NMOS_VTL
M$8 10 2 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 9 3 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 7 4 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.93,0.2975 NMOS_VTL
M$11 8 5 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND4_X2

* cell AND2_X1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X1 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 7 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 5 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND2_X1

* cell AOI221_X2
* pin B1
* pin B2
* pin A
* pin C2
* pin C1
* pin ZN
* pin NWELL,VDD
* pin PWELL,VSS
.SUBCKT AOI221_X2 1 2 3 4 5 6 8 9
* net 1 B1
* net 2 B2
* net 3 A
* net 4 C2
* net 5 C1
* net 6 ZN
* net 8 NWELL,VDD
* net 9 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 3 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.09135P PS=2.24U PD=1.55U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 1 7 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 2 8 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.32,0.995 PMOS_VTL
M$7 6 4 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.09135P AD=0.11025P PS=1.55U PD=2.24U
* device instance $8 r0 *1 1.51,0.995 PMOS_VTL
M$8 10 5 6 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 6 3 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.060175P PS=1.595U
+ PD=1.12U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 14 1 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 9 2 14 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 13 2 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 6 1 13 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 1.32,0.2975 NMOS_VTL
M$17 12 4 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.031125P AD=0.02905P PS=0.565U
+ PD=0.555U
* device instance $18 r0 *1 1.51,0.2975 NMOS_VTL
M$18 6 5 12 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.7,0.2975 NMOS_VTL
M$19 11 5 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.89,0.2975 NMOS_VTL
M$20 9 4 11 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI221_X2

* cell OR3_X2
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X2 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 9 1 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 2 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 5 1 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 4 2 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 5 3 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 7 4 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS OR3_X2

* cell OAI22_X2
* pin B2
* pin B1
* pin A2
* pin A1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI22_X2 1 2 3 4 6 7 8
* net 1 B2
* net 2 B1
* net 3 A2
* net 4 A1
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 9 2 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 1 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 12 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 4 12 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 11 4 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 6 3 11 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 7 1 5 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $10 r0 *1 0.36,0.2975 NMOS_VTL
M$10 5 2 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.93,0.2975 NMOS_VTL
M$13 8 3 5 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $14 r0 *1 1.12,0.2975 NMOS_VTL
M$14 5 4 8 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI22_X2

* cell AOI22_X1
* pin B2
* pin B1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI22_X1 1 2 3 4 5 7 8
* net 1 B2
* net 2 B1
* net 3 A1
* net 4 A2
* net 5 PWELL,VSS
* net 7 NWELL,VDD
* net 8 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 7 1 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 6 2 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 8 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 6 4 8 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.185,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.375,0.2975 NMOS_VTL
M$6 8 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.565,0.2975 NMOS_VTL
M$7 9 3 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.755,0.2975 NMOS_VTL
M$8 5 4 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI22_X1

* cell NOR3_X2
* pin A3
* pin A2
* pin A1
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT NOR3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 NWELL,VDD
* net 5 ZN
* net 6 PWELL,VSS
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 10 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 9 2 10 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 5 3 9 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 8 3 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 4 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 5 1 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 6 2 5 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 5 3 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS NOR3_X2

* cell AND2_X2
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X2 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 3 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 3 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND2_X2

* cell NOR2_X4
* pin A2
* pin A1
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT NOR2_X4 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 ZN
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 9 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 3 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 8 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 1 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 3 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 6 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 1 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 3 1 4 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 4 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS NOR2_X4

* cell AOI211_X2
* pin B
* pin A
* pin C2
* pin C1
* pin ZN
* pin NWELL,VDD
* pin PWELL,VSS
.SUBCKT AOI211_X2 1 2 3 4 6 7 8
* net 1 B
* net 2 A
* net 3 C2
* net 4 C1
* net 6 ZN
* net 7 NWELL,VDD
* net 8 PWELL,VSS
* device instance $1 r0 *1 0.175,0.995 PMOS_VTL
M$1 10 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.365,0.995 PMOS_VTL
M$2 7 2 10 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.555,0.995 PMOS_VTL
M$3 9 2 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.745,0.995 PMOS_VTL
M$4 5 1 9 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.055125P PS=0.77U PD=0.805U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 6 3 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.099225P AD=0.11025P PS=1.575U PD=2.24U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 5 4 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.175,0.2975 NMOS_VTL
M$9 6 1 8 8 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0653625P PS=1.595U
+ PD=1.145U
* device instance $10 r0 *1 0.365,0.2975 NMOS_VTL
M$10 8 2 6 8 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 11 3 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.0363125P AD=0.02905P PS=0.59U
+ PD=0.555U
* device instance $14 r0 *1 1.16,0.2975 NMOS_VTL
M$14 6 4 11 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.35,0.2975 NMOS_VTL
M$15 12 4 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.54,0.2975 NMOS_VTL
M$16 8 3 12 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI211_X2

* cell AOI211_X4
* pin C1
* pin C2
* pin B
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI211_X4 1 2 3 4 8 9 10
* net 1 C1
* net 2 C2
* net 3 B
* net 4 A
* net 8 PWELL,VSS
* net 9 NWELL,VDD
* net 10 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 7 9 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 6 9 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 11 3 7 9 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 9 4 11 9 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 5 6 9 9 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 5 9 9 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 12 1 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 8 2 12 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 6 3 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 8 4 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 5 6 8 8 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.31,0.2975 NMOS_VTL
M$17 10 5 8 8 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U
+ PD=2.705U
.ENDS AOI211_X4

* cell AOI21_X2
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X2 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 7 1 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 9 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X2

* cell BUF_X8
* pin PWELL,VSS
* pin Z
* pin NWELL,VDD
* pin A
.SUBCKT BUF_X8 1 3 4 5
* net 1 PWELL,VSS
* net 3 Z
* net 4 NWELL,VDD
* net 5 A
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 5 4 4 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 3 2 4 4 PMOS_VTL L=0.05U W=5.04U AS=0.3528P AD=0.37485P PS=6.16U PD=6.86U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 5 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=3.32U AS=0.2324P AD=0.246925P PS=4.44U PD=4.925U
.ENDS BUF_X8

* cell DFFR_X2
* pin PWELL,VSS
* pin CK
* pin D
* pin RN
* pin QN
* pin Q
* pin NWELL,VDD
.SUBCKT DFFR_X2 1 3 5 9 11 12 19
* net 1 PWELL,VSS
* net 3 CK
* net 5 D
* net 9 RN
* net 11 QN
* net 12 Q
* net 19 NWELL,VDD
* device instance $1 r0 *1 2.51,1.025 PMOS_VTL
M$1 23 4 8 19 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $2 r0 *1 2.7,1.025 PMOS_VTL
M$2 23 10 19 19 PMOS_VTL L=0.05U W=0.09U AS=0.0252P AD=0.0063P PS=0.77U PD=0.23U
* device instance $3 r0 *1 1.875,1.0125 PMOS_VTL
M$3 19 6 7 19 PMOS_VTL L=0.05U W=0.315U AS=0.04725P AD=0.0322875P PS=0.93U
+ PD=0.52U
* device instance $4 r0 *1 2.13,1.0125 PMOS_VTL
M$4 22 6 19 19 PMOS_VTL L=0.05U W=0.315U AS=0.0322875P AD=0.02205P PS=0.52U
+ PD=0.455U
* device instance $5 r0 *1 2.32,1.0125 PMOS_VTL
M$5 8 2 22 19 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $6 r0 *1 2.89,0.995 PMOS_VTL
M$6 10 9 19 19 PMOS_VTL L=0.05U W=0.63U AS=0.0252P AD=0.048825P PS=0.77U
+ PD=0.785U
* device instance $7 r0 *1 3.095,0.995 PMOS_VTL
M$7 19 8 10 19 PMOS_VTL L=0.05U W=0.63U AS=0.048825P AD=0.06615P PS=0.785U
+ PD=0.84U
* device instance $8 r0 *1 3.355,0.995 PMOS_VTL
M$8 11 8 19 19 PMOS_VTL L=0.05U W=1.26U AS=0.1323P AD=0.11025P PS=1.68U PD=1.61U
* device instance $10 r0 *1 3.805,0.995 PMOS_VTL
M$10 12 10 19 19 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U
+ PD=2.24U
* device instance $12 r0 *1 1.1,1.065 PMOS_VTL
M$12 20 2 6 19 PMOS_VTL L=0.05U W=0.09U AS=0.01785P AD=0.0063P PS=0.56U PD=0.23U
* device instance $13 r0 *1 1.29,1.065 PMOS_VTL
M$13 19 7 20 19 PMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.0063P PS=0.23U PD=0.23U
* device instance $14 r0 *1 1.48,1.065 PMOS_VTL
M$14 20 9 19 19 PMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.01035P PS=0.23U
+ PD=0.41U
* device instance $15 r0 *1 0.72,1.05 PMOS_VTL
M$15 21 5 19 19 PMOS_VTL L=0.05U W=0.42U AS=0.0441P AD=0.0294P PS=1.05U PD=0.56U
* device instance $16 r0 *1 0.91,1.05 PMOS_VTL
M$16 6 4 21 19 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.01785P PS=0.56U PD=0.56U
* device instance $17 r0 *1 0.19,1.0325 PMOS_VTL
M$17 19 3 2 19 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $18 r0 *1 0.38,1.0325 PMOS_VTL
M$18 4 2 19 19 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $19 r0 *1 3.425,0.2975 NMOS_VTL
M$19 11 8 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U
+ PD=1.11U
* device instance $21 r0 *1 3.805,0.2975 NMOS_VTL
M$21 12 10 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U
+ PD=1.595U
* device instance $23 r0 *1 2.445,0.26 NMOS_VTL
M$23 18 2 8 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $24 r0 *1 2.635,0.26 NMOS_VTL
M$24 18 10 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.017675P AD=0.0063P PS=0.555U
+ PD=0.23U
* device instance $25 r0 *1 1.875,0.32 NMOS_VTL
M$25 1 6 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $26 r0 *1 2.065,0.32 NMOS_VTL
M$26 16 6 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $27 r0 *1 2.255,0.32 NMOS_VTL
M$27 8 4 16 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $28 r0 *1 2.825,0.2975 NMOS_VTL
M$28 17 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.017675P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $29 r0 *1 3.015,0.2975 NMOS_VTL
M$29 10 8 17 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $30 r0 *1 0.19,0.245 NMOS_VTL
M$30 1 3 2 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $31 r0 *1 0.38,0.245 NMOS_VTL
M$31 4 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $32 r0 *1 1.1,0.35 NMOS_VTL
M$32 15 4 6 1 NMOS_VTL L=0.05U W=0.09U AS=0.012775P AD=0.0063P PS=0.415U
+ PD=0.23U
* device instance $33 r0 *1 1.29,0.35 NMOS_VTL
M$33 14 7 15 1 NMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.0063P PS=0.23U PD=0.23U
* device instance $34 r0 *1 1.48,0.35 NMOS_VTL
M$34 1 9 14 1 NMOS_VTL L=0.05U W=0.09U AS=0.0063P AD=0.00945P PS=0.23U PD=0.39U
* device instance $35 r0 *1 0.72,0.3525 NMOS_VTL
M$35 13 5 1 1 NMOS_VTL L=0.05U W=0.275U AS=0.028875P AD=0.01925P PS=0.76U
+ PD=0.415U
* device instance $36 r0 *1 0.91,0.3525 NMOS_VTL
M$36 6 2 13 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.012775P PS=0.415U
+ PD=0.415U
.ENDS DFFR_X2

* cell HA_X1
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin CO
.SUBCKT HA_X1 1 2 4 5 6 9
* net 1 A
* net 2 B
* net 4 S
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 9 CO
* device instance $1 r0 *1 0.785,1.0275 PMOS_VTL
M$1 10 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $2 r0 *1 0.975,1.0275 PMOS_VTL
M$2 7 1 10 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $3 r0 *1 0.21,0.995 PMOS_VTL
M$3 4 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $4 r0 *1 0.4,0.995 PMOS_VTL
M$4 3 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.59,0.995 PMOS_VTL
M$5 5 7 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0338625P PS=0.77U PD=0.775U
* device instance $6 r0 *1 1.345,1.0275 PMOS_VTL
M$6 8 1 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $7 r0 *1 1.535,1.0275 PMOS_VTL
M$7 8 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $8 r0 *1 1.725,0.995 PMOS_VTL
M$8 9 8 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.345,0.195 NMOS_VTL
M$9 12 1 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $10 r0 *1 1.535,0.195 NMOS_VTL
M$10 6 2 12 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $11 r0 *1 1.725,0.2975 NMOS_VTL
M$11 9 8 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $12 r0 *1 0.785,0.195 NMOS_VTL
M$12 7 2 6 6 NMOS_VTL L=0.05U W=0.21U AS=0.0224P AD=0.0147P PS=0.56U PD=0.35U
* device instance $13 r0 *1 0.975,0.195 NMOS_VTL
M$13 6 1 7 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $14 r0 *1 0.21,0.2975 NMOS_VTL
M$14 11 2 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $15 r0 *1 0.4,0.2975 NMOS_VTL
M$15 4 1 11 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.59,0.2975 NMOS_VTL
M$16 6 7 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0224P PS=0.555U PD=0.56U
.ENDS HA_X1

* cell AOI221_X1
* pin B2
* pin B1
* pin A
* pin C2
* pin C1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI221_X1 1 2 3 4 5 6 8 9
* net 1 B2
* net 2 B1
* net 3 A
* net 4 C2
* net 5 C1
* net 6 PWELL,VSS
* net 8 NWELL,VDD
* net 9 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 7 8 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 10 3 7 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 9 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 10 5 9 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 12 1 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 9 2 12 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 6 3 9 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 11 4 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 9 5 11 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI221_X1

* cell OR4_X1
* pin A1
* pin A2
* pin A3
* pin A4
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR4_X1 1 2 3 4 5 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 5 PWELL,VSS
* net 7 NWELL,VDD
* net 8 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 10 1 6 7 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 2 10 7 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 11 3 9 7 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 11 4 7 7 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 6 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 6 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 5 2 6 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $8 r0 *1 0.55,0.195 NMOS_VTL
M$8 6 3 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.74,0.195 NMOS_VTL
M$9 5 4 6 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 8 6 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR4_X1

* cell AOI22_X4
* pin PWELL,VSS
* pin B2
* pin B1
* pin ZN
* pin A2
* pin A1
* pin NWELL,VDD
.SUBCKT AOI22_X4 1 2 3 4 5 6 16
* net 1 PWELL,VSS
* net 2 B2
* net 3 B1
* net 4 ZN
* net 5 A2
* net 6 A1
* net 16 NWELL,VDD
* device instance $1 r0 *1 0.175,0.995 PMOS_VTL
M$1 16 2 15 16 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $2 r0 *1 0.365,0.995 PMOS_VTL
M$2 15 3 16 16 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $9 r0 *1 1.695,0.995 PMOS_VTL
M$9 4 5 15 16 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $10 r0 *1 1.885,0.995 PMOS_VTL
M$10 15 6 4 16 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $17 r0 *1 0.175,0.2975 NMOS_VTL
M$17 7 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $18 r0 *1 0.365,0.2975 NMOS_VTL
M$18 4 3 7 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 0.555,0.2975 NMOS_VTL
M$19 10 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 0.745,0.2975 NMOS_VTL
M$20 1 2 10 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 0.935,0.2975 NMOS_VTL
M$21 8 2 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.125,0.2975 NMOS_VTL
M$22 4 3 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 1.315,0.2975 NMOS_VTL
M$23 12 3 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 1.505,0.2975 NMOS_VTL
M$24 1 2 12 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $25 r0 *1 1.695,0.2975 NMOS_VTL
M$25 13 5 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $26 r0 *1 1.885,0.2975 NMOS_VTL
M$26 4 6 13 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $27 r0 *1 2.075,0.2975 NMOS_VTL
M$27 11 6 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $28 r0 *1 2.265,0.2975 NMOS_VTL
M$28 1 5 11 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $29 r0 *1 2.455,0.2975 NMOS_VTL
M$29 14 5 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $30 r0 *1 2.645,0.2975 NMOS_VTL
M$30 4 6 14 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $31 r0 *1 2.835,0.2975 NMOS_VTL
M$31 9 6 4 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $32 r0 *1 3.025,0.2975 NMOS_VTL
M$32 1 5 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI22_X4

* cell OR4_X2
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OR4_X2 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 ZN
* net 8 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 11 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 10 2 11 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 9 3 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 7 5 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 5 1 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.36,0.2975 NMOS_VTL
M$8 8 2 5 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 5 3 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 8 4 5 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.93,0.2975 NMOS_VTL
M$11 7 5 8 8 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS OR4_X2

* cell MUX2_X1
* pin A
* pin S
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT MUX2_X1 1 2 3 5 6 8
* net 1 A
* net 2 S
* net 3 B
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 8 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 6 2 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 7 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 10 4 7 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $5 r0 *1 0.93,1.1525 PMOS_VTL
M$5 10 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 7 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.195 NMOS_VTL
M$7 5 2 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $8 r0 *1 0.36,0.195 NMOS_VTL
M$8 12 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.55,0.195 NMOS_VTL
M$9 7 4 12 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $10 r0 *1 0.74,0.195 NMOS_VTL
M$10 11 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $11 r0 *1 0.93,0.195 NMOS_VTL
M$11 5 3 11 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 8 7 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS MUX2_X1

* cell NOR3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 6 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 4 2 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR3_X1

* cell NAND3_X2
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 10 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 9 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 1 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X2

* cell NOR4_X4
* pin PWELL,VSS
* pin A1
* pin A2
* pin A3
* pin A4
* pin ZN
* pin NWELL,VDD
.SUBCKT NOR4_X4 1 2 3 4 5 6 10
* net 1 PWELL,VSS
* net 2 A1
* net 3 A2
* net 4 A3
* net 5 A4
* net 6 ZN
* net 10 NWELL,VDD
* device instance $1 r0 *1 1.92,0.995 PMOS_VTL
M$1 8 4 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 2.68,0.995 PMOS_VTL
M$5 10 5 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.17,0.995 PMOS_VTL
M$9 6 2 7 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $13 r0 *1 0.93,0.995 PMOS_VTL
M$13 8 3 7 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $17 r0 *1 1.92,0.2975 NMOS_VTL
M$17 1 4 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 2.68,0.2975 NMOS_VTL
M$21 1 5 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $25 r0 *1 0.17,0.2975 NMOS_VTL
M$25 6 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $29 r0 *1 0.93,0.2975 NMOS_VTL
M$29 6 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NOR4_X4

* cell OAI221_X2
* pin C2
* pin C1
* pin B1
* pin B2
* pin A
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT OAI221_X2 1 2 3 4 5 7 9 10
* net 1 C2
* net 2 C1
* net 3 B1
* net 4 B2
* net 5 A
* net 7 ZN
* net 9 PWELL,VSS
* net 10 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 12 1 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 7 2 12 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 11 2 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 10 1 11 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 5 10 10 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 14 3 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 10 4 14 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 13 4 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.73,0.995 PMOS_VTL
M$9 7 3 13 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 0.21,0.2975 NMOS_VTL
M$11 7 1 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $12 r0 *1 0.4,0.2975 NMOS_VTL
M$12 6 2 7 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $15 r0 *1 0.97,0.2975 NMOS_VTL
M$15 8 5 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $16 r0 *1 1.16,0.2975 NMOS_VTL
M$16 9 3 8 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.35,0.2975 NMOS_VTL
M$17 8 4 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI221_X2

* cell OAI21_X1
* pin B2
* pin B1
* pin A
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OAI21_X1 1 2 3 5 6 7
* net 1 B2
* net 2 B1
* net 3 A
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 6 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.575,0.995 PMOS_VTL
M$3 5 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.195,0.2975 NMOS_VTL
M$4 6 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.385,0.2975 NMOS_VTL
M$5 4 2 6 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.575,0.2975 NMOS_VTL
M$6 7 3 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X1

* cell NAND3_X4
* pin A2
* pin A1
* pin A3
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND3_X4 1 2 3 4 5 6
* net 1 A2
* net 2 A1
* net 3 A3
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 3 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 6 1 5 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $13 r0 *1 0.21,0.2975 NMOS_VTL
M$13 13 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $14 r0 *1 0.4,0.2975 NMOS_VTL
M$14 12 1 13 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.59,0.2975 NMOS_VTL
M$15 5 2 12 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.78,0.2975 NMOS_VTL
M$16 10 2 5 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 0.97,0.2975 NMOS_VTL
M$17 8 1 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.16,0.2975 NMOS_VTL
M$18 4 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.35,0.2975 NMOS_VTL
M$19 9 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.54,0.2975 NMOS_VTL
M$20 7 1 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.73,0.2975 NMOS_VTL
M$21 5 2 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.92,0.2975 NMOS_VTL
M$22 14 2 5 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.11,0.2975 NMOS_VTL
M$23 11 1 14 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.3,0.2975 NMOS_VTL
M$24 4 3 11 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X4

* cell MUX2_X2
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin Z
.SUBCKT MUX2_X2 1 2 3 6 7 8
* net 1 A
* net 2 B
* net 3 S
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 Z
* device instance $1 r0 *1 1.16,0.995 PMOS_VTL
M$1 8 4 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.077175P PS=2.24U PD=1.54U
* device instance $3 r0 *1 1.54,1.1525 PMOS_VTL
M$3 9 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $4 r0 *1 0.215,0.995 PMOS_VTL
M$4 6 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $5 r0 *1 0.405,0.995 PMOS_VTL
M$5 5 9 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 0.595,0.995 PMOS_VTL
M$6 4 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.045675P PS=0.77U PD=0.775U
* device instance $7 r0 *1 0.79,0.995 PMOS_VTL
M$7 5 3 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.045675P AD=0.0693P PS=0.775U PD=1.48U
* device instance $8 r0 *1 1.54,0.195 NMOS_VTL
M$8 9 3 7 7 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.02205P PS=0.555U PD=0.63U
* device instance $9 r0 *1 1.16,0.2975 NMOS_VTL
M$9 8 4 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.050925P PS=1.595U
+ PD=1.11U
* device instance $11 r0 *1 0.215,0.2975 NMOS_VTL
M$11 11 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.405,0.2975 NMOS_VTL
M$12 7 9 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.595,0.2975 NMOS_VTL
M$13 10 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P PS=0.555U
+ PD=0.56U
* device instance $14 r0 *1 0.79,0.2975 NMOS_VTL
M$14 4 3 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.043575P PS=0.56U
+ PD=1.04U
.ENDS MUX2_X2

* cell NAND3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 8 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X1

* cell OR2_X1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X1 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 7 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 4 1 3 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 3 2 4 3 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 4 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR2_X1

* cell XOR2_X2
* pin B
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT XOR2_X2 1 2 4 5 7
* net 1 B
* net 2 A
* net 4 NWELL,VDD
* net 5 Z
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.2,0.995 PMOS_VTL
M$1 8 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.39,0.995 PMOS_VTL
M$2 4 1 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.58,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.77,0.995 PMOS_VTL
M$4 5 2 6 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.96,0.995 PMOS_VTL
M$5 6 1 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.2,0.2975 NMOS_VTL
M$9 3 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.39,0.2975 NMOS_VTL
M$10 7 1 3 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.58,0.2975 NMOS_VTL
M$11 5 3 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $12 r0 *1 0.77,0.2975 NMOS_VTL
M$12 10 2 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.96,0.2975 NMOS_VTL
M$13 7 1 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.15,0.2975 NMOS_VTL
M$14 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.34,0.2975 NMOS_VTL
M$15 5 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
.ENDS XOR2_X2

* cell NOR2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 7 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 4 1 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.21,0.2975 NMOS_VTL
M$5 5 1 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $6 r0 *1 0.4,0.2975 NMOS_VTL
M$6 3 2 5 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS NOR2_X2

* cell NOR2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 6 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 5 2 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 5 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 3 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR2_X1

* cell OAI21_X4
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X4 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 11 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 7 3 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 5 2 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 9 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 7 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 8 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 5 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 6 1 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 7 2 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $18 r0 *1 1.12,0.2975 NMOS_VTL
M$18 4 3 7 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI21_X4

* cell NAND2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.195,0.2975 NMOS_VTL
M$5 7 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.385,0.2975 NMOS_VTL
M$6 5 2 7 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.575,0.2975 NMOS_VTL
M$7 6 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.765,0.2975 NMOS_VTL
M$8 3 1 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X2

* cell XNOR2_X2
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT XNOR2_X2 2 3 4 5 7
* net 2 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 1.135,0.995 PMOS_VTL
M$1 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 1.325,0.995 PMOS_VTL
M$2 9 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 1.515,0.995 PMOS_VTL
M$3 5 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 1.705,0.995 PMOS_VTL
M$4 8 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.18,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $7 r0 *1 0.56,0.995 PMOS_VTL
M$7 1 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 0.75,0.995 PMOS_VTL
M$8 5 2 1 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.135,0.2975 NMOS_VTL
M$9 6 2 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $11 r0 *1 1.515,0.2975 NMOS_VTL
M$11 6 3 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $13 r0 *1 0.18,0.2975 NMOS_VTL
M$13 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $15 r0 *1 0.56,0.2975 NMOS_VTL
M$15 10 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.75,0.2975 NMOS_VTL
M$16 1 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X2

* cell NAND4_X2
* pin A3
* pin A2
* pin A1
* pin A4
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND4_X2 1 2 3 4 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 A4
* net 5 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 4 7 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 7 1 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 7 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 7 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 13 4 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 12 1 13 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.59,0.2975 NMOS_VTL
M$11 11 2 12 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 6 3 11 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 8 3 6 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.16,0.2975 NMOS_VTL
M$14 10 2 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.35,0.2975 NMOS_VTL
M$15 9 1 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.54,0.2975 NMOS_VTL
M$16 5 4 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X2

* cell OAI211_X4
* pin PWELL,VSS
* pin A
* pin B
* pin C2
* pin ZN
* pin C1
* pin NWELL,VDD
.SUBCKT OAI211_X4 1 3 4 5 6 7 12
* net 1 PWELL,VSS
* net 3 A
* net 4 B
* net 5 C2
* net 6 ZN
* net 7 C1
* net 12 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 3 12 12 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 12 4 6 12 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 13 5 12 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 6 7 13 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 15 7 6 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 12 5 15 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $13 r0 *1 2.45,0.995 PMOS_VTL
M$13 14 5 12 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $14 r0 *1 2.64,0.995 PMOS_VTL
M$14 6 7 14 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $15 r0 *1 2.83,0.995 PMOS_VTL
M$15 16 7 6 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $16 r0 *1 3.02,0.995 PMOS_VTL
M$16 12 5 16 12 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 8 3 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $18 r0 *1 0.36,0.2975 NMOS_VTL
M$18 1 4 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 0.55,0.2975 NMOS_VTL
M$19 10 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 0.74,0.2975 NMOS_VTL
M$20 2 3 10 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 0.93,0.2975 NMOS_VTL
M$21 9 3 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.12,0.2975 NMOS_VTL
M$22 1 4 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 1.31,0.2975 NMOS_VTL
M$23 11 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 1.5,0.2975 NMOS_VTL
M$24 2 3 11 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $25 r0 *1 1.69,0.2975 NMOS_VTL
M$25 6 5 2 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $26 r0 *1 1.88,0.2975 NMOS_VTL
M$26 2 7 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI211_X4

* cell OAI21_X2
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X2 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 3 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 5 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 6 1 4 6 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 7 2 4 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 4 3 7 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI21_X2

* cell OAI211_X2
* pin A
* pin B
* pin C2
* pin C1
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT OAI211_X2 1 2 3 4 6 7 8
* net 1 A
* net 2 B
* net 3 C2
* net 4 C1
* net 6 ZN
* net 7 PWELL,VSS
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.205,0.995 PMOS_VTL
M$1 6 1 8 8 PMOS_VTL L=0.05U W=1.26U AS=0.111825P AD=0.0882P PS=2.245U PD=1.54U
* device instance $2 r0 *1 0.395,0.995 PMOS_VTL
M$2 8 2 6 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.089775P PS=1.54U PD=1.545U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 10 3 8 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 6 4 10 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 9 4 6 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 8 3 9 8 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.205,0.2975 NMOS_VTL
M$9 12 1 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.395,0.2975 NMOS_VTL
M$10 7 2 12 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.585,0.2975 NMOS_VTL
M$11 11 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P PS=0.555U
+ PD=0.56U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 5 1 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.02905P PS=0.56U
+ PD=0.555U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 6 3 5 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $14 r0 *1 1.16,0.2975 NMOS_VTL
M$14 5 4 6 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI211_X2

* cell NAND2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 6 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 5 2 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X1

* cell AOI21_X4
* pin PWELL,VSS
* pin ZN
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
.SUBCKT AOI21_X4 1 2 3 4 5 11
* net 1 PWELL,VSS
* net 2 ZN
* net 3 A
* net 4 B2
* net 5 B1
* net 11 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 11 3 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 2 4 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 10 5 2 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $13 r0 *1 0.185,0.2975 NMOS_VTL
M$13 2 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.945,0.2975 NMOS_VTL
M$17 8 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.135,0.2975 NMOS_VTL
M$18 2 5 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.325,0.2975 NMOS_VTL
M$19 9 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.515,0.2975 NMOS_VTL
M$20 1 4 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.705,0.2975 NMOS_VTL
M$21 6 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.895,0.2975 NMOS_VTL
M$22 2 5 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.085,0.2975 NMOS_VTL
M$23 7 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.275,0.2975 NMOS_VTL
M$24 1 4 7 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X4

* cell BUF_X4
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT BUF_X4 1 3 4 5
* net 1 A
* net 3 NWELL,VDD
* net 4 Z
* net 5 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 2 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 4 2 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS BUF_X4

* cell AOI21_X1
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X1 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 2 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 7 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 8 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 6 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.59,0.2975 NMOS_VTL
M$6 4 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X1

* cell BUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS BUF_X2
