module parameterized_clock_gating (clk_in,
    clk_out,
    enable,
    test_mode);
 input clk_in;
 output clk_out;
 input enable;
 input test_mode;

 wire _0_;
 wire enable_final;
 wire enable_latch;
 wire \gen_sync.enable_sync_reg[0] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;

 sky130_fd_sc_hd__or2_0 _1_ (.A(net3),
    .B(enable_final),
    .X(_0_));
 sky130_fd_sc_hd__and2_0 _2_ (.A(enable_latch),
    .B(net1),
    .X(net4));
 sky130_fd_sc_hd__dlxtn_1 \enable_latch$_DLATCH_N_  (.D(_0_),
    .Q(enable_latch),
    .GATE_N(net1));
 sky130_fd_sc_hd__dfxtp_1 \gen_sync.enable_sync_reg[0]$_DFF_P_  (.D(net2),
    .Q(\gen_sync.enable_sync_reg[0] ),
    .CLK(net1));
 sky130_fd_sc_hd__dfxtp_1 \gen_sync.enable_sync_reg[1]$_DFF_P_  (.D(\gen_sync.enable_sync_reg[0] ),
    .Q(enable_final),
    .CLK(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_146 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(clk_in),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(enable),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(test_mode),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 output4 (.A(net4),
    .X(clk_out));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
endmodule
