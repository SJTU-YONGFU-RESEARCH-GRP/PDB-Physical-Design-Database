module fair_priority_arbiter (clk,
    rst_n,
    valid,
    grant,
    grant_idx,
    priorities,
    request);
 input clk;
 input rst_n;
 output valid;
 output [3:0] grant;
 output [1:0] grant_idx;
 input [7:0] priorities;
 input [3:0] request;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire net1;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net74;
 wire net75;
 wire net76;
 wire net37;
 wire net38;

 sky130_fd_sc_hd__a222oi_1 _132_ (.A1(net8),
    .A2(_108_),
    .B1(_120_),
    .B2(net6),
    .C1(_116_),
    .C2(net10),
    .Y(_053_));
 sky130_fd_sc_hd__inv_1 _133_ (.A(net4),
    .Y(_054_));
 sky130_fd_sc_hd__mux2i_4 _134_ (.A0(_053_),
    .A1(_054_),
    .S(_114_),
    .Y(_055_));
 sky130_fd_sc_hd__inv_1 _135_ (.A(_055_),
    .Y(_103_));
 sky130_fd_sc_hd__buf_2 _136_ (.A(request[1]),
    .X(_056_));
 sky130_fd_sc_hd__buf_2 _137_ (.A(request[3]),
    .X(_057_));
 sky130_fd_sc_hd__dlymetal6s2s_1 split1 (.A(net23),
    .X(net1));
 sky130_fd_sc_hd__mux2i_1 _139_ (.A0(_056_),
    .A1(_057_),
    .S(_109_),
    .Y(_059_));
 sky130_fd_sc_hd__mux2i_1 _140_ (.A0(net12),
    .A1(net13),
    .S(_109_),
    .Y(_060_));
 sky130_fd_sc_hd__or2_4 _141_ (.A(_122_),
    .B(net21),
    .X(_061_));
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__mux2_4 _143_ (.A0(_059_),
    .A1(_060_),
    .S(_061_),
    .X(_063_));
 sky130_fd_sc_hd__a222oi_1 _144_ (.A1(_112_),
    .A2(net11),
    .B1(net9),
    .B2(_116_),
    .C1(net7),
    .C2(_108_),
    .Y(_064_));
 sky130_fd_sc_hd__nand2_1 _145_ (.A(net36),
    .B(net5),
    .Y(_065_));
 sky130_fd_sc_hd__o21ai_1 _146_ (.A1(net36),
    .A2(_064_),
    .B1(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__nand2b_4 _147_ (.A_N(_063_),
    .B(_066_),
    .Y(_099_));
 sky130_fd_sc_hd__a222oi_1 _148_ (.A1(net11),
    .A2(_110_),
    .B1(_112_),
    .B2(net7),
    .C1(_120_),
    .C2(net9),
    .Y(_067_));
 sky130_fd_sc_hd__inv_1 _149_ (.A(net5),
    .Y(_068_));
 sky130_fd_sc_hd__mux2_1 _150_ (.A0(_067_),
    .A1(_068_),
    .S(_118_),
    .X(_124_));
 sky130_fd_sc_hd__inv_1 _151_ (.A(_110_),
    .Y(_069_));
 sky130_fd_sc_hd__a222oi_1 _152_ (.A1(net9),
    .A2(_112_),
    .B1(_116_),
    .B2(net7),
    .C1(_120_),
    .C2(net11),
    .Y(_070_));
 sky130_fd_sc_hd__nand2_1 _153_ (.A(_069_),
    .B(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__o21ai_0 _154_ (.A1(net5),
    .A2(_069_),
    .B1(_071_),
    .Y(_128_));
 sky130_fd_sc_hd__buf_2 _155_ (.A(_109_),
    .X(_072_));
 sky130_fd_sc_hd__mux4_1 _156_ (.A0(net12),
    .A1(net13),
    .A2(_057_),
    .A3(_056_),
    .S0(_072_),
    .S1(_061_),
    .X(_073_));
 sky130_fd_sc_hd__nand2b_1 _157_ (.A_N(_057_),
    .B(_109_),
    .Y(_074_));
 sky130_fd_sc_hd__o21bai_1 _158_ (.A1(net2),
    .A2(net1),
    .B1_N(_072_),
    .Y(_075_));
 sky130_fd_sc_hd__o22ai_1 _159_ (.A1(_061_),
    .A2(_074_),
    .B1(_075_),
    .B2(net13),
    .Y(_076_));
 sky130_fd_sc_hd__nor2_1 _160_ (.A(net12),
    .B(_056_),
    .Y(_077_));
 sky130_fd_sc_hd__or4_1 _161_ (.A(_056_),
    .B(net2),
    .C(net1),
    .D(_109_),
    .X(_078_));
 sky130_fd_sc_hd__o21ai_1 _162_ (.A1(net2),
    .A2(net1),
    .B1(_072_),
    .Y(_079_));
 sky130_fd_sc_hd__or3_1 _163_ (.A(net12),
    .B(net13),
    .C(_057_),
    .X(_080_));
 sky130_fd_sc_hd__o32ai_2 _164_ (.A1(net13),
    .A2(_057_),
    .A3(_078_),
    .B1(_079_),
    .B2(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__a21oi_1 _165_ (.A1(_076_),
    .A2(_077_),
    .B1(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__nor2_1 _166_ (.A(_073_),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__inv_1 _167_ (.A(_083_),
    .Y(_004_));
 sky130_fd_sc_hd__nor2_2 _168_ (.A(net2),
    .B(net22),
    .Y(_084_));
 sky130_fd_sc_hd__mux4_2 _169_ (.A0(_056_),
    .A1(net13),
    .A2(_057_),
    .A3(net12),
    .S0(_084_),
    .S1(_109_),
    .X(_085_));
 sky130_fd_sc_hd__nor2b_4 _170_ (.A(_104_),
    .B_N(_101_),
    .Y(_086_));
 sky130_fd_sc_hd__a2bb2oi_2 _171_ (.A1_N(_086_),
    .A2_N(_100_),
    .B1(net34),
    .B2(_105_),
    .Y(_087_));
 sky130_fd_sc_hd__a222oi_1 _172_ (.A1(net10),
    .A2(_112_),
    .B1(_116_),
    .B2(net8),
    .C1(net6),
    .C2(_108_),
    .Y(_088_));
 sky130_fd_sc_hd__and2b_2 _173_ (.A_N(net36),
    .B(_088_),
    .X(_089_));
 sky130_fd_sc_hd__nor2b_1 _174_ (.A(net4),
    .B_N(net36),
    .Y(_090_));
 sky130_fd_sc_hd__a2111oi_2 _175_ (.A1(_085_),
    .A2(net31),
    .B1(_063_),
    .C1(_089_),
    .D1(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__o21a_2 _176_ (.A1(_087_),
    .A2(_063_),
    .B1(_085_),
    .X(_092_));
 sky130_fd_sc_hd__nor3_4 _177_ (.A(_063_),
    .B(_089_),
    .C(_090_),
    .Y(_102_));
 sky130_fd_sc_hd__o22ai_4 _178_ (.A1(_055_),
    .A2(_091_),
    .B1(_092_),
    .B2(net75),
    .Y(_093_));
 sky130_fd_sc_hd__inv_1 _179_ (.A(net13),
    .Y(_094_));
 sky130_fd_sc_hd__o21ai_1 _180_ (.A1(_057_),
    .A2(_079_),
    .B1(_078_),
    .Y(_095_));
 sky130_fd_sc_hd__o22ai_2 _181_ (.A1(_061_),
    .A2(_074_),
    .B1(_075_),
    .B2(_056_),
    .Y(_096_));
 sky130_fd_sc_hd__inv_1 _182_ (.A(net12),
    .Y(_097_));
 sky130_fd_sc_hd__nor2_4 _183_ (.A(_126_),
    .B(_127_),
    .Y(_007_));
 sky130_fd_sc_hd__a221oi_4 _184_ (.A1(_094_),
    .A2(_095_),
    .B1(_096_),
    .B2(_097_),
    .C1(_007_),
    .Y(_008_));
 sky130_fd_sc_hd__mux4_1 _185_ (.A0(net13),
    .A1(_057_),
    .A2(net12),
    .A3(_056_),
    .S0(_084_),
    .S1(_072_),
    .X(_009_));
 sky130_fd_sc_hd__inv_1 _186_ (.A(_009_),
    .Y(_010_));
 sky130_fd_sc_hd__nor2_1 _187_ (.A(_131_),
    .B(_130_),
    .Y(_011_));
 sky130_fd_sc_hd__a211oi_2 _188_ (.A1(_076_),
    .A2(_077_),
    .B1(_081_),
    .C1(_011_),
    .Y(_012_));
 sky130_fd_sc_hd__o21ai_1 _189_ (.A1(_008_),
    .A2(_010_),
    .B1(_012_),
    .Y(_013_));
 sky130_fd_sc_hd__a222oi_1 _190_ (.A1(net10),
    .A2(_110_),
    .B1(_112_),
    .B2(net6),
    .C1(_120_),
    .C2(net8),
    .Y(_014_));
 sky130_fd_sc_hd__mux2i_2 _191_ (.A0(_014_),
    .A1(_054_),
    .S(_118_),
    .Y(_015_));
 sky130_fd_sc_hd__a222oi_1 _192_ (.A1(net8),
    .A2(_112_),
    .B1(_116_),
    .B2(net6),
    .C1(_120_),
    .C2(net10),
    .Y(_016_));
 sky130_fd_sc_hd__nor2b_1 _193_ (.A(net4),
    .B_N(_110_),
    .Y(_017_));
 sky130_fd_sc_hd__a211o_1 _194_ (.A1(_069_),
    .A2(_016_),
    .B1(_017_),
    .C1(_130_),
    .X(_018_));
 sky130_fd_sc_hd__a21o_1 _195_ (.A1(_015_),
    .A2(_009_),
    .B1(_018_),
    .X(_019_));
 sky130_fd_sc_hd__inv_1 _196_ (.A(_126_),
    .Y(_020_));
 sky130_fd_sc_hd__a2111o_1 _197_ (.A1(_069_),
    .A2(_016_),
    .B1(_017_),
    .C1(_130_),
    .D1(_020_),
    .X(_021_));
 sky130_fd_sc_hd__a221o_1 _198_ (.A1(_094_),
    .A2(_095_),
    .B1(_096_),
    .B2(_097_),
    .C1(_021_),
    .X(_022_));
 sky130_fd_sc_hd__nand3_2 _199_ (.A(_012_),
    .B(_022_),
    .C(_019_),
    .Y(_023_));
 sky130_fd_sc_hd__o211ai_2 _200_ (.A1(_013_),
    .A2(_093_),
    .B1(_073_),
    .C1(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__and2_0 _201_ (.A(_020_),
    .B(_015_),
    .X(_025_));
 sky130_fd_sc_hd__a21boi_0 _202_ (.A1(_093_),
    .A2(_025_),
    .B1_N(_008_),
    .Y(_026_));
 sky130_fd_sc_hd__nor2_1 _203_ (.A(_072_),
    .B(_084_),
    .Y(_027_));
 sky130_fd_sc_hd__nor2b_1 _204_ (.A(net30),
    .B_N(_057_),
    .Y(_028_));
 sky130_fd_sc_hd__nor3_1 _205_ (.A(_097_),
    .B(_061_),
    .C(_028_),
    .Y(_029_));
 sky130_fd_sc_hd__o21ai_1 _206_ (.A1(_063_),
    .A2(net30),
    .B1(_085_),
    .Y(_030_));
 sky130_fd_sc_hd__a221oi_1 _207_ (.A1(_056_),
    .A2(_027_),
    .B1(_029_),
    .B2(_072_),
    .C1(_030_),
    .Y(_031_));
 sky130_fd_sc_hd__o21ai_1 _208_ (.A1(_026_),
    .A2(_010_),
    .B1(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__nor2_1 _209_ (.A(_010_),
    .B(_008_),
    .Y(_033_));
 sky130_fd_sc_hd__a41o_1 _210_ (.A1(_020_),
    .A2(_093_),
    .A3(_015_),
    .A4(_009_),
    .B1(_033_),
    .X(_034_));
 sky130_fd_sc_hd__nand2_1 _211_ (.A(_057_),
    .B(_084_),
    .Y(_035_));
 sky130_fd_sc_hd__o21ai_0 _212_ (.A1(_094_),
    .A2(_084_),
    .B1(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__nand2_1 _213_ (.A(_072_),
    .B(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__nand2b_1 _214_ (.A_N(_072_),
    .B(_036_),
    .Y(_038_));
 sky130_fd_sc_hd__o32a_1 _215_ (.A1(_034_),
    .A2(_029_),
    .A3(_037_),
    .B1(_038_),
    .B2(_026_),
    .X(_039_));
 sky130_fd_sc_hd__nand3_1 _216_ (.A(_056_),
    .B(_072_),
    .C(net35),
    .Y(_040_));
 sky130_fd_sc_hd__o31ai_2 _217_ (.A1(_097_),
    .A2(_072_),
    .A3(net35),
    .B1(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__o2bb2ai_1 _218_ (.A1_N(_019_),
    .A2_N(_022_),
    .B1(_033_),
    .B2(_093_),
    .Y(_042_));
 sky130_fd_sc_hd__nand2_1 _219_ (.A(_012_),
    .B(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__a32oi_4 _220_ (.A1(net37),
    .A2(_032_),
    .A3(_039_),
    .B1(_041_),
    .B2(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__nor2_1 _221_ (.A(_059_),
    .B(_092_),
    .Y(_045_));
 sky130_fd_sc_hd__o21a_1 _222_ (.A1(_034_),
    .A2(_045_),
    .B1(_024_),
    .X(_046_));
 sky130_fd_sc_hd__o21ai_1 _223_ (.A1(_030_),
    .A2(_034_),
    .B1(_024_),
    .Y(_047_));
 sky130_fd_sc_hd__mux2_4 _224_ (.A0(_046_),
    .A1(_047_),
    .S(net35),
    .X(_048_));
 sky130_fd_sc_hd__nor3_2 _225_ (.A(_083_),
    .B(_048_),
    .C(_044_),
    .Y(_000_));
 sky130_fd_sc_hd__mux2i_2 _226_ (.A0(_046_),
    .A1(_047_),
    .S(net35),
    .Y(_049_));
 sky130_fd_sc_hd__nor2_1 _227_ (.A(_049_),
    .B(_044_),
    .Y(_001_));
 sky130_fd_sc_hd__and2_4 _228_ (.A(_049_),
    .B(_044_),
    .X(_002_));
 sky130_fd_sc_hd__and2_4 _229_ (.A(_048_),
    .B(_044_),
    .X(_003_));
 sky130_fd_sc_hd__a222oi_1 _230_ (.A1(net9),
    .A2(_108_),
    .B1(_120_),
    .B2(net7),
    .C1(_116_),
    .C2(net11),
    .Y(_050_));
 sky130_fd_sc_hd__mux2i_2 _231_ (.A0(_050_),
    .A1(_068_),
    .S(_114_),
    .Y(_098_));
 sky130_fd_sc_hd__inv_4 _232_ (.A(net18),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _233_ (.A(net19),
    .Y(_107_));
 sky130_fd_sc_hd__nand2_2 _234_ (.A(_092_),
    .B(_098_),
    .Y(_051_));
 sky130_fd_sc_hd__o21ai_4 _235_ (.A1(_092_),
    .A2(_099_),
    .B1(_051_),
    .Y(_125_));
 sky130_fd_sc_hd__nor2_1 _236_ (.A(_034_),
    .B(_125_),
    .Y(_052_));
 sky130_fd_sc_hd__a21oi_1 _237_ (.A1(_124_),
    .A2(_034_),
    .B1(_052_),
    .Y(_129_));
 sky130_fd_sc_hd__o21ai_1 _238_ (.A1(_106_),
    .A2(_004_),
    .B1(_049_),
    .Y(_005_));
 sky130_fd_sc_hd__a21o_1 _239_ (.A1(net25),
    .A2(_083_),
    .B1(_044_),
    .X(_006_));
 sky130_fd_sc_hd__ha_4 _240_ (.A(_099_),
    .B(_098_),
    .COUT(_100_),
    .SUM(_101_));
 sky130_fd_sc_hd__ha_2 _241_ (.A(_102_),
    .B(_103_),
    .COUT(_104_),
    .SUM(_105_));
 sky130_fd_sc_hd__ha_4 _242_ (.A(_106_),
    .B(_107_),
    .COUT(_108_),
    .SUM(_109_));
 sky130_fd_sc_hd__ha_1 _243_ (.A(_106_),
    .B(_107_),
    .COUT(_110_),
    .SUM(_111_));
 sky130_fd_sc_hd__ha_4 _244_ (.A(_106_),
    .B(net26),
    .COUT(_112_),
    .SUM(_113_));
 sky130_fd_sc_hd__ha_2 _245_ (.A(_106_),
    .B(net27),
    .COUT(_114_),
    .SUM(_115_));
 sky130_fd_sc_hd__ha_2 _246_ (.A(net24),
    .B(_107_),
    .COUT(_116_),
    .SUM(_117_));
 sky130_fd_sc_hd__ha_1 _247_ (.A(net1),
    .B(_107_),
    .COUT(_118_),
    .SUM(_119_));
 sky130_fd_sc_hd__ha_2 _248_ (.A(net33),
    .B(net26),
    .COUT(_120_),
    .SUM(_121_));
 sky130_fd_sc_hd__ha_4 _249_ (.A(net19),
    .B(net18),
    .COUT(_122_),
    .SUM(_123_));
 sky130_fd_sc_hd__ha_4 _250_ (.A(_125_),
    .B(_124_),
    .COUT(_126_),
    .SUM(_127_));
 sky130_fd_sc_hd__ha_2 _251_ (.A(_128_),
    .B(_129_),
    .COUT(_130_),
    .SUM(_131_));
 sky130_fd_sc_hd__dfrtp_1 \grant[0]$_DFF_PN0_  (.D(_000_),
    .Q(net14),
    .RESET_B(net3),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \grant[1]$_DFF_PN0_  (.D(_001_),
    .Q(net15),
    .RESET_B(net3),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \grant[2]$_DFF_PN0_  (.D(_002_),
    .Q(net16),
    .RESET_B(net3),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \grant[3]$_DFF_PN0_  (.D(_003_),
    .Q(net17),
    .RESET_B(net3),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \last_grant_idx[0]$_DFFE_PN0P_  (.D(_005_),
    .Q(net18),
    .RESET_B(net3),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \last_grant_idx[1]$_DFFE_PN0P_  (.D(_006_),
    .Q(net19),
    .RESET_B(net3),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid$_DFF_PN0_  (.D(_004_),
    .Q(net20),
    .RESET_B(net3),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlymetal6s2s_1 split2 (.A(_122_),
    .X(net2));
 sky130_fd_sc_hd__buf_2 hold3 (.A(net76),
    .X(net3));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_49 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(priorities[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(priorities[1]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(priorities[2]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(priorities[3]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(priorities[4]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(priorities[5]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(priorities[6]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(priorities[7]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(request[0]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(request[2]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net14),
    .X(grant[0]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net15),
    .X(grant[1]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net16),
    .X(grant[2]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net17),
    .X(grant[3]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net32),
    .X(grant_idx[0]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net28),
    .X(grant_idx[1]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net20),
    .X(valid));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__buf_6 rebuffer1 (.A(net18),
    .X(net21));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net21),
    .X(net22));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net22),
    .X(net23));
 sky130_fd_sc_hd__buf_1 rebuffer4 (.A(net21),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net19),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 rebuffer6 (.A(net19),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net26),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net19),
    .X(net28));
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(_087_),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(_087_),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net57),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net18),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer14 (.A(_101_),
    .X(net34));
 sky130_fd_sc_hd__buf_2 clone15 (.A(_061_),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(_122_),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net74),
    .X(net70));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__clkbuf_2 rebuffer54 (.A(net38),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(_102_),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(rst_n),
    .X(net76));
 sky130_fd_sc_hd__buf_2 rebuffer15 (.A(_024_),
    .X(net37));
 sky130_fd_sc_hd__buf_6 rebuffer17 (.A(net18),
    .X(net38));
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_142 ();
endmodule
