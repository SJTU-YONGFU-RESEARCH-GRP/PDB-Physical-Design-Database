module shift_register_left (clk,
    en,
    load,
    rst_n,
    serial_in,
    serial_out,
    parallel_in,
    parallel_out);
 input clk;
 input en;
 input load;
 input rst_n;
 input serial_in;
 output serial_out;
 input [7:0] parallel_in;
 output [7:0] parallel_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net21;

 sky130_fd_sc_hd__buf_6 _26_ (.A(net2),
    .X(_08_));
 sky130_fd_sc_hd__buf_6 _27_ (.A(en),
    .X(_09_));
 sky130_fd_sc_hd__mux2i_1 _28_ (.A0(net12),
    .A1(net11),
    .S(_09_),
    .Y(_10_));
 sky130_fd_sc_hd__nand2_1 _29_ (.A(_08_),
    .B(net3),
    .Y(_11_));
 sky130_fd_sc_hd__o21ai_0 _30_ (.A1(_08_),
    .A2(_10_),
    .B1(_11_),
    .Y(_00_));
 sky130_fd_sc_hd__mux2i_1 _31_ (.A0(net13),
    .A1(net12),
    .S(_09_),
    .Y(_12_));
 sky130_fd_sc_hd__nand2_1 _32_ (.A(_08_),
    .B(net4),
    .Y(_13_));
 sky130_fd_sc_hd__o21ai_0 _33_ (.A1(_08_),
    .A2(_12_),
    .B1(_13_),
    .Y(_01_));
 sky130_fd_sc_hd__mux2i_1 _34_ (.A0(net14),
    .A1(net13),
    .S(_09_),
    .Y(_14_));
 sky130_fd_sc_hd__nand2_1 _35_ (.A(_08_),
    .B(net5),
    .Y(_15_));
 sky130_fd_sc_hd__o21ai_0 _36_ (.A1(net2),
    .A2(_14_),
    .B1(_15_),
    .Y(_02_));
 sky130_fd_sc_hd__mux2i_1 _37_ (.A0(net15),
    .A1(net14),
    .S(_09_),
    .Y(_16_));
 sky130_fd_sc_hd__nand2_1 _38_ (.A(_08_),
    .B(net6),
    .Y(_17_));
 sky130_fd_sc_hd__o21ai_0 _39_ (.A1(net2),
    .A2(_16_),
    .B1(_17_),
    .Y(_03_));
 sky130_fd_sc_hd__mux2i_1 _40_ (.A0(net16),
    .A1(net15),
    .S(_09_),
    .Y(_18_));
 sky130_fd_sc_hd__nand2_1 _41_ (.A(_08_),
    .B(net7),
    .Y(_19_));
 sky130_fd_sc_hd__o21ai_0 _42_ (.A1(net2),
    .A2(_18_),
    .B1(_19_),
    .Y(_04_));
 sky130_fd_sc_hd__mux2i_1 _43_ (.A0(net17),
    .A1(net16),
    .S(_09_),
    .Y(_20_));
 sky130_fd_sc_hd__nand2_1 _44_ (.A(_08_),
    .B(net8),
    .Y(_21_));
 sky130_fd_sc_hd__o21ai_0 _45_ (.A1(net2),
    .A2(_20_),
    .B1(_21_),
    .Y(_05_));
 sky130_fd_sc_hd__mux2i_1 _46_ (.A0(net18),
    .A1(net17),
    .S(_09_),
    .Y(_22_));
 sky130_fd_sc_hd__nand2_1 _47_ (.A(_08_),
    .B(net9),
    .Y(_23_));
 sky130_fd_sc_hd__o21ai_0 _48_ (.A1(net2),
    .A2(_22_),
    .B1(_23_),
    .Y(_06_));
 sky130_fd_sc_hd__mux2i_1 _49_ (.A0(net20),
    .A1(net18),
    .S(_09_),
    .Y(_24_));
 sky130_fd_sc_hd__nand2_1 _50_ (.A(_08_),
    .B(net10),
    .Y(_25_));
 sky130_fd_sc_hd__o21ai_0 _51_ (.A1(net2),
    .A2(_24_),
    .B1(_25_),
    .Y(_07_));
 sky130_fd_sc_hd__clkbuf_1 _52_ (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[0]$_DFFE_PN0P_  (.D(_00_),
    .Q(net12),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[1]$_DFFE_PN0P_  (.D(_01_),
    .Q(net13),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[2]$_DFFE_PN0P_  (.D(_02_),
    .Q(net14),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[3]$_DFFE_PN0P_  (.D(_03_),
    .Q(net15),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[4]$_DFFE_PN0P_  (.D(_04_),
    .Q(net16),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[5]$_DFFE_PN0P_  (.D(_05_),
    .Q(net17),
    .RESET_B(net1),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[6]$_DFFE_PN0P_  (.D(_06_),
    .Q(net18),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \parallel_out[7]$_DFFE_PN0P_  (.D(_07_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 hold1 (.A(net21),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_24 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(load),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(parallel_in[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(parallel_in[1]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(parallel_in[2]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(parallel_in[3]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(parallel_in[4]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(parallel_in[5]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(parallel_in[6]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(parallel_in[7]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(serial_in),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net12),
    .X(parallel_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(parallel_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(parallel_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(parallel_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(parallel_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(parallel_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(parallel_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(parallel_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(serial_out));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net21));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_91 ();
endmodule
