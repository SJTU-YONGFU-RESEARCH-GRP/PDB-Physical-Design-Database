module parameterized_johnson_updown_counter (clk,
    enable,
    rst_n,
    up_down,
    count);
 input clk;
 input enable;
 input rst_n;
 input up_down;
 output [3:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X4 _23_ (.A(enable),
    .Z(_06_));
 OAI21_X1 _24_ (.A(net1),
    .B1(_06_),
    .B2(net2),
    .ZN(_07_));
 BUF_X4 _25_ (.A(up_down),
    .Z(_08_));
 MUX2_X1 _26_ (.A(_00_),
    .B(net3),
    .S(_08_),
    .Z(_09_));
 INV_X1 _27_ (.A(_09_),
    .ZN(_10_));
 AOI21_X1 _28_ (.A(_07_),
    .B1(_10_),
    .B2(_06_),
    .ZN(_02_));
 OAI21_X1 _29_ (.A(net1),
    .B1(_06_),
    .B2(net3),
    .ZN(_11_));
 MUX2_X1 _30_ (.A(net2),
    .B(net4),
    .S(_08_),
    .Z(_12_));
 INV_X1 _31_ (.A(_12_),
    .ZN(_13_));
 AOI21_X1 _32_ (.A(_11_),
    .B1(_13_),
    .B2(_06_),
    .ZN(_03_));
 OAI21_X1 _33_ (.A(net1),
    .B1(_06_),
    .B2(net4),
    .ZN(_14_));
 MUX2_X1 _34_ (.A(net3),
    .B(net5),
    .S(_08_),
    .Z(_15_));
 INV_X1 _35_ (.A(_15_),
    .ZN(_16_));
 AOI21_X1 _36_ (.A(_14_),
    .B1(_16_),
    .B2(_06_),
    .ZN(_04_));
 NOR2_X1 _37_ (.A1(net5),
    .A2(_06_),
    .ZN(_17_));
 INV_X1 _38_ (.A(_06_),
    .ZN(_18_));
 MUX2_X1 _39_ (.A(net4),
    .B(_01_),
    .S(_08_),
    .Z(_19_));
 NOR2_X1 _40_ (.A1(_18_),
    .A2(_19_),
    .ZN(_20_));
 OAI21_X1 _41_ (.A(net1),
    .B1(_17_),
    .B2(_20_),
    .ZN(_05_));
 DFF_X1 \counter_reg[0]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net2),
    .QN(_01_));
 DFF_X1 \counter_reg[1]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net3),
    .QN(_22_));
 DFF_X1 \counter_reg[2]$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net4),
    .QN(_21_));
 DFF_X1 \counter_reg[3]$_SDFFE_PN1P_  (.D(_05_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net5),
    .QN(_00_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_63 ();
 BUF_X1 input1 (.A(rst_n),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(count[0]));
 BUF_X1 output3 (.A(net3),
    .Z(count[1]));
 BUF_X1 output4 (.A(net4),
    .Z(count[2]));
 BUF_X1 output5 (.A(net5),
    .Z(count[3]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X16 FILLER_0_97 ();
 FILLCELL_X1 FILLER_0_113 ();
 FILLCELL_X32 FILLER_0_117 ();
 FILLCELL_X32 FILLER_0_149 ();
 FILLCELL_X32 FILLER_0_181 ();
 FILLCELL_X16 FILLER_0_213 ();
 FILLCELL_X8 FILLER_0_229 ();
 FILLCELL_X1 FILLER_0_237 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X16 FILLER_1_97 ();
 FILLCELL_X4 FILLER_1_113 ();
 FILLCELL_X2 FILLER_1_117 ();
 FILLCELL_X1 FILLER_1_119 ();
 FILLCELL_X32 FILLER_1_123 ();
 FILLCELL_X32 FILLER_1_155 ();
 FILLCELL_X32 FILLER_1_187 ();
 FILLCELL_X16 FILLER_1_219 ();
 FILLCELL_X2 FILLER_1_235 ();
 FILLCELL_X1 FILLER_1_237 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X8 FILLER_2_225 ();
 FILLCELL_X4 FILLER_2_233 ();
 FILLCELL_X1 FILLER_2_237 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X8 FILLER_3_225 ();
 FILLCELL_X4 FILLER_3_233 ();
 FILLCELL_X1 FILLER_3_237 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X8 FILLER_4_225 ();
 FILLCELL_X4 FILLER_4_233 ();
 FILLCELL_X1 FILLER_4_237 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X8 FILLER_5_225 ();
 FILLCELL_X4 FILLER_5_233 ();
 FILLCELL_X1 FILLER_5_237 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X8 FILLER_6_225 ();
 FILLCELL_X4 FILLER_6_233 ();
 FILLCELL_X1 FILLER_6_237 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X8 FILLER_7_225 ();
 FILLCELL_X4 FILLER_7_233 ();
 FILLCELL_X1 FILLER_7_237 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X8 FILLER_8_225 ();
 FILLCELL_X4 FILLER_8_233 ();
 FILLCELL_X1 FILLER_8_237 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X8 FILLER_9_225 ();
 FILLCELL_X4 FILLER_9_233 ();
 FILLCELL_X1 FILLER_9_237 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X8 FILLER_10_225 ();
 FILLCELL_X4 FILLER_10_233 ();
 FILLCELL_X1 FILLER_10_237 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X8 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_142 ();
 FILLCELL_X32 FILLER_11_174 ();
 FILLCELL_X32 FILLER_11_206 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X8 FILLER_12_225 ();
 FILLCELL_X4 FILLER_12_233 ();
 FILLCELL_X1 FILLER_12_237 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X16 FILLER_13_97 ();
 FILLCELL_X2 FILLER_13_113 ();
 FILLCELL_X1 FILLER_13_115 ();
 FILLCELL_X8 FILLER_13_133 ();
 FILLCELL_X32 FILLER_13_158 ();
 FILLCELL_X4 FILLER_13_190 ();
 FILLCELL_X2 FILLER_13_194 ();
 FILLCELL_X1 FILLER_13_196 ();
 FILLCELL_X32 FILLER_13_204 ();
 FILLCELL_X2 FILLER_13_236 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X16 FILLER_14_97 ();
 FILLCELL_X8 FILLER_14_113 ();
 FILLCELL_X2 FILLER_14_121 ();
 FILLCELL_X4 FILLER_14_127 ();
 FILLCELL_X2 FILLER_14_131 ();
 FILLCELL_X1 FILLER_14_133 ();
 FILLCELL_X4 FILLER_14_141 ();
 FILLCELL_X2 FILLER_14_145 ();
 FILLCELL_X32 FILLER_14_158 ();
 FILLCELL_X8 FILLER_14_190 ();
 FILLCELL_X4 FILLER_14_198 ();
 FILLCELL_X2 FILLER_14_202 ();
 FILLCELL_X1 FILLER_14_204 ();
 FILLCELL_X16 FILLER_14_208 ();
 FILLCELL_X8 FILLER_14_224 ();
 FILLCELL_X4 FILLER_14_232 ();
 FILLCELL_X2 FILLER_14_236 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X16 FILLER_15_97 ();
 FILLCELL_X8 FILLER_15_113 ();
 FILLCELL_X4 FILLER_15_121 ();
 FILLCELL_X1 FILLER_15_125 ();
 FILLCELL_X8 FILLER_15_130 ();
 FILLCELL_X4 FILLER_15_140 ();
 FILLCELL_X1 FILLER_15_148 ();
 FILLCELL_X2 FILLER_15_151 ();
 FILLCELL_X1 FILLER_15_153 ();
 FILLCELL_X32 FILLER_15_159 ();
 FILLCELL_X32 FILLER_15_191 ();
 FILLCELL_X8 FILLER_15_223 ();
 FILLCELL_X4 FILLER_15_231 ();
 FILLCELL_X2 FILLER_15_235 ();
 FILLCELL_X1 FILLER_15_237 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X8 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_144 ();
 FILLCELL_X32 FILLER_16_176 ();
 FILLCELL_X16 FILLER_16_208 ();
 FILLCELL_X8 FILLER_16_224 ();
 FILLCELL_X4 FILLER_16_232 ();
 FILLCELL_X2 FILLER_16_236 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X16 FILLER_17_97 ();
 FILLCELL_X8 FILLER_17_113 ();
 FILLCELL_X2 FILLER_17_121 ();
 FILLCELL_X4 FILLER_17_131 ();
 FILLCELL_X4 FILLER_17_142 ();
 FILLCELL_X1 FILLER_17_146 ();
 FILLCELL_X1 FILLER_17_157 ();
 FILLCELL_X2 FILLER_17_162 ();
 FILLCELL_X32 FILLER_17_171 ();
 FILLCELL_X32 FILLER_17_203 ();
 FILLCELL_X2 FILLER_17_235 ();
 FILLCELL_X1 FILLER_17_237 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X16 FILLER_18_97 ();
 FILLCELL_X4 FILLER_18_113 ();
 FILLCELL_X2 FILLER_18_117 ();
 FILLCELL_X1 FILLER_18_119 ();
 FILLCELL_X32 FILLER_18_154 ();
 FILLCELL_X32 FILLER_18_186 ();
 FILLCELL_X16 FILLER_18_218 ();
 FILLCELL_X4 FILLER_18_234 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X8 FILLER_19_225 ();
 FILLCELL_X4 FILLER_19_233 ();
 FILLCELL_X1 FILLER_19_237 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X8 FILLER_20_225 ();
 FILLCELL_X4 FILLER_20_233 ();
 FILLCELL_X1 FILLER_20_237 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X8 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_142 ();
 FILLCELL_X32 FILLER_21_174 ();
 FILLCELL_X32 FILLER_21_206 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X8 FILLER_22_225 ();
 FILLCELL_X4 FILLER_22_233 ();
 FILLCELL_X1 FILLER_22_237 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X8 FILLER_23_225 ();
 FILLCELL_X4 FILLER_23_233 ();
 FILLCELL_X1 FILLER_23_237 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X8 FILLER_24_225 ();
 FILLCELL_X4 FILLER_24_233 ();
 FILLCELL_X1 FILLER_24_237 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X8 FILLER_25_225 ();
 FILLCELL_X4 FILLER_25_233 ();
 FILLCELL_X1 FILLER_25_237 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X8 FILLER_26_225 ();
 FILLCELL_X4 FILLER_26_233 ();
 FILLCELL_X1 FILLER_26_237 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X8 FILLER_27_225 ();
 FILLCELL_X4 FILLER_27_233 ();
 FILLCELL_X1 FILLER_27_237 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X8 FILLER_28_225 ();
 FILLCELL_X4 FILLER_28_233 ();
 FILLCELL_X1 FILLER_28_237 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X8 FILLER_29_225 ();
 FILLCELL_X4 FILLER_29_233 ();
 FILLCELL_X1 FILLER_29_237 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X8 FILLER_30_225 ();
 FILLCELL_X4 FILLER_30_233 ();
 FILLCELL_X1 FILLER_30_237 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X16 FILLER_31_97 ();
 FILLCELL_X8 FILLER_31_113 ();
 FILLCELL_X4 FILLER_31_121 ();
 FILLCELL_X2 FILLER_31_125 ();
 FILLCELL_X1 FILLER_31_127 ();
 FILLCELL_X8 FILLER_31_131 ();
 FILLCELL_X32 FILLER_31_142 ();
 FILLCELL_X32 FILLER_31_174 ();
 FILLCELL_X32 FILLER_31_206 ();
endmodule
