module configurable_kogge_stone_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _327_ (.I(net1),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _328_ (.I(net33),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _329_ (.I(net65),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _330_ (.I(_004_),
    .ZN(net67));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _331_ (.I(_005_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _332_ (.A1(_014_),
    .A2(_016_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _333_ (.A1(_010_),
    .A2(_012_),
    .A3(_070_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _334_ (.A1(_066_),
    .A2(_067_),
    .A3(_064_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _335_ (.A1(_064_),
    .A2(_065_),
    .B(_063_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _336_ (.A1(_062_),
    .A2(_060_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _337_ (.A1(_056_),
    .A2(_058_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _338_ (.A1(_072_),
    .A2(_073_),
    .B(_074_),
    .C(_075_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _339_ (.A1(_060_),
    .A2(_061_),
    .B(_059_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _340_ (.A1(_056_),
    .A2(_057_),
    .B(_055_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _341_ (.A1(_075_),
    .A2(_077_),
    .B(_078_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _342_ (.I(_050_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _343_ (.I(_049_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _344_ (.I(_048_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _345_ (.A1(_080_),
    .A2(_081_),
    .B(_082_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _346_ (.A1(_052_),
    .A2(_054_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _347_ (.A1(_076_),
    .A2(_079_),
    .B1(_083_),
    .B2(_047_),
    .C(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _348_ (.A1(_052_),
    .A2(_053_),
    .B(_051_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _349_ (.A1(_048_),
    .A2(_049_),
    .B(_047_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _350_ (.A1(_082_),
    .A2(_080_),
    .A3(_086_),
    .B(_087_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _351_ (.A1(_028_),
    .A2(_029_),
    .B(_027_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _352_ (.A1(_043_),
    .A2(_045_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _353_ (.A1(_040_),
    .A2(_041_),
    .B(_039_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _354_ (.A1(_089_),
    .A2(_090_),
    .A3(_091_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _355_ (.A1(_032_),
    .A2(_034_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _356_ (.A1(_036_),
    .A2(_037_),
    .B(_035_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _357_ (.A1(_032_),
    .A2(_033_),
    .B(_031_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _358_ (.A1(_093_),
    .A2(_094_),
    .B(_095_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _359_ (.A1(_088_),
    .A2(_092_),
    .A3(_096_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _360_ (.A1(_085_),
    .A2(_097_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _361_ (.A1(_028_),
    .A2(_030_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _362_ (.A1(_046_),
    .A2(_043_),
    .A3(_045_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _363_ (.A1(_028_),
    .A2(_030_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _364_ (.A1(_091_),
    .A2(_100_),
    .B(_101_),
    .C(_093_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _365_ (.A1(_044_),
    .A2(_043_),
    .B(_040_),
    .C(_042_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _366_ (.A1(_036_),
    .A2(_038_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _367_ (.A1(_091_),
    .A2(_103_),
    .B(_104_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _368_ (.I(_089_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _369_ (.A1(_096_),
    .A2(_099_),
    .B1(_102_),
    .B2(_105_),
    .C(_106_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _370_ (.A1(_098_),
    .A2(_107_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _371_ (.A1(_024_),
    .A2(_026_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _372_ (.A1(_018_),
    .A2(_020_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _373_ (.A1(_022_),
    .A2(_109_),
    .A3(_110_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _374_ (.A1(_024_),
    .A2(_025_),
    .B(_023_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _375_ (.I(_112_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _376_ (.A1(_022_),
    .A2(_113_),
    .B(_021_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _377_ (.A1(_018_),
    .A2(_020_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _378_ (.A1(_018_),
    .A2(_019_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _379_ (.A1(_017_),
    .A2(_116_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _380_ (.I(_117_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _381_ (.A1(_108_),
    .A2(_111_),
    .B1(_114_),
    .B2(_115_),
    .C(_118_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _382_ (.A1(_012_),
    .A2(_013_),
    .B(_011_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _383_ (.I(_120_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _384_ (.A1(_010_),
    .A2(_121_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _385_ (.A1(_010_),
    .A2(_012_),
    .A3(_014_),
    .A4(_015_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _386_ (.A1(_009_),
    .A2(_122_),
    .A3(_123_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _387_ (.A1(_071_),
    .A2(_119_),
    .B(_124_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _388_ (.A1(_066_),
    .A2(_064_),
    .A3(_068_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _389_ (.A1(_062_),
    .A2(_060_),
    .A3(_126_),
    .Z(_127_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _390_ (.I(_003_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _391_ (.A1(_061_),
    .A2(_063_),
    .Z(_129_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _392_ (.A1(_067_),
    .A2(_128_),
    .A3(_065_),
    .A4(_129_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _393_ (.A1(_066_),
    .A2(_067_),
    .B(_065_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _394_ (.A1(_062_),
    .A2(_060_),
    .A3(_064_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _395_ (.A1(_062_),
    .A2(_060_),
    .A3(_063_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _396_ (.A1(_131_),
    .A2(_132_),
    .B(_133_),
    .C(_077_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _397_ (.A1(_127_),
    .A2(_130_),
    .B(_134_),
    .C(_057_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _398_ (.A1(_062_),
    .A2(_056_),
    .A3(_058_),
    .A4(_060_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _399_ (.A1(_136_),
    .A2(_126_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _400_ (.A1(_050_),
    .A2(_052_),
    .A3(_054_),
    .Z(_138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _401_ (.A1(_137_),
    .A2(_138_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _402_ (.A1(_080_),
    .A2(_086_),
    .B(_081_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _403_ (.A1(_045_),
    .A2(_047_),
    .A3(_140_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _404_ (.A1(_076_),
    .A2(_079_),
    .B(_138_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _405_ (.A1(_135_),
    .A2(_139_),
    .B(_141_),
    .C(_142_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _406_ (.A1(_044_),
    .A2(_043_),
    .Z(_144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _407_ (.A1(_042_),
    .A2(_144_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _408_ (.I(_046_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _409_ (.A1(_146_),
    .A2(_087_),
    .B(_090_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _410_ (.I(_057_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _411_ (.A1(_054_),
    .A2(_055_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _412_ (.A1(_051_),
    .A2(_053_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _413_ (.A1(_148_),
    .A2(_149_),
    .A3(_150_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _414_ (.A1(_058_),
    .A2(_134_),
    .B(_147_),
    .C(_151_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _415_ (.A1(_056_),
    .A2(_055_),
    .B(_054_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _416_ (.A1(_052_),
    .A2(_051_),
    .B(_048_),
    .C(_050_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _417_ (.A1(_150_),
    .A2(_153_),
    .B(_154_),
    .C(_146_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _418_ (.A1(_147_),
    .A2(_155_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _419_ (.A1(_145_),
    .A2(_152_),
    .A3(_156_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _420_ (.A1(_041_),
    .A2(_043_),
    .Z(_158_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _421_ (.A1(_036_),
    .A2(_038_),
    .A3(_040_),
    .A4(_042_),
    .Z(_159_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _422_ (.A1(_044_),
    .A2(_046_),
    .Z(_160_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _423_ (.A1(_048_),
    .A2(_050_),
    .A3(_052_),
    .A4(_054_),
    .Z(_161_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _424_ (.A1(_136_),
    .A2(_126_),
    .A3(_160_),
    .A4(_161_),
    .Z(_162_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _425_ (.A1(_159_),
    .A2(_162_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _426_ (.A1(_143_),
    .A2(_157_),
    .A3(_158_),
    .B(_163_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _427_ (.A1(_036_),
    .A2(_037_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _428_ (.A1(_091_),
    .A2(_104_),
    .B(_165_),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _429_ (.A1(_035_),
    .A2(_166_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _430_ (.A1(_048_),
    .A2(_045_),
    .A3(_047_),
    .Z(_168_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _431_ (.A1(_046_),
    .A2(_045_),
    .Z(_169_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _432_ (.A1(_044_),
    .A2(_168_),
    .A3(_169_),
    .Z(_170_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _433_ (.A1(_159_),
    .A2(_138_),
    .Z(_171_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _434_ (.A1(_076_),
    .A2(_079_),
    .B(_170_),
    .C(_171_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _435_ (.A1(_045_),
    .A2(_047_),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _436_ (.A1(_080_),
    .A2(_086_),
    .B(_173_),
    .C(_081_),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _437_ (.A1(_044_),
    .A2(_159_),
    .A3(_168_),
    .A4(_169_),
    .Z(_175_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _438_ (.A1(_043_),
    .A2(_159_),
    .B1(_174_),
    .B2(_175_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _439_ (.A1(_167_),
    .A2(_172_),
    .A3(_176_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _440_ (.A1(_030_),
    .A2(_032_),
    .Z(_178_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _441_ (.A1(_026_),
    .A2(_028_),
    .A3(_178_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _442_ (.A1(_034_),
    .A2(_035_),
    .Z(_180_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _443_ (.A1(_034_),
    .A2(_166_),
    .B(_180_),
    .C(_033_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _444_ (.I(_028_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _445_ (.A1(_030_),
    .A2(_031_),
    .B(_029_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _446_ (.I(_027_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _447_ (.A1(_182_),
    .A2(_183_),
    .B(_184_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _448_ (.A1(_026_),
    .A2(_185_),
    .B(_025_),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _449_ (.I(_019_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _450_ (.A1(_187_),
    .A2(_089_),
    .Z(_188_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _451_ (.A1(_179_),
    .A2(_181_),
    .B(_186_),
    .C(_188_),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _452_ (.A1(_034_),
    .A2(_036_),
    .A3(_038_),
    .A4(_040_),
    .Z(_190_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _453_ (.A1(_042_),
    .A2(_144_),
    .A3(_190_),
    .Z(_191_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _454_ (.A1(_147_),
    .A2(_155_),
    .B(_191_),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _455_ (.A1(_152_),
    .A2(_192_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _456_ (.I(_096_),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _457_ (.A1(_194_),
    .A2(_183_),
    .A3(_181_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _458_ (.A1(_177_),
    .A2(_189_),
    .A3(_193_),
    .A4(_195_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _459_ (.A1(_022_),
    .A2(_024_),
    .A3(_110_),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _460_ (.A1(_179_),
    .A2(_197_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _461_ (.A1(_042_),
    .A2(_190_),
    .A3(_162_),
    .Z(_199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _462_ (.A1(_198_),
    .A2(_199_),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _463_ (.A1(_164_),
    .A2(_196_),
    .B(_200_),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _464_ (.A1(_071_),
    .A2(_190_),
    .Z(_202_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _465_ (.A1(_093_),
    .A2(_101_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _466_ (.A1(_022_),
    .A2(_024_),
    .A3(_026_),
    .Z(_204_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _467_ (.A1(_020_),
    .A2(_204_),
    .Z(_205_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _468_ (.A1(_012_),
    .A2(_018_),
    .A3(_070_),
    .Z(_206_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _469_ (.A1(_203_),
    .A2(_159_),
    .A3(_205_),
    .A4(_206_),
    .Z(_207_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _470_ (.A1(_202_),
    .A2(_162_),
    .A3(_198_),
    .A4(_207_),
    .Z(_208_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _471_ (.A1(_119_),
    .A2(_201_),
    .B(_208_),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _472_ (.I(_008_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _473_ (.A1(_125_),
    .A2(_209_),
    .B(_210_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _474_ (.A1(_007_),
    .A2(_211_),
    .B(_006_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _475_ (.A1(_069_),
    .A2(_212_),
    .ZN(net66));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _476_ (.I(_138_),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _477_ (.A1(_127_),
    .A2(_130_),
    .B(_134_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _478_ (.A1(_148_),
    .A2(_214_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _479_ (.A1(_137_),
    .A2(_215_),
    .B(_076_),
    .C(_079_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _480_ (.A1(_213_),
    .A2(_216_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _481_ (.A1(_140_),
    .A2(_217_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _482_ (.A1(_048_),
    .A2(_218_),
    .ZN(net68));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _483_ (.A1(_048_),
    .A2(_140_),
    .B(_047_),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _484_ (.A1(_085_),
    .A2(_219_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _485_ (.A1(_137_),
    .A2(_161_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _486_ (.A1(_221_),
    .A2(_218_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _487_ (.A1(_220_),
    .A2(_222_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _488_ (.A1(_046_),
    .A2(_223_),
    .ZN(net69));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _489_ (.A1(_135_),
    .A2(_139_),
    .Z(_224_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _490_ (.A1(_141_),
    .A2(_142_),
    .A3(_224_),
    .Z(_225_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _491_ (.A1(_085_),
    .A2(_219_),
    .A3(_221_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _492_ (.A1(_046_),
    .A2(_226_),
    .B(_045_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _493_ (.A1(_225_),
    .A2(_227_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _494_ (.A1(_044_),
    .A2(_228_),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _495_ (.A1(_044_),
    .A2(_168_),
    .A3(_169_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _496_ (.A1(_141_),
    .A2(_142_),
    .B(_229_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _497_ (.A1(_043_),
    .A2(_230_),
    .Z(_231_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _498_ (.A1(_162_),
    .A2(_228_),
    .B(_231_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _499_ (.A1(_042_),
    .A2(_232_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _500_ (.A1(_042_),
    .A2(_162_),
    .Z(_233_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _501_ (.A1(_043_),
    .A2(_230_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _502_ (.A1(_225_),
    .A2(_227_),
    .B(_234_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _503_ (.A1(_233_),
    .A2(_235_),
    .B(_041_),
    .C(_157_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _504_ (.A1(_040_),
    .A2(_236_),
    .ZN(net72));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _505_ (.I(_040_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _506_ (.I(_039_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _507_ (.A1(_237_),
    .A2(_236_),
    .B(_238_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _508_ (.A1(_038_),
    .A2(_239_),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _509_ (.A1(_038_),
    .A2(_239_),
    .B(_037_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _510_ (.A1(_036_),
    .A2(_240_),
    .ZN(net74));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _511_ (.A1(_164_),
    .A2(_167_),
    .A3(_172_),
    .A4(_176_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _512_ (.A1(_034_),
    .A2(_241_),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _513_ (.I(_181_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _514_ (.A1(_242_),
    .A2(_193_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _515_ (.A1(_241_),
    .A2(_199_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _516_ (.A1(_243_),
    .A2(_244_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _517_ (.A1(_032_),
    .A2(_245_),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _518_ (.A1(_032_),
    .A2(_034_),
    .A3(_163_),
    .Z(_246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _519_ (.A1(_046_),
    .A2(_220_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _520_ (.A1(_090_),
    .A2(_091_),
    .A3(_247_),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _521_ (.A1(_032_),
    .A2(_034_),
    .A3(_105_),
    .A4(_248_),
    .Z(_249_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _522_ (.A1(_245_),
    .A2(_246_),
    .B(_249_),
    .C(_096_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _523_ (.A1(_030_),
    .A2(_250_),
    .ZN(net77));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _524_ (.A1(_066_),
    .A2(_003_),
    .ZN(net78));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _525_ (.A1(_177_),
    .A2(_193_),
    .A3(_195_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _526_ (.A1(_190_),
    .A2(_233_),
    .Z(_252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _527_ (.A1(_178_),
    .A2(_252_),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _528_ (.I(_178_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _529_ (.A1(_254_),
    .A2(_181_),
    .Z(_255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _530_ (.A1(_178_),
    .A2(_191_),
    .ZN(_256_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _531_ (.A1(_152_),
    .A2(_156_),
    .A3(_256_),
    .Z(_257_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _532_ (.A1(_183_),
    .A2(_255_),
    .A3(_257_),
    .Z(_258_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _533_ (.A1(_164_),
    .A2(_251_),
    .B1(_253_),
    .B2(_258_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _534_ (.A1(_182_),
    .A2(_259_),
    .ZN(net79));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _535_ (.A1(_203_),
    .A2(_163_),
    .Z(_260_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _536_ (.A1(_085_),
    .A2(_097_),
    .B(_107_),
    .ZN(_261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _537_ (.A1(_260_),
    .A2(_259_),
    .B(_261_),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _538_ (.A1(_026_),
    .A2(_262_),
    .ZN(net80));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _539_ (.I(_186_),
    .ZN(_263_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _540_ (.A1(_261_),
    .A2(_260_),
    .B(_199_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _541_ (.A1(_243_),
    .A2(_264_),
    .B(_179_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _542_ (.A1(_106_),
    .A2(_263_),
    .A3(_242_),
    .Z(_266_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _543_ (.A1(_263_),
    .A2(_265_),
    .B1(_266_),
    .B2(_259_),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _544_ (.A1(_024_),
    .A2(_267_),
    .ZN(net81));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _545_ (.A1(_263_),
    .A2(_265_),
    .B1(_266_),
    .B2(_259_),
    .C(_260_),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _546_ (.A1(_108_),
    .A2(_268_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _547_ (.A1(_109_),
    .A2(_269_),
    .B(_113_),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _548_ (.A1(_022_),
    .A2(_270_),
    .ZN(net82));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _549_ (.A1(_261_),
    .A2(_204_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _550_ (.A1(_114_),
    .A2(_271_),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _551_ (.A1(_022_),
    .A2(_024_),
    .A3(_026_),
    .A4(_028_),
    .Z(_273_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _552_ (.A1(_178_),
    .A2(_252_),
    .A3(_273_),
    .Z(_274_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _553_ (.A1(_108_),
    .A2(_112_),
    .A3(_114_),
    .A4(_268_),
    .ZN(_275_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _554_ (.A1(_272_),
    .A2(_274_),
    .B(_275_),
    .ZN(_276_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _555_ (.A1(_020_),
    .A2(_276_),
    .ZN(net83));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _556_ (.A1(_205_),
    .A2(_260_),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _557_ (.A1(_164_),
    .A2(_196_),
    .B1(_277_),
    .B2(_187_),
    .ZN(_278_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _558_ (.A1(_020_),
    .A2(_272_),
    .B(_278_),
    .ZN(_279_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _559_ (.A1(_018_),
    .A2(_279_),
    .ZN(net84));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _560_ (.I(_016_),
    .ZN(_280_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _561_ (.A1(_119_),
    .A2(_201_),
    .ZN(_281_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _562_ (.A1(_016_),
    .A2(_204_),
    .A3(_260_),
    .Z(_282_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _563_ (.A1(_117_),
    .A2(_272_),
    .A3(_282_),
    .ZN(_283_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _564_ (.A1(_110_),
    .A2(_117_),
    .B(_016_),
    .ZN(_284_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _565_ (.A1(_281_),
    .A2(_283_),
    .A3(_284_),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _566_ (.A1(_280_),
    .A2(_281_),
    .B(_285_),
    .ZN(net85));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _567_ (.A1(_015_),
    .A2(_285_),
    .ZN(_286_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _568_ (.A1(_014_),
    .A2(_286_),
    .ZN(net86));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _569_ (.A1(_070_),
    .A2(_110_),
    .Z(_287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _570_ (.A1(_274_),
    .A2(_287_),
    .ZN(_288_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _571_ (.A1(_015_),
    .A2(_274_),
    .A3(_287_),
    .Z(_289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _572_ (.A1(_272_),
    .A2(_287_),
    .B(_289_),
    .ZN(_290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _573_ (.A1(_016_),
    .A2(_117_),
    .Z(_291_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _574_ (.A1(_015_),
    .A2(_291_),
    .Z(_292_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _575_ (.A1(_014_),
    .A2(_292_),
    .B(_013_),
    .ZN(_293_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _576_ (.A1(_281_),
    .A2(_288_),
    .B(_290_),
    .C(_293_),
    .ZN(_294_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _577_ (.A1(_012_),
    .A2(_294_),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _578_ (.I(_020_),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _579_ (.I(_205_),
    .ZN(_296_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _580_ (.I(_035_),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _581_ (.A1(_091_),
    .A2(_104_),
    .B(_165_),
    .C(_297_),
    .ZN(_298_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _582_ (.I(_030_),
    .ZN(_299_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _583_ (.I(_029_),
    .ZN(_300_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _584_ (.A1(_299_),
    .A2(_095_),
    .B(_300_),
    .ZN(_301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _585_ (.A1(_203_),
    .A2(_298_),
    .B1(_301_),
    .B2(_028_),
    .C(_027_),
    .ZN(_302_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _586_ (.A1(_295_),
    .A2(_114_),
    .B1(_296_),
    .B2(_302_),
    .C(_187_),
    .ZN(_303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _587_ (.A1(_016_),
    .A2(_018_),
    .Z(_304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _588_ (.A1(_016_),
    .A2(_017_),
    .B1(_303_),
    .B2(_304_),
    .C(_015_),
    .ZN(_305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _589_ (.A1(_012_),
    .A2(_014_),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _590_ (.A1(_305_),
    .A2(_306_),
    .B(_120_),
    .ZN(_307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _591_ (.A1(_234_),
    .A2(_293_),
    .ZN(_308_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _592_ (.A1(_307_),
    .A2(_308_),
    .ZN(_309_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _593_ (.A1(_281_),
    .A2(_288_),
    .B(_290_),
    .C(_309_),
    .ZN(_310_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _594_ (.A1(_162_),
    .A2(_231_),
    .A3(_307_),
    .Z(_311_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _595_ (.A1(_207_),
    .A2(_307_),
    .B(_310_),
    .C(_311_),
    .ZN(_312_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _596_ (.A1(_010_),
    .A2(_312_),
    .ZN(net88));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _597_ (.A1(_128_),
    .A2(_068_),
    .Z(_313_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _598_ (.A1(_067_),
    .A2(_313_),
    .Z(_314_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _599_ (.A1(_066_),
    .A2(_314_),
    .B(_065_),
    .ZN(_315_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _600_ (.A1(_064_),
    .A2(_315_),
    .ZN(net89));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _601_ (.A1(_210_),
    .A2(_125_),
    .A3(_209_),
    .Z(_316_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _602_ (.A1(_211_),
    .A2(_316_),
    .ZN(net90));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _603_ (.A1(_006_),
    .A2(_007_),
    .A3(_211_),
    .Z(_317_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _604_ (.A1(_212_),
    .A2(_317_),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _605_ (.A1(_067_),
    .A2(_128_),
    .A3(_065_),
    .B(_126_),
    .ZN(_318_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _606_ (.A1(_072_),
    .A2(_073_),
    .A3(_318_),
    .ZN(_319_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _607_ (.A1(_062_),
    .A2(_319_),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _608_ (.A1(_062_),
    .A2(_319_),
    .B(_061_),
    .ZN(_320_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _609_ (.A1(_060_),
    .A2(_320_),
    .ZN(net93));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _610_ (.A1(_058_),
    .A2(_214_),
    .ZN(net94));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _611_ (.I(_214_),
    .ZN(_321_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _612_ (.A1(_058_),
    .A2(_321_),
    .B(_057_),
    .ZN(_322_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _613_ (.A1(_056_),
    .A2(_322_),
    .ZN(net95));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _614_ (.A1(_054_),
    .A2(_216_),
    .ZN(net96));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _615_ (.I(_054_),
    .ZN(_323_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _616_ (.I(_053_),
    .ZN(_324_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _617_ (.A1(_323_),
    .A2(_216_),
    .B(_324_),
    .ZN(_325_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _618_ (.A1(_052_),
    .A2(_325_),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _619_ (.A1(_052_),
    .A2(_325_),
    .B(_051_),
    .ZN(_326_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _620_ (.A1(_050_),
    .A2(_326_),
    .ZN(net98));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _621_ (.A(_000_),
    .B(_001_),
    .CI(_002_),
    .CO(_003_),
    .S(_004_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _622_ (.A(net25),
    .B(net57),
    .CO(_005_),
    .S(_006_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _623_ (.A(net24),
    .B(net56),
    .CO(_007_),
    .S(_008_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _624_ (.A(net22),
    .B(net54),
    .CO(_009_),
    .S(_010_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _625_ (.A(net21),
    .B(net53),
    .CO(_011_),
    .S(_012_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _626_ (.A(net20),
    .B(net52),
    .CO(_013_),
    .S(_014_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _627_ (.A(net19),
    .B(net51),
    .CO(_015_),
    .S(_016_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _628_ (.A(net18),
    .B(net50),
    .CO(_017_),
    .S(_018_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _629_ (.A(net17),
    .B(net49),
    .CO(_019_),
    .S(_020_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _630_ (.A(net16),
    .B(net48),
    .CO(_021_),
    .S(_022_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _631_ (.A(net15),
    .B(net47),
    .CO(_023_),
    .S(_024_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _632_ (.A(net14),
    .B(net46),
    .CO(_025_),
    .S(_026_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _633_ (.A(net13),
    .B(net45),
    .CO(_027_),
    .S(_028_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _634_ (.A(net11),
    .B(net43),
    .CO(_029_),
    .S(_030_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _635_ (.A(net10),
    .B(net42),
    .CO(_031_),
    .S(_032_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _636_ (.A(net9),
    .B(net41),
    .CO(_033_),
    .S(_034_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _637_ (.A(net8),
    .B(net40),
    .CO(_035_),
    .S(_036_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _638_ (.A(net7),
    .B(net39),
    .CO(_037_),
    .S(_038_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _639_ (.A(net6),
    .B(net38),
    .CO(_039_),
    .S(_040_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _640_ (.A(net5),
    .B(net37),
    .CO(_041_),
    .S(_042_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _641_ (.A(net4),
    .B(net36),
    .CO(_043_),
    .S(_044_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _642_ (.A(net3),
    .B(net35),
    .CO(_045_),
    .S(_046_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _643_ (.A(net2),
    .B(net34),
    .CO(_047_),
    .S(_048_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _644_ (.A(net32),
    .B(net64),
    .CO(_049_),
    .S(_050_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _645_ (.A(net31),
    .B(net63),
    .CO(_051_),
    .S(_052_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _646_ (.A(net30),
    .B(net62),
    .CO(_053_),
    .S(_054_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _647_ (.A(net29),
    .B(net61),
    .CO(_055_),
    .S(_056_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _648_ (.A(net28),
    .B(net60),
    .CO(_057_),
    .S(_058_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _649_ (.A(net27),
    .B(net59),
    .CO(_059_),
    .S(_060_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _650_ (.A(net26),
    .B(net58),
    .CO(_061_),
    .S(_062_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _651_ (.A(net23),
    .B(net55),
    .CO(_063_),
    .S(_064_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _652_ (.A(net12),
    .B(net44),
    .CO(_065_),
    .S(_066_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _653_ (.A(net1),
    .B(net33),
    .CO(_067_),
    .S(_068_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(a[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(a[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(a[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(a[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(a[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(a[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(a[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(a[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(a[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(a[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(a[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(a[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(a[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(a[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(a[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(a[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(a[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(a[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(a[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(a[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(a[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(a[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(a[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(a[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(a[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(a[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(a[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(a[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(a[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(a[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(a[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(a[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input33 (.I(b[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(b[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(b[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(b[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(b[13]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(b[14]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input39 (.I(b[15]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input40 (.I(b[16]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(b[17]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(b[18]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(b[19]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input44 (.I(b[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(b[20]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input46 (.I(b[21]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input47 (.I(b[22]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(b[23]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(b[24]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input50 (.I(b[25]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input51 (.I(b[26]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(b[27]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(b[28]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input54 (.I(b[29]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input55 (.I(b[2]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input56 (.I(b[30]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input57 (.I(b[31]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input58 (.I(b[3]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input59 (.I(b[4]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input60 (.I(b[5]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input61 (.I(b[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input62 (.I(b[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input63 (.I(b[8]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input64 (.I(b[9]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input65 (.I(cin),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net66),
    .Z(cout));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net67),
    .Z(sum[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net68),
    .Z(sum[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net69),
    .Z(sum[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net70),
    .Z(sum[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net71),
    .Z(sum[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net72),
    .Z(sum[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net73),
    .Z(sum[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net74),
    .Z(sum[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net75),
    .Z(sum[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net76),
    .Z(sum[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net77),
    .Z(sum[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net78),
    .Z(sum[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net79),
    .Z(sum[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net80),
    .Z(sum[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net81),
    .Z(sum[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net82),
    .Z(sum[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net83),
    .Z(sum[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output84 (.I(net84),
    .Z(sum[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output85 (.I(net85),
    .Z(sum[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output86 (.I(net86),
    .Z(sum[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output87 (.I(net87),
    .Z(sum[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output88 (.I(net88),
    .Z(sum[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net89),
    .Z(sum[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output90 (.I(net90),
    .Z(sum[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output91 (.I(net91),
    .Z(sum[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net92),
    .Z(sum[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net93),
    .Z(sum[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net94),
    .Z(sum[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net95),
    .Z(sum[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net96),
    .Z(sum[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net97),
    .Z(sum[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net98),
    .Z(sum[9]));
endmodule
