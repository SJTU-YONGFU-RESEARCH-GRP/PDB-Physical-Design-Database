module hamming_code (single_bit_error,
    corrected_code,
    data_in,
    data_out,
    encoded_out,
    received_in);
 output single_bit_error;
 output [6:0] corrected_code;
 input [3:0] data_in;
 output [3:0] data_out;
 output [6:0] encoded_out;
 input [6:0] received_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire p1;
 wire p2;
 wire p3;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;

 gf180mcu_fd_sc_mcu9t5v0__buf_4 _075_ (.I(net10),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _076_ (.A1(_004_),
    .A2(net8),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _077_ (.I(net11),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _078_ (.A1(net9),
    .A2(_006_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _079_ (.A1(_005_),
    .A2(_007_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _080_ (.A1(_005_),
    .A2(_007_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _081_ (.A1(net7),
    .A2(net5),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _082_ (.I(_010_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _083_ (.I0(_008_),
    .I1(_009_),
    .S(_011_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _084_ (.A1(net7),
    .A2(net6),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _085_ (.A1(net11),
    .A2(net10),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _086_ (.A1(_013_),
    .A2(_014_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _087_ (.A1(_012_),
    .A2(_015_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _088_ (.A1(net5),
    .A2(_016_),
    .ZN(net12));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _089_ (.A1(net7),
    .A2(_014_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _090_ (.A1(net7),
    .A2(net5),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _091_ (.I(_018_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _092_ (.I0(_008_),
    .I1(_009_),
    .S(_019_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _093_ (.I0(net6),
    .I1(_017_),
    .S(_020_),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _094_ (.A1(net6),
    .A2(_014_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _095_ (.I0(net7),
    .I1(_021_),
    .S(_012_),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _096_ (.I(net8),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _097_ (.I(_013_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _098_ (.A1(_019_),
    .A2(_023_),
    .B(_022_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _099_ (.A1(_022_),
    .A2(_011_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _100_ (.A1(_004_),
    .A2(_024_),
    .B(_025_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _101_ (.I(_006_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _102_ (.A1(net7),
    .A2(net6),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _103_ (.I(net8),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _104_ (.A1(_019_),
    .A2(_028_),
    .B(_029_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _105_ (.I(_004_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _106_ (.A1(_031_),
    .A2(_011_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _107_ (.A1(_006_),
    .A2(_030_),
    .A3(_032_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _108_ (.A1(_022_),
    .A2(_023_),
    .B1(_026_),
    .B2(_027_),
    .C(_033_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _109_ (.A1(_019_),
    .A2(_028_),
    .B(_022_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _110_ (.A1(_004_),
    .A2(_035_),
    .B(_025_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _111_ (.A1(_019_),
    .A2(_013_),
    .B(_029_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _112_ (.A1(_027_),
    .A2(_032_),
    .A3(_037_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _113_ (.A1(_022_),
    .A2(_028_),
    .B1(_036_),
    .B2(_006_),
    .C(_038_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _114_ (.I0(_034_),
    .I1(_039_),
    .S(net9),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _115_ (.A1(_029_),
    .A2(_013_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _116_ (.I(net9),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _117_ (.A1(_041_),
    .A2(_031_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _118_ (.A1(_040_),
    .A2(_042_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _119_ (.A1(_031_),
    .A2(_022_),
    .A3(_019_),
    .A4(_023_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _120_ (.A1(_041_),
    .A2(_019_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _121_ (.A1(_029_),
    .A2(_023_),
    .B(_041_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _122_ (.A1(_022_),
    .A2(_011_),
    .A3(_013_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _123_ (.A1(_046_),
    .A2(_047_),
    .B(_031_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _124_ (.A1(_043_),
    .A2(_044_),
    .A3(_045_),
    .A4(_048_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _125_ (.A1(_011_),
    .A2(_023_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _126_ (.A1(_029_),
    .A2(_050_),
    .B1(_040_),
    .B2(net9),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _127_ (.A1(_022_),
    .A2(_018_),
    .A3(_013_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _128_ (.A1(_046_),
    .A2(_052_),
    .B(_004_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _129_ (.A1(_041_),
    .A2(_011_),
    .B1(_051_),
    .B2(_004_),
    .C(_053_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _130_ (.I0(_049_),
    .I1(_054_),
    .S(_006_),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _131_ (.A1(_029_),
    .A2(_019_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _132_ (.A1(net9),
    .A2(_031_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _133_ (.A1(_041_),
    .A2(_029_),
    .A3(_011_),
    .A4(_023_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _134_ (.A1(_004_),
    .A2(_023_),
    .B1(_055_),
    .B2(_056_),
    .C(_057_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _135_ (.A1(_031_),
    .A2(_025_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _136_ (.A1(_052_),
    .A2(_059_),
    .B(net9),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _137_ (.A1(net9),
    .A2(net8),
    .A3(_010_),
    .A4(_028_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _138_ (.A1(_004_),
    .A2(_028_),
    .B1(_055_),
    .B2(_042_),
    .C(_061_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _139_ (.A1(net9),
    .A2(_031_),
    .A3(_025_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _140_ (.A1(net9),
    .A2(_029_),
    .A3(_011_),
    .A4(_023_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _141_ (.A1(_006_),
    .A2(_062_),
    .A3(_063_),
    .A4(_064_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _142_ (.A1(_027_),
    .A2(_058_),
    .A3(_060_),
    .B(_065_),
    .ZN(net17));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _143_ (.A1(_031_),
    .A2(_023_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _144_ (.A1(_031_),
    .A2(_029_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _145_ (.A1(_067_),
    .A2(_019_),
    .B(_006_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _146_ (.A1(_067_),
    .A2(_050_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _147_ (.A1(_019_),
    .A2(_023_),
    .B(_006_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _148_ (.A1(_004_),
    .A2(_022_),
    .A3(_070_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _149_ (.A1(_041_),
    .A2(_068_),
    .A3(_069_),
    .A4(_071_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _150_ (.A1(_011_),
    .A2(_013_),
    .B(_006_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _151_ (.A1(_004_),
    .A2(_029_),
    .A3(_073_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _152_ (.A1(_031_),
    .A2(_022_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _153_ (.A1(_011_),
    .A2(_000_),
    .B(_006_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _154_ (.A1(net9),
    .A2(_044_),
    .A3(_074_),
    .A4(_001_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _155_ (.A1(_027_),
    .A2(_066_),
    .B1(_072_),
    .B2(_002_),
    .ZN(net18));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _156_ (.A1(net4),
    .A2(net2),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _157_ (.A1(net1),
    .A2(_003_),
    .ZN(p1));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _158_ (.A1(net4),
    .A2(net1),
    .A3(net3),
    .Z(p2));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _159_ (.A1(net3),
    .A2(_003_),
    .ZN(p3));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _160_ (.A1(_015_),
    .A2(_020_),
    .ZN(net30));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _161_ (.I(net14),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _162_ (.I(net16),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _163_ (.I(net17),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _164_ (.I(net18),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _165_ (.I(p1),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _166_ (.I(p2),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _167_ (.I(net1),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _168_ (.I(p3),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _169_ (.I(net2),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _170_ (.I(net3),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 _171_ (.I(net4),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_67 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_68 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_69 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_70 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_71 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_72 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_73 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_74 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_75 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_76 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_77 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(data_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(data_in[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(data_in[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(data_in[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(received_in[0]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input6 (.I(received_in[1]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input7 (.I(received_in[2]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input8 (.I(received_in[3]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input9 (.I(received_in[4]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(received_in[5]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(received_in[6]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net12),
    .Z(corrected_code[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net13),
    .Z(corrected_code[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net14),
    .Z(corrected_code[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net15),
    .Z(corrected_code[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net16),
    .Z(corrected_code[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net17),
    .Z(corrected_code[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net18),
    .Z(corrected_code[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net19),
    .Z(data_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net20),
    .Z(data_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net21),
    .Z(data_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net22),
    .Z(data_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net23),
    .Z(encoded_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net24),
    .Z(encoded_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output25 (.I(net25),
    .Z(encoded_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output26 (.I(net26),
    .Z(encoded_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output27 (.I(net27),
    .Z(encoded_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output28 (.I(net28),
    .Z(encoded_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output29 (.I(net29),
    .Z(encoded_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output30 (.I(net30),
    .Z(single_bit_error));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_11 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_290 ();
endmodule
