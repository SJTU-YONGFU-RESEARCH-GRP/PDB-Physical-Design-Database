module parameterized_gray_counter (clk,
    enable,
    rst_n,
    binary_out,
    gray_out);
 input clk;
 input enable;
 input rst_n;
 output [3:0] binary_out;
 output [3:0] gray_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _12_ (.A1(net3),
    .A2(net1),
    .Z(_04_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13_ (.A1(net2),
    .A2(_04_),
    .Z(_00_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14_ (.I0(net4),
    .I1(net7),
    .S(net1),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15_ (.A1(net2),
    .A2(_05_),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16_ (.A1(_10_),
    .A2(net1),
    .ZN(_06_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17_ (.A1(net5),
    .A2(_06_),
    .ZN(_07_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18_ (.A1(net2),
    .A2(_07_),
    .Z(_02_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19_ (.A1(net3),
    .A2(_11_),
    .A3(net1),
    .Z(_08_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20_ (.A1(net6),
    .A2(_08_),
    .Z(_09_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21_ (.A1(net2),
    .A2(_09_),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22_ (.A1(net5),
    .A2(net6),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _23_ (.A(net3),
    .B(net4),
    .CO(_10_),
    .S(net7));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _24_ (.A(net4),
    .B(net5),
    .CO(_11_),
    .S(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _25_ (.I(net6),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \binary_count[0]$_SDFFE_PN0P_  (.D(_00_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net3));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \binary_count[1]$_SDFFE_PN0P_  (.D(_01_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \binary_count[2]$_SDFFE_PN0P_  (.D(_02_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \binary_count[3]$_SDFFE_PN0P_  (.D(_03_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_57 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(enable),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(rst_n),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output3 (.I(net3),
    .Z(binary_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output4 (.I(net4),
    .Z(binary_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output5 (.I(net5),
    .Z(binary_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output6 (.I(net6),
    .Z(binary_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output7 (.I(net7),
    .Z(gray_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output8 (.I(net8),
    .Z(gray_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output9 (.I(net9),
    .Z(gray_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output10 (.I(net10),
    .Z(gray_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_218 ();
endmodule
