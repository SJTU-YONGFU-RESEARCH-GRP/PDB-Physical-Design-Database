module register_file (clk,
    read_en1,
    read_en2,
    rst_n,
    write_en,
    read_addr1,
    read_addr2,
    read_data1,
    read_data2,
    write_addr,
    write_data);
 input clk;
 input read_en1;
 input read_en2;
 input rst_n;
 input write_en;
 input [4:0] read_addr1;
 input [4:0] read_addr2;
 output [31:0] read_data1;
 output [31:0] read_data2;
 input [4:0] write_addr;
 input [31:0] write_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire \registers[0][0] ;
 wire \registers[0][10] ;
 wire \registers[0][11] ;
 wire \registers[0][12] ;
 wire \registers[0][13] ;
 wire \registers[0][14] ;
 wire \registers[0][15] ;
 wire \registers[0][16] ;
 wire \registers[0][17] ;
 wire \registers[0][18] ;
 wire \registers[0][19] ;
 wire \registers[0][1] ;
 wire \registers[0][20] ;
 wire \registers[0][21] ;
 wire \registers[0][22] ;
 wire \registers[0][23] ;
 wire \registers[0][24] ;
 wire \registers[0][25] ;
 wire \registers[0][26] ;
 wire \registers[0][27] ;
 wire \registers[0][28] ;
 wire \registers[0][29] ;
 wire \registers[0][2] ;
 wire \registers[0][30] ;
 wire \registers[0][31] ;
 wire \registers[0][3] ;
 wire \registers[0][4] ;
 wire \registers[0][5] ;
 wire \registers[0][6] ;
 wire \registers[0][7] ;
 wire \registers[0][8] ;
 wire \registers[0][9] ;
 wire \registers[10][0] ;
 wire \registers[10][10] ;
 wire \registers[10][11] ;
 wire \registers[10][12] ;
 wire \registers[10][13] ;
 wire \registers[10][14] ;
 wire \registers[10][15] ;
 wire \registers[10][16] ;
 wire \registers[10][17] ;
 wire \registers[10][18] ;
 wire \registers[10][19] ;
 wire \registers[10][1] ;
 wire \registers[10][20] ;
 wire \registers[10][21] ;
 wire \registers[10][22] ;
 wire \registers[10][23] ;
 wire \registers[10][24] ;
 wire \registers[10][25] ;
 wire \registers[10][26] ;
 wire \registers[10][27] ;
 wire \registers[10][28] ;
 wire \registers[10][29] ;
 wire \registers[10][2] ;
 wire \registers[10][30] ;
 wire \registers[10][31] ;
 wire \registers[10][3] ;
 wire \registers[10][4] ;
 wire \registers[10][5] ;
 wire \registers[10][6] ;
 wire \registers[10][7] ;
 wire \registers[10][8] ;
 wire \registers[10][9] ;
 wire \registers[11][0] ;
 wire \registers[11][10] ;
 wire \registers[11][11] ;
 wire \registers[11][12] ;
 wire \registers[11][13] ;
 wire \registers[11][14] ;
 wire \registers[11][15] ;
 wire \registers[11][16] ;
 wire \registers[11][17] ;
 wire \registers[11][18] ;
 wire \registers[11][19] ;
 wire \registers[11][1] ;
 wire \registers[11][20] ;
 wire \registers[11][21] ;
 wire \registers[11][22] ;
 wire \registers[11][23] ;
 wire \registers[11][24] ;
 wire \registers[11][25] ;
 wire \registers[11][26] ;
 wire \registers[11][27] ;
 wire \registers[11][28] ;
 wire \registers[11][29] ;
 wire \registers[11][2] ;
 wire \registers[11][30] ;
 wire \registers[11][31] ;
 wire \registers[11][3] ;
 wire \registers[11][4] ;
 wire \registers[11][5] ;
 wire \registers[11][6] ;
 wire \registers[11][7] ;
 wire \registers[11][8] ;
 wire \registers[11][9] ;
 wire \registers[12][0] ;
 wire \registers[12][10] ;
 wire \registers[12][11] ;
 wire \registers[12][12] ;
 wire \registers[12][13] ;
 wire \registers[12][14] ;
 wire \registers[12][15] ;
 wire \registers[12][16] ;
 wire \registers[12][17] ;
 wire \registers[12][18] ;
 wire \registers[12][19] ;
 wire \registers[12][1] ;
 wire \registers[12][20] ;
 wire \registers[12][21] ;
 wire \registers[12][22] ;
 wire \registers[12][23] ;
 wire \registers[12][24] ;
 wire \registers[12][25] ;
 wire \registers[12][26] ;
 wire \registers[12][27] ;
 wire \registers[12][28] ;
 wire \registers[12][29] ;
 wire \registers[12][2] ;
 wire \registers[12][30] ;
 wire \registers[12][31] ;
 wire \registers[12][3] ;
 wire \registers[12][4] ;
 wire \registers[12][5] ;
 wire \registers[12][6] ;
 wire \registers[12][7] ;
 wire \registers[12][8] ;
 wire \registers[12][9] ;
 wire \registers[13][0] ;
 wire \registers[13][10] ;
 wire \registers[13][11] ;
 wire \registers[13][12] ;
 wire \registers[13][13] ;
 wire \registers[13][14] ;
 wire \registers[13][15] ;
 wire \registers[13][16] ;
 wire \registers[13][17] ;
 wire \registers[13][18] ;
 wire \registers[13][19] ;
 wire \registers[13][1] ;
 wire \registers[13][20] ;
 wire \registers[13][21] ;
 wire \registers[13][22] ;
 wire \registers[13][23] ;
 wire \registers[13][24] ;
 wire \registers[13][25] ;
 wire \registers[13][26] ;
 wire \registers[13][27] ;
 wire \registers[13][28] ;
 wire \registers[13][29] ;
 wire \registers[13][2] ;
 wire \registers[13][30] ;
 wire \registers[13][31] ;
 wire \registers[13][3] ;
 wire \registers[13][4] ;
 wire \registers[13][5] ;
 wire \registers[13][6] ;
 wire \registers[13][7] ;
 wire \registers[13][8] ;
 wire \registers[13][9] ;
 wire \registers[14][0] ;
 wire \registers[14][10] ;
 wire \registers[14][11] ;
 wire \registers[14][12] ;
 wire \registers[14][13] ;
 wire \registers[14][14] ;
 wire \registers[14][15] ;
 wire \registers[14][16] ;
 wire \registers[14][17] ;
 wire \registers[14][18] ;
 wire \registers[14][19] ;
 wire \registers[14][1] ;
 wire \registers[14][20] ;
 wire \registers[14][21] ;
 wire \registers[14][22] ;
 wire \registers[14][23] ;
 wire \registers[14][24] ;
 wire \registers[14][25] ;
 wire \registers[14][26] ;
 wire \registers[14][27] ;
 wire \registers[14][28] ;
 wire \registers[14][29] ;
 wire \registers[14][2] ;
 wire \registers[14][30] ;
 wire \registers[14][31] ;
 wire \registers[14][3] ;
 wire \registers[14][4] ;
 wire \registers[14][5] ;
 wire \registers[14][6] ;
 wire \registers[14][7] ;
 wire \registers[14][8] ;
 wire \registers[14][9] ;
 wire \registers[15][0] ;
 wire \registers[15][10] ;
 wire \registers[15][11] ;
 wire \registers[15][12] ;
 wire \registers[15][13] ;
 wire \registers[15][14] ;
 wire \registers[15][15] ;
 wire \registers[15][16] ;
 wire \registers[15][17] ;
 wire \registers[15][18] ;
 wire \registers[15][19] ;
 wire \registers[15][1] ;
 wire \registers[15][20] ;
 wire \registers[15][21] ;
 wire \registers[15][22] ;
 wire \registers[15][23] ;
 wire \registers[15][24] ;
 wire \registers[15][25] ;
 wire \registers[15][26] ;
 wire \registers[15][27] ;
 wire \registers[15][28] ;
 wire \registers[15][29] ;
 wire \registers[15][2] ;
 wire \registers[15][30] ;
 wire \registers[15][31] ;
 wire \registers[15][3] ;
 wire \registers[15][4] ;
 wire \registers[15][5] ;
 wire \registers[15][6] ;
 wire \registers[15][7] ;
 wire \registers[15][8] ;
 wire \registers[15][9] ;
 wire \registers[16][0] ;
 wire \registers[16][10] ;
 wire \registers[16][11] ;
 wire \registers[16][12] ;
 wire \registers[16][13] ;
 wire \registers[16][14] ;
 wire \registers[16][15] ;
 wire \registers[16][16] ;
 wire \registers[16][17] ;
 wire \registers[16][18] ;
 wire \registers[16][19] ;
 wire \registers[16][1] ;
 wire \registers[16][20] ;
 wire \registers[16][21] ;
 wire \registers[16][22] ;
 wire \registers[16][23] ;
 wire \registers[16][24] ;
 wire \registers[16][25] ;
 wire \registers[16][26] ;
 wire \registers[16][27] ;
 wire \registers[16][28] ;
 wire \registers[16][29] ;
 wire \registers[16][2] ;
 wire \registers[16][30] ;
 wire \registers[16][31] ;
 wire \registers[16][3] ;
 wire \registers[16][4] ;
 wire \registers[16][5] ;
 wire \registers[16][6] ;
 wire \registers[16][7] ;
 wire \registers[16][8] ;
 wire \registers[16][9] ;
 wire \registers[17][0] ;
 wire \registers[17][10] ;
 wire \registers[17][11] ;
 wire \registers[17][12] ;
 wire \registers[17][13] ;
 wire \registers[17][14] ;
 wire \registers[17][15] ;
 wire \registers[17][16] ;
 wire \registers[17][17] ;
 wire \registers[17][18] ;
 wire \registers[17][19] ;
 wire \registers[17][1] ;
 wire \registers[17][20] ;
 wire \registers[17][21] ;
 wire \registers[17][22] ;
 wire \registers[17][23] ;
 wire \registers[17][24] ;
 wire \registers[17][25] ;
 wire \registers[17][26] ;
 wire \registers[17][27] ;
 wire \registers[17][28] ;
 wire \registers[17][29] ;
 wire \registers[17][2] ;
 wire \registers[17][30] ;
 wire \registers[17][31] ;
 wire \registers[17][3] ;
 wire \registers[17][4] ;
 wire \registers[17][5] ;
 wire \registers[17][6] ;
 wire \registers[17][7] ;
 wire \registers[17][8] ;
 wire \registers[17][9] ;
 wire \registers[18][0] ;
 wire \registers[18][10] ;
 wire \registers[18][11] ;
 wire \registers[18][12] ;
 wire \registers[18][13] ;
 wire \registers[18][14] ;
 wire \registers[18][15] ;
 wire \registers[18][16] ;
 wire \registers[18][17] ;
 wire \registers[18][18] ;
 wire \registers[18][19] ;
 wire \registers[18][1] ;
 wire \registers[18][20] ;
 wire \registers[18][21] ;
 wire \registers[18][22] ;
 wire \registers[18][23] ;
 wire \registers[18][24] ;
 wire \registers[18][25] ;
 wire \registers[18][26] ;
 wire \registers[18][27] ;
 wire \registers[18][28] ;
 wire \registers[18][29] ;
 wire \registers[18][2] ;
 wire \registers[18][30] ;
 wire \registers[18][31] ;
 wire \registers[18][3] ;
 wire \registers[18][4] ;
 wire \registers[18][5] ;
 wire \registers[18][6] ;
 wire \registers[18][7] ;
 wire \registers[18][8] ;
 wire \registers[18][9] ;
 wire \registers[19][0] ;
 wire \registers[19][10] ;
 wire \registers[19][11] ;
 wire \registers[19][12] ;
 wire \registers[19][13] ;
 wire \registers[19][14] ;
 wire \registers[19][15] ;
 wire \registers[19][16] ;
 wire \registers[19][17] ;
 wire \registers[19][18] ;
 wire \registers[19][19] ;
 wire \registers[19][1] ;
 wire \registers[19][20] ;
 wire \registers[19][21] ;
 wire \registers[19][22] ;
 wire \registers[19][23] ;
 wire \registers[19][24] ;
 wire \registers[19][25] ;
 wire \registers[19][26] ;
 wire \registers[19][27] ;
 wire \registers[19][28] ;
 wire \registers[19][29] ;
 wire \registers[19][2] ;
 wire \registers[19][30] ;
 wire \registers[19][31] ;
 wire \registers[19][3] ;
 wire \registers[19][4] ;
 wire \registers[19][5] ;
 wire \registers[19][6] ;
 wire \registers[19][7] ;
 wire \registers[19][8] ;
 wire \registers[19][9] ;
 wire \registers[1][0] ;
 wire \registers[1][10] ;
 wire \registers[1][11] ;
 wire \registers[1][12] ;
 wire \registers[1][13] ;
 wire \registers[1][14] ;
 wire \registers[1][15] ;
 wire \registers[1][16] ;
 wire \registers[1][17] ;
 wire \registers[1][18] ;
 wire \registers[1][19] ;
 wire \registers[1][1] ;
 wire \registers[1][20] ;
 wire \registers[1][21] ;
 wire \registers[1][22] ;
 wire \registers[1][23] ;
 wire \registers[1][24] ;
 wire \registers[1][25] ;
 wire \registers[1][26] ;
 wire \registers[1][27] ;
 wire \registers[1][28] ;
 wire \registers[1][29] ;
 wire \registers[1][2] ;
 wire \registers[1][30] ;
 wire \registers[1][31] ;
 wire \registers[1][3] ;
 wire \registers[1][4] ;
 wire \registers[1][5] ;
 wire \registers[1][6] ;
 wire \registers[1][7] ;
 wire \registers[1][8] ;
 wire \registers[1][9] ;
 wire \registers[20][0] ;
 wire \registers[20][10] ;
 wire \registers[20][11] ;
 wire \registers[20][12] ;
 wire \registers[20][13] ;
 wire \registers[20][14] ;
 wire \registers[20][15] ;
 wire \registers[20][16] ;
 wire \registers[20][17] ;
 wire \registers[20][18] ;
 wire \registers[20][19] ;
 wire \registers[20][1] ;
 wire \registers[20][20] ;
 wire \registers[20][21] ;
 wire \registers[20][22] ;
 wire \registers[20][23] ;
 wire \registers[20][24] ;
 wire \registers[20][25] ;
 wire \registers[20][26] ;
 wire \registers[20][27] ;
 wire \registers[20][28] ;
 wire \registers[20][29] ;
 wire \registers[20][2] ;
 wire \registers[20][30] ;
 wire \registers[20][31] ;
 wire \registers[20][3] ;
 wire \registers[20][4] ;
 wire \registers[20][5] ;
 wire \registers[20][6] ;
 wire \registers[20][7] ;
 wire \registers[20][8] ;
 wire \registers[20][9] ;
 wire \registers[21][0] ;
 wire \registers[21][10] ;
 wire \registers[21][11] ;
 wire \registers[21][12] ;
 wire \registers[21][13] ;
 wire \registers[21][14] ;
 wire \registers[21][15] ;
 wire \registers[21][16] ;
 wire \registers[21][17] ;
 wire \registers[21][18] ;
 wire \registers[21][19] ;
 wire \registers[21][1] ;
 wire \registers[21][20] ;
 wire \registers[21][21] ;
 wire \registers[21][22] ;
 wire \registers[21][23] ;
 wire \registers[21][24] ;
 wire \registers[21][25] ;
 wire \registers[21][26] ;
 wire \registers[21][27] ;
 wire \registers[21][28] ;
 wire \registers[21][29] ;
 wire \registers[21][2] ;
 wire \registers[21][30] ;
 wire \registers[21][31] ;
 wire \registers[21][3] ;
 wire \registers[21][4] ;
 wire \registers[21][5] ;
 wire \registers[21][6] ;
 wire \registers[21][7] ;
 wire \registers[21][8] ;
 wire \registers[21][9] ;
 wire \registers[22][0] ;
 wire \registers[22][10] ;
 wire \registers[22][11] ;
 wire \registers[22][12] ;
 wire \registers[22][13] ;
 wire \registers[22][14] ;
 wire \registers[22][15] ;
 wire \registers[22][16] ;
 wire \registers[22][17] ;
 wire \registers[22][18] ;
 wire \registers[22][19] ;
 wire \registers[22][1] ;
 wire \registers[22][20] ;
 wire \registers[22][21] ;
 wire \registers[22][22] ;
 wire \registers[22][23] ;
 wire \registers[22][24] ;
 wire \registers[22][25] ;
 wire \registers[22][26] ;
 wire \registers[22][27] ;
 wire \registers[22][28] ;
 wire \registers[22][29] ;
 wire \registers[22][2] ;
 wire \registers[22][30] ;
 wire \registers[22][31] ;
 wire \registers[22][3] ;
 wire \registers[22][4] ;
 wire \registers[22][5] ;
 wire \registers[22][6] ;
 wire \registers[22][7] ;
 wire \registers[22][8] ;
 wire \registers[22][9] ;
 wire \registers[23][0] ;
 wire \registers[23][10] ;
 wire \registers[23][11] ;
 wire \registers[23][12] ;
 wire \registers[23][13] ;
 wire \registers[23][14] ;
 wire \registers[23][15] ;
 wire \registers[23][16] ;
 wire \registers[23][17] ;
 wire \registers[23][18] ;
 wire \registers[23][19] ;
 wire \registers[23][1] ;
 wire \registers[23][20] ;
 wire \registers[23][21] ;
 wire \registers[23][22] ;
 wire \registers[23][23] ;
 wire \registers[23][24] ;
 wire \registers[23][25] ;
 wire \registers[23][26] ;
 wire \registers[23][27] ;
 wire \registers[23][28] ;
 wire \registers[23][29] ;
 wire \registers[23][2] ;
 wire \registers[23][30] ;
 wire \registers[23][31] ;
 wire \registers[23][3] ;
 wire \registers[23][4] ;
 wire \registers[23][5] ;
 wire \registers[23][6] ;
 wire \registers[23][7] ;
 wire \registers[23][8] ;
 wire \registers[23][9] ;
 wire \registers[24][0] ;
 wire \registers[24][10] ;
 wire \registers[24][11] ;
 wire \registers[24][12] ;
 wire \registers[24][13] ;
 wire \registers[24][14] ;
 wire \registers[24][15] ;
 wire \registers[24][16] ;
 wire \registers[24][17] ;
 wire \registers[24][18] ;
 wire \registers[24][19] ;
 wire \registers[24][1] ;
 wire \registers[24][20] ;
 wire \registers[24][21] ;
 wire \registers[24][22] ;
 wire \registers[24][23] ;
 wire \registers[24][24] ;
 wire \registers[24][25] ;
 wire \registers[24][26] ;
 wire \registers[24][27] ;
 wire \registers[24][28] ;
 wire \registers[24][29] ;
 wire \registers[24][2] ;
 wire \registers[24][30] ;
 wire \registers[24][31] ;
 wire \registers[24][3] ;
 wire \registers[24][4] ;
 wire \registers[24][5] ;
 wire \registers[24][6] ;
 wire \registers[24][7] ;
 wire \registers[24][8] ;
 wire \registers[24][9] ;
 wire \registers[25][0] ;
 wire \registers[25][10] ;
 wire \registers[25][11] ;
 wire \registers[25][12] ;
 wire \registers[25][13] ;
 wire \registers[25][14] ;
 wire \registers[25][15] ;
 wire \registers[25][16] ;
 wire \registers[25][17] ;
 wire \registers[25][18] ;
 wire \registers[25][19] ;
 wire \registers[25][1] ;
 wire \registers[25][20] ;
 wire \registers[25][21] ;
 wire \registers[25][22] ;
 wire \registers[25][23] ;
 wire \registers[25][24] ;
 wire \registers[25][25] ;
 wire \registers[25][26] ;
 wire \registers[25][27] ;
 wire \registers[25][28] ;
 wire \registers[25][29] ;
 wire \registers[25][2] ;
 wire \registers[25][30] ;
 wire \registers[25][31] ;
 wire \registers[25][3] ;
 wire \registers[25][4] ;
 wire \registers[25][5] ;
 wire \registers[25][6] ;
 wire \registers[25][7] ;
 wire \registers[25][8] ;
 wire \registers[25][9] ;
 wire \registers[26][0] ;
 wire \registers[26][10] ;
 wire \registers[26][11] ;
 wire \registers[26][12] ;
 wire \registers[26][13] ;
 wire \registers[26][14] ;
 wire \registers[26][15] ;
 wire \registers[26][16] ;
 wire \registers[26][17] ;
 wire \registers[26][18] ;
 wire \registers[26][19] ;
 wire \registers[26][1] ;
 wire \registers[26][20] ;
 wire \registers[26][21] ;
 wire \registers[26][22] ;
 wire \registers[26][23] ;
 wire \registers[26][24] ;
 wire \registers[26][25] ;
 wire \registers[26][26] ;
 wire \registers[26][27] ;
 wire \registers[26][28] ;
 wire \registers[26][29] ;
 wire \registers[26][2] ;
 wire \registers[26][30] ;
 wire \registers[26][31] ;
 wire \registers[26][3] ;
 wire \registers[26][4] ;
 wire \registers[26][5] ;
 wire \registers[26][6] ;
 wire \registers[26][7] ;
 wire \registers[26][8] ;
 wire \registers[26][9] ;
 wire \registers[27][0] ;
 wire \registers[27][10] ;
 wire \registers[27][11] ;
 wire \registers[27][12] ;
 wire \registers[27][13] ;
 wire \registers[27][14] ;
 wire \registers[27][15] ;
 wire \registers[27][16] ;
 wire \registers[27][17] ;
 wire \registers[27][18] ;
 wire \registers[27][19] ;
 wire \registers[27][1] ;
 wire \registers[27][20] ;
 wire \registers[27][21] ;
 wire \registers[27][22] ;
 wire \registers[27][23] ;
 wire \registers[27][24] ;
 wire \registers[27][25] ;
 wire \registers[27][26] ;
 wire \registers[27][27] ;
 wire \registers[27][28] ;
 wire \registers[27][29] ;
 wire \registers[27][2] ;
 wire \registers[27][30] ;
 wire \registers[27][31] ;
 wire \registers[27][3] ;
 wire \registers[27][4] ;
 wire \registers[27][5] ;
 wire \registers[27][6] ;
 wire \registers[27][7] ;
 wire \registers[27][8] ;
 wire \registers[27][9] ;
 wire \registers[28][0] ;
 wire \registers[28][10] ;
 wire \registers[28][11] ;
 wire \registers[28][12] ;
 wire \registers[28][13] ;
 wire \registers[28][14] ;
 wire \registers[28][15] ;
 wire \registers[28][16] ;
 wire \registers[28][17] ;
 wire \registers[28][18] ;
 wire \registers[28][19] ;
 wire \registers[28][1] ;
 wire \registers[28][20] ;
 wire \registers[28][21] ;
 wire \registers[28][22] ;
 wire \registers[28][23] ;
 wire \registers[28][24] ;
 wire \registers[28][25] ;
 wire \registers[28][26] ;
 wire \registers[28][27] ;
 wire \registers[28][28] ;
 wire \registers[28][29] ;
 wire \registers[28][2] ;
 wire \registers[28][30] ;
 wire \registers[28][31] ;
 wire \registers[28][3] ;
 wire \registers[28][4] ;
 wire \registers[28][5] ;
 wire \registers[28][6] ;
 wire \registers[28][7] ;
 wire \registers[28][8] ;
 wire \registers[28][9] ;
 wire \registers[29][0] ;
 wire \registers[29][10] ;
 wire \registers[29][11] ;
 wire \registers[29][12] ;
 wire \registers[29][13] ;
 wire \registers[29][14] ;
 wire \registers[29][15] ;
 wire \registers[29][16] ;
 wire \registers[29][17] ;
 wire \registers[29][18] ;
 wire \registers[29][19] ;
 wire \registers[29][1] ;
 wire \registers[29][20] ;
 wire \registers[29][21] ;
 wire \registers[29][22] ;
 wire \registers[29][23] ;
 wire \registers[29][24] ;
 wire \registers[29][25] ;
 wire \registers[29][26] ;
 wire \registers[29][27] ;
 wire \registers[29][28] ;
 wire \registers[29][29] ;
 wire \registers[29][2] ;
 wire \registers[29][30] ;
 wire \registers[29][31] ;
 wire \registers[29][3] ;
 wire \registers[29][4] ;
 wire \registers[29][5] ;
 wire \registers[29][6] ;
 wire \registers[29][7] ;
 wire \registers[29][8] ;
 wire \registers[29][9] ;
 wire \registers[2][0] ;
 wire \registers[2][10] ;
 wire \registers[2][11] ;
 wire \registers[2][12] ;
 wire \registers[2][13] ;
 wire \registers[2][14] ;
 wire \registers[2][15] ;
 wire \registers[2][16] ;
 wire \registers[2][17] ;
 wire \registers[2][18] ;
 wire \registers[2][19] ;
 wire \registers[2][1] ;
 wire \registers[2][20] ;
 wire \registers[2][21] ;
 wire \registers[2][22] ;
 wire \registers[2][23] ;
 wire \registers[2][24] ;
 wire \registers[2][25] ;
 wire \registers[2][26] ;
 wire \registers[2][27] ;
 wire \registers[2][28] ;
 wire \registers[2][29] ;
 wire \registers[2][2] ;
 wire \registers[2][30] ;
 wire \registers[2][31] ;
 wire \registers[2][3] ;
 wire \registers[2][4] ;
 wire \registers[2][5] ;
 wire \registers[2][6] ;
 wire \registers[2][7] ;
 wire \registers[2][8] ;
 wire \registers[2][9] ;
 wire \registers[30][0] ;
 wire \registers[30][10] ;
 wire \registers[30][11] ;
 wire \registers[30][12] ;
 wire \registers[30][13] ;
 wire \registers[30][14] ;
 wire \registers[30][15] ;
 wire \registers[30][16] ;
 wire \registers[30][17] ;
 wire \registers[30][18] ;
 wire \registers[30][19] ;
 wire \registers[30][1] ;
 wire \registers[30][20] ;
 wire \registers[30][21] ;
 wire \registers[30][22] ;
 wire \registers[30][23] ;
 wire \registers[30][24] ;
 wire \registers[30][25] ;
 wire \registers[30][26] ;
 wire \registers[30][27] ;
 wire \registers[30][28] ;
 wire \registers[30][29] ;
 wire \registers[30][2] ;
 wire \registers[30][30] ;
 wire \registers[30][31] ;
 wire \registers[30][3] ;
 wire \registers[30][4] ;
 wire \registers[30][5] ;
 wire \registers[30][6] ;
 wire \registers[30][7] ;
 wire \registers[30][8] ;
 wire \registers[30][9] ;
 wire \registers[31][0] ;
 wire \registers[31][10] ;
 wire \registers[31][11] ;
 wire \registers[31][12] ;
 wire \registers[31][13] ;
 wire \registers[31][14] ;
 wire \registers[31][15] ;
 wire \registers[31][16] ;
 wire \registers[31][17] ;
 wire \registers[31][18] ;
 wire \registers[31][19] ;
 wire \registers[31][1] ;
 wire \registers[31][20] ;
 wire \registers[31][21] ;
 wire \registers[31][22] ;
 wire \registers[31][23] ;
 wire \registers[31][24] ;
 wire \registers[31][25] ;
 wire \registers[31][26] ;
 wire \registers[31][27] ;
 wire \registers[31][28] ;
 wire \registers[31][29] ;
 wire \registers[31][2] ;
 wire \registers[31][30] ;
 wire \registers[31][31] ;
 wire \registers[31][3] ;
 wire \registers[31][4] ;
 wire \registers[31][5] ;
 wire \registers[31][6] ;
 wire \registers[31][7] ;
 wire \registers[31][8] ;
 wire \registers[31][9] ;
 wire \registers[3][0] ;
 wire \registers[3][10] ;
 wire \registers[3][11] ;
 wire \registers[3][12] ;
 wire \registers[3][13] ;
 wire \registers[3][14] ;
 wire \registers[3][15] ;
 wire \registers[3][16] ;
 wire \registers[3][17] ;
 wire \registers[3][18] ;
 wire \registers[3][19] ;
 wire \registers[3][1] ;
 wire \registers[3][20] ;
 wire \registers[3][21] ;
 wire \registers[3][22] ;
 wire \registers[3][23] ;
 wire \registers[3][24] ;
 wire \registers[3][25] ;
 wire \registers[3][26] ;
 wire \registers[3][27] ;
 wire \registers[3][28] ;
 wire \registers[3][29] ;
 wire \registers[3][2] ;
 wire \registers[3][30] ;
 wire \registers[3][31] ;
 wire \registers[3][3] ;
 wire \registers[3][4] ;
 wire \registers[3][5] ;
 wire \registers[3][6] ;
 wire \registers[3][7] ;
 wire \registers[3][8] ;
 wire \registers[3][9] ;
 wire \registers[4][0] ;
 wire \registers[4][10] ;
 wire \registers[4][11] ;
 wire \registers[4][12] ;
 wire \registers[4][13] ;
 wire \registers[4][14] ;
 wire \registers[4][15] ;
 wire \registers[4][16] ;
 wire \registers[4][17] ;
 wire \registers[4][18] ;
 wire \registers[4][19] ;
 wire \registers[4][1] ;
 wire \registers[4][20] ;
 wire \registers[4][21] ;
 wire \registers[4][22] ;
 wire \registers[4][23] ;
 wire \registers[4][24] ;
 wire \registers[4][25] ;
 wire \registers[4][26] ;
 wire \registers[4][27] ;
 wire \registers[4][28] ;
 wire \registers[4][29] ;
 wire \registers[4][2] ;
 wire \registers[4][30] ;
 wire \registers[4][31] ;
 wire \registers[4][3] ;
 wire \registers[4][4] ;
 wire \registers[4][5] ;
 wire \registers[4][6] ;
 wire \registers[4][7] ;
 wire \registers[4][8] ;
 wire \registers[4][9] ;
 wire \registers[5][0] ;
 wire \registers[5][10] ;
 wire \registers[5][11] ;
 wire \registers[5][12] ;
 wire \registers[5][13] ;
 wire \registers[5][14] ;
 wire \registers[5][15] ;
 wire \registers[5][16] ;
 wire \registers[5][17] ;
 wire \registers[5][18] ;
 wire \registers[5][19] ;
 wire \registers[5][1] ;
 wire \registers[5][20] ;
 wire \registers[5][21] ;
 wire \registers[5][22] ;
 wire \registers[5][23] ;
 wire \registers[5][24] ;
 wire \registers[5][25] ;
 wire \registers[5][26] ;
 wire \registers[5][27] ;
 wire \registers[5][28] ;
 wire \registers[5][29] ;
 wire \registers[5][2] ;
 wire \registers[5][30] ;
 wire \registers[5][31] ;
 wire \registers[5][3] ;
 wire \registers[5][4] ;
 wire \registers[5][5] ;
 wire \registers[5][6] ;
 wire \registers[5][7] ;
 wire \registers[5][8] ;
 wire \registers[5][9] ;
 wire \registers[6][0] ;
 wire \registers[6][10] ;
 wire \registers[6][11] ;
 wire \registers[6][12] ;
 wire \registers[6][13] ;
 wire \registers[6][14] ;
 wire \registers[6][15] ;
 wire \registers[6][16] ;
 wire \registers[6][17] ;
 wire \registers[6][18] ;
 wire \registers[6][19] ;
 wire \registers[6][1] ;
 wire \registers[6][20] ;
 wire \registers[6][21] ;
 wire \registers[6][22] ;
 wire \registers[6][23] ;
 wire \registers[6][24] ;
 wire \registers[6][25] ;
 wire \registers[6][26] ;
 wire \registers[6][27] ;
 wire \registers[6][28] ;
 wire \registers[6][29] ;
 wire \registers[6][2] ;
 wire \registers[6][30] ;
 wire \registers[6][31] ;
 wire \registers[6][3] ;
 wire \registers[6][4] ;
 wire \registers[6][5] ;
 wire \registers[6][6] ;
 wire \registers[6][7] ;
 wire \registers[6][8] ;
 wire \registers[6][9] ;
 wire \registers[7][0] ;
 wire \registers[7][10] ;
 wire \registers[7][11] ;
 wire \registers[7][12] ;
 wire \registers[7][13] ;
 wire \registers[7][14] ;
 wire \registers[7][15] ;
 wire \registers[7][16] ;
 wire \registers[7][17] ;
 wire \registers[7][18] ;
 wire \registers[7][19] ;
 wire \registers[7][1] ;
 wire \registers[7][20] ;
 wire \registers[7][21] ;
 wire \registers[7][22] ;
 wire \registers[7][23] ;
 wire \registers[7][24] ;
 wire \registers[7][25] ;
 wire \registers[7][26] ;
 wire \registers[7][27] ;
 wire \registers[7][28] ;
 wire \registers[7][29] ;
 wire \registers[7][2] ;
 wire \registers[7][30] ;
 wire \registers[7][31] ;
 wire \registers[7][3] ;
 wire \registers[7][4] ;
 wire \registers[7][5] ;
 wire \registers[7][6] ;
 wire \registers[7][7] ;
 wire \registers[7][8] ;
 wire \registers[7][9] ;
 wire \registers[8][0] ;
 wire \registers[8][10] ;
 wire \registers[8][11] ;
 wire \registers[8][12] ;
 wire \registers[8][13] ;
 wire \registers[8][14] ;
 wire \registers[8][15] ;
 wire \registers[8][16] ;
 wire \registers[8][17] ;
 wire \registers[8][18] ;
 wire \registers[8][19] ;
 wire \registers[8][1] ;
 wire \registers[8][20] ;
 wire \registers[8][21] ;
 wire \registers[8][22] ;
 wire \registers[8][23] ;
 wire \registers[8][24] ;
 wire \registers[8][25] ;
 wire \registers[8][26] ;
 wire \registers[8][27] ;
 wire \registers[8][28] ;
 wire \registers[8][29] ;
 wire \registers[8][2] ;
 wire \registers[8][30] ;
 wire \registers[8][31] ;
 wire \registers[8][3] ;
 wire \registers[8][4] ;
 wire \registers[8][5] ;
 wire \registers[8][6] ;
 wire \registers[8][7] ;
 wire \registers[8][8] ;
 wire \registers[8][9] ;
 wire \registers[9][0] ;
 wire \registers[9][10] ;
 wire \registers[9][11] ;
 wire \registers[9][12] ;
 wire \registers[9][13] ;
 wire \registers[9][14] ;
 wire \registers[9][15] ;
 wire \registers[9][16] ;
 wire \registers[9][17] ;
 wire \registers[9][18] ;
 wire \registers[9][19] ;
 wire \registers[9][1] ;
 wire \registers[9][20] ;
 wire \registers[9][21] ;
 wire \registers[9][22] ;
 wire \registers[9][23] ;
 wire \registers[9][24] ;
 wire \registers[9][25] ;
 wire \registers[9][26] ;
 wire \registers[9][27] ;
 wire \registers[9][28] ;
 wire \registers[9][29] ;
 wire \registers[9][2] ;
 wire \registers[9][30] ;
 wire \registers[9][31] ;
 wire \registers[9][3] ;
 wire \registers[9][4] ;
 wire \registers[9][5] ;
 wire \registers[9][6] ;
 wire \registers[9][7] ;
 wire \registers[9][8] ;
 wire \registers[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;

 sky130_fd_sc_hd__a221oi_2 _2566_ (.A1(_1828_),
    .A2(_1910_),
    .B1(_1911_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_1912_));
 sky130_fd_sc_hd__o21ai_0 _2567_ (.A1(_1800_),
    .A2(_1909_),
    .B1(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__mux4_1 _2568_ (.A0(\registers[24][15] ),
    .A1(\registers[26][15] ),
    .A2(\registers[28][15] ),
    .A3(\registers[30][15] ),
    .S0(_1764_),
    .S1(_1877_),
    .X(_1914_));
 sky130_fd_sc_hd__mux4_1 _2569_ (.A0(\registers[25][15] ),
    .A1(\registers[27][15] ),
    .A2(\registers[29][15] ),
    .A3(\registers[31][15] ),
    .S0(_1839_),
    .S1(_1879_),
    .X(_1915_));
 sky130_fd_sc_hd__a22oi_2 _2570_ (.A1(_1836_),
    .A2(_1914_),
    .B1(_1915_),
    .B2(_1812_),
    .Y(_1916_));
 sky130_fd_sc_hd__mux4_1 _2571_ (.A0(\registers[8][15] ),
    .A1(\registers[9][15] ),
    .A2(\registers[10][15] ),
    .A3(\registers[11][15] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_1917_));
 sky130_fd_sc_hd__mux4_1 _2572_ (.A0(\registers[12][15] ),
    .A1(\registers[13][15] ),
    .A2(\registers[14][15] ),
    .A3(\registers[15][15] ),
    .S0(_1862_),
    .S1(_1816_),
    .X(_1918_));
 sky130_fd_sc_hd__mux2i_2 _2573_ (.A0(_1917_),
    .A1(_1918_),
    .S(_1845_),
    .Y(_1919_));
 sky130_fd_sc_hd__mux4_1 _2574_ (.A0(\registers[1][15] ),
    .A1(\registers[3][15] ),
    .A2(\registers[5][15] ),
    .A3(\registers[7][15] ),
    .S0(_1865_),
    .S1(_1885_),
    .X(_1920_));
 sky130_fd_sc_hd__mux4_1 _2575_ (.A0(\registers[0][15] ),
    .A1(\registers[2][15] ),
    .A2(\registers[4][15] ),
    .A3(\registers[6][15] ),
    .S0(_1848_),
    .S1(_1867_),
    .X(_1921_));
 sky130_fd_sc_hd__mux2i_1 _2576_ (.A0(_1920_),
    .A1(_1921_),
    .S(_1750_),
    .Y(_1922_));
 sky130_fd_sc_hd__buf_8 _2577_ (.A(_1792_),
    .X(_1923_));
 sky130_fd_sc_hd__a221o_2 _2578_ (.A1(_1785_),
    .A2(_1919_),
    .B1(_1922_),
    .B2(_1923_),
    .C1(_1798_),
    .X(_1924_));
 sky130_fd_sc_hd__a31oi_1 _2579_ (.A1(_1746_),
    .A2(_1913_),
    .A3(_1916_),
    .B1(_1924_),
    .Y(_0072_));
 sky130_fd_sc_hd__mux4_1 _2580_ (.A0(\registers[17][16] ),
    .A1(\registers[19][16] ),
    .A2(\registers[21][16] ),
    .A3(\registers[23][16] ),
    .S0(_1801_),
    .S1(_1871_),
    .X(_1925_));
 sky130_fd_sc_hd__mux2i_1 _2581_ (.A0(\registers[18][16] ),
    .A1(\registers[22][16] ),
    .S(_1829_),
    .Y(_1926_));
 sky130_fd_sc_hd__mux2i_1 _2582_ (.A0(\registers[16][16] ),
    .A1(\registers[20][16] ),
    .S(_1776_),
    .Y(_1927_));
 sky130_fd_sc_hd__a221oi_1 _2583_ (.A1(_1828_),
    .A2(_1926_),
    .B1(_1927_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_1928_));
 sky130_fd_sc_hd__o21ai_0 _2584_ (.A1(_1800_),
    .A2(_1925_),
    .B1(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__mux4_1 _2585_ (.A0(\registers[24][16] ),
    .A1(\registers[26][16] ),
    .A2(\registers[28][16] ),
    .A3(\registers[30][16] ),
    .S0(_1764_),
    .S1(_1877_),
    .X(_1930_));
 sky130_fd_sc_hd__mux4_1 _2586_ (.A0(\registers[25][16] ),
    .A1(\registers[27][16] ),
    .A2(\registers[29][16] ),
    .A3(\registers[31][16] ),
    .S0(_1839_),
    .S1(_1879_),
    .X(_1931_));
 sky130_fd_sc_hd__a22oi_2 _2587_ (.A1(_1836_),
    .A2(_1930_),
    .B1(_1931_),
    .B2(_1812_),
    .Y(_1932_));
 sky130_fd_sc_hd__mux4_1 _2588_ (.A0(\registers[0][16] ),
    .A1(\registers[1][16] ),
    .A2(\registers[2][16] ),
    .A3(\registers[3][16] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_1933_));
 sky130_fd_sc_hd__mux4_1 _2589_ (.A0(\registers[4][16] ),
    .A1(\registers[5][16] ),
    .A2(\registers[6][16] ),
    .A3(\registers[7][16] ),
    .S0(_1862_),
    .S1(_1816_),
    .X(_1934_));
 sky130_fd_sc_hd__mux2i_1 _2590_ (.A0(_1933_),
    .A1(_1934_),
    .S(_1845_),
    .Y(_1935_));
 sky130_fd_sc_hd__mux4_1 _2591_ (.A0(\registers[9][16] ),
    .A1(\registers[11][16] ),
    .A2(\registers[13][16] ),
    .A3(\registers[15][16] ),
    .S0(_1865_),
    .S1(_1885_),
    .X(_1936_));
 sky130_fd_sc_hd__mux4_1 _2592_ (.A0(\registers[8][16] ),
    .A1(\registers[10][16] ),
    .A2(\registers[12][16] ),
    .A3(\registers[14][16] ),
    .S0(_1848_),
    .S1(_1867_),
    .X(_1937_));
 sky130_fd_sc_hd__buf_16 _2593_ (.A(_1749_),
    .X(_1938_));
 sky130_fd_sc_hd__mux2i_4 _2594_ (.A0(_1936_),
    .A1(_1937_),
    .S(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__a221o_2 _2595_ (.A1(_1793_),
    .A2(_1935_),
    .B1(_1939_),
    .B2(_1825_),
    .C1(_1798_),
    .X(_1940_));
 sky130_fd_sc_hd__a31oi_1 _2596_ (.A1(_1746_),
    .A2(_1929_),
    .A3(_1932_),
    .B1(_1940_),
    .Y(_0073_));
 sky130_fd_sc_hd__mux4_1 _2597_ (.A0(\registers[17][17] ),
    .A1(\registers[19][17] ),
    .A2(\registers[21][17] ),
    .A3(\registers[23][17] ),
    .S0(_1801_),
    .S1(_1871_),
    .X(_1941_));
 sky130_fd_sc_hd__mux2i_1 _2598_ (.A0(\registers[18][17] ),
    .A1(\registers[22][17] ),
    .S(_1829_),
    .Y(_1942_));
 sky130_fd_sc_hd__buf_6 _2599_ (.A(_1819_),
    .X(_1943_));
 sky130_fd_sc_hd__mux2i_1 _2600_ (.A0(\registers[16][17] ),
    .A1(\registers[20][17] ),
    .S(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__a221oi_2 _2601_ (.A1(_1828_),
    .A2(_1942_),
    .B1(_1944_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_1945_));
 sky130_fd_sc_hd__o21ai_0 _2602_ (.A1(_1800_),
    .A2(_1941_),
    .B1(_1945_),
    .Y(_1946_));
 sky130_fd_sc_hd__mux4_1 _2603_ (.A0(\registers[24][17] ),
    .A1(\registers[26][17] ),
    .A2(\registers[28][17] ),
    .A3(\registers[30][17] ),
    .S0(_1764_),
    .S1(_1877_),
    .X(_1947_));
 sky130_fd_sc_hd__mux4_1 _2604_ (.A0(\registers[25][17] ),
    .A1(\registers[27][17] ),
    .A2(\registers[29][17] ),
    .A3(\registers[31][17] ),
    .S0(_1839_),
    .S1(_1879_),
    .X(_1948_));
 sky130_fd_sc_hd__a22oi_2 _2605_ (.A1(_1836_),
    .A2(_1947_),
    .B1(_1948_),
    .B2(_1812_),
    .Y(_1949_));
 sky130_fd_sc_hd__mux4_1 _2606_ (.A0(\registers[8][17] ),
    .A1(\registers[9][17] ),
    .A2(\registers[10][17] ),
    .A3(\registers[11][17] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_1950_));
 sky130_fd_sc_hd__mux4_1 _2607_ (.A0(\registers[12][17] ),
    .A1(\registers[13][17] ),
    .A2(\registers[14][17] ),
    .A3(\registers[15][17] ),
    .S0(_1862_),
    .S1(_1816_),
    .X(_1951_));
 sky130_fd_sc_hd__mux2i_2 _2608_ (.A0(_1950_),
    .A1(_1951_),
    .S(_1845_),
    .Y(_1952_));
 sky130_fd_sc_hd__mux4_1 _2609_ (.A0(\registers[1][17] ),
    .A1(\registers[3][17] ),
    .A2(\registers[5][17] ),
    .A3(\registers[7][17] ),
    .S0(_1865_),
    .S1(_1885_),
    .X(_1953_));
 sky130_fd_sc_hd__mux4_1 _2610_ (.A0(\registers[0][17] ),
    .A1(\registers[2][17] ),
    .A2(\registers[4][17] ),
    .A3(\registers[6][17] ),
    .S0(_1848_),
    .S1(_1867_),
    .X(_1954_));
 sky130_fd_sc_hd__mux2i_1 _2611_ (.A0(_1953_),
    .A1(_1954_),
    .S(_1938_),
    .Y(_1955_));
 sky130_fd_sc_hd__a221o_2 _2612_ (.A1(_1785_),
    .A2(_1952_),
    .B1(_1955_),
    .B2(_1923_),
    .C1(_1798_),
    .X(_1956_));
 sky130_fd_sc_hd__a31oi_2 _2613_ (.A1(_1746_),
    .A2(_1946_),
    .A3(_1949_),
    .B1(_1956_),
    .Y(_0074_));
 sky130_fd_sc_hd__mux4_1 _2614_ (.A0(\registers[17][18] ),
    .A1(\registers[19][18] ),
    .A2(\registers[21][18] ),
    .A3(\registers[23][18] ),
    .S0(_1801_),
    .S1(_1871_),
    .X(_1957_));
 sky130_fd_sc_hd__mux2i_1 _2615_ (.A0(\registers[18][18] ),
    .A1(\registers[22][18] ),
    .S(_1829_),
    .Y(_1958_));
 sky130_fd_sc_hd__mux2i_1 _2616_ (.A0(\registers[16][18] ),
    .A1(\registers[20][18] ),
    .S(_1943_),
    .Y(_1959_));
 sky130_fd_sc_hd__a221oi_1 _2617_ (.A1(_1828_),
    .A2(_1958_),
    .B1(_1959_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_1960_));
 sky130_fd_sc_hd__o21ai_0 _2618_ (.A1(_1800_),
    .A2(_1957_),
    .B1(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__buf_8 _2619_ (.A(_1753_),
    .X(_1962_));
 sky130_fd_sc_hd__mux4_1 _2620_ (.A0(\registers[24][18] ),
    .A1(\registers[26][18] ),
    .A2(\registers[28][18] ),
    .A3(\registers[30][18] ),
    .S0(_1962_),
    .S1(_1877_),
    .X(_1963_));
 sky130_fd_sc_hd__mux4_1 _2621_ (.A0(\registers[25][18] ),
    .A1(\registers[27][18] ),
    .A2(\registers[29][18] ),
    .A3(\registers[31][18] ),
    .S0(_1839_),
    .S1(_1879_),
    .X(_1964_));
 sky130_fd_sc_hd__a22oi_4 _2622_ (.A1(_1836_),
    .A2(_1963_),
    .B1(_1964_),
    .B2(_1812_),
    .Y(_1965_));
 sky130_fd_sc_hd__mux4_1 _2623_ (.A0(\registers[0][18] ),
    .A1(\registers[1][18] ),
    .A2(\registers[2][18] ),
    .A3(\registers[3][18] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_1966_));
 sky130_fd_sc_hd__mux4_1 _2624_ (.A0(\registers[4][18] ),
    .A1(\registers[5][18] ),
    .A2(\registers[6][18] ),
    .A3(\registers[7][18] ),
    .S0(_1862_),
    .S1(_1816_),
    .X(_1967_));
 sky130_fd_sc_hd__mux2i_1 _2625_ (.A0(_1966_),
    .A1(_1967_),
    .S(_1845_),
    .Y(_1968_));
 sky130_fd_sc_hd__mux4_1 _2626_ (.A0(\registers[9][18] ),
    .A1(\registers[11][18] ),
    .A2(\registers[13][18] ),
    .A3(\registers[15][18] ),
    .S0(_1865_),
    .S1(_1885_),
    .X(_1969_));
 sky130_fd_sc_hd__mux4_1 _2627_ (.A0(\registers[8][18] ),
    .A1(\registers[10][18] ),
    .A2(\registers[12][18] ),
    .A3(\registers[14][18] ),
    .S0(_1848_),
    .S1(_1867_),
    .X(_1970_));
 sky130_fd_sc_hd__mux2i_4 _2628_ (.A0(_1969_),
    .A1(_1970_),
    .S(_1938_),
    .Y(_1971_));
 sky130_fd_sc_hd__a221o_1 _2629_ (.A1(_1793_),
    .A2(_1968_),
    .B1(_1971_),
    .B2(_1825_),
    .C1(_1798_),
    .X(_1972_));
 sky130_fd_sc_hd__a31oi_1 _2630_ (.A1(_1746_),
    .A2(_1961_),
    .A3(_1965_),
    .B1(_1972_),
    .Y(_0075_));
 sky130_fd_sc_hd__buf_8 _2631_ (.A(_1745_),
    .X(_1973_));
 sky130_fd_sc_hd__mux4_1 _2632_ (.A0(\registers[25][19] ),
    .A1(\registers[27][19] ),
    .A2(\registers[29][19] ),
    .A3(\registers[31][19] ),
    .S0(_1754_),
    .S1(_1757_),
    .X(_1974_));
 sky130_fd_sc_hd__mux2i_1 _2633_ (.A0(\registers[24][19] ),
    .A1(\registers[28][19] ),
    .S(_1840_),
    .Y(_1975_));
 sky130_fd_sc_hd__nand2_1 _2634_ (.A(_1766_),
    .B(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__mux2i_1 _2635_ (.A0(\registers[26][19] ),
    .A1(\registers[30][19] ),
    .S(_1760_),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _2636_ (.A(_1770_),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__o2111ai_4 _2637_ (.A1(_1751_),
    .A2(_1974_),
    .B1(_1976_),
    .C1(_1978_),
    .D1(_1773_),
    .Y(_1979_));
 sky130_fd_sc_hd__mux4_1 _2638_ (.A0(\registers[16][19] ),
    .A1(\registers[18][19] ),
    .A2(\registers[20][19] ),
    .A3(\registers[22][19] ),
    .S0(_1962_),
    .S1(_1877_),
    .X(_1980_));
 sky130_fd_sc_hd__mux4_1 _2639_ (.A0(\registers[17][19] ),
    .A1(\registers[19][19] ),
    .A2(\registers[21][19] ),
    .A3(\registers[23][19] ),
    .S0(_1839_),
    .S1(_1879_),
    .X(_1981_));
 sky130_fd_sc_hd__a22oi_1 _2640_ (.A1(_1778_),
    .A2(_1980_),
    .B1(_1981_),
    .B2(_1779_),
    .Y(_1982_));
 sky130_fd_sc_hd__mux4_1 _2641_ (.A0(\registers[8][19] ),
    .A1(\registers[9][19] ),
    .A2(\registers[10][19] ),
    .A3(\registers[11][19] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_1983_));
 sky130_fd_sc_hd__mux4_1 _2642_ (.A0(\registers[12][19] ),
    .A1(\registers[13][19] ),
    .A2(\registers[14][19] ),
    .A3(\registers[15][19] ),
    .S0(_1862_),
    .S1(_1816_),
    .X(_1984_));
 sky130_fd_sc_hd__mux2i_2 _2643_ (.A0(_1983_),
    .A1(_1984_),
    .S(_1845_),
    .Y(_1985_));
 sky130_fd_sc_hd__mux4_1 _2644_ (.A0(\registers[1][19] ),
    .A1(\registers[3][19] ),
    .A2(\registers[5][19] ),
    .A3(\registers[7][19] ),
    .S0(_1865_),
    .S1(_1885_),
    .X(_1986_));
 sky130_fd_sc_hd__mux4_1 _2645_ (.A0(\registers[0][19] ),
    .A1(\registers[2][19] ),
    .A2(\registers[4][19] ),
    .A3(\registers[6][19] ),
    .S0(_1848_),
    .S1(_1867_),
    .X(_1987_));
 sky130_fd_sc_hd__mux2i_1 _2646_ (.A0(_1986_),
    .A1(_1987_),
    .S(_1938_),
    .Y(_1988_));
 sky130_fd_sc_hd__buf_6 _2647_ (.A(_1797_),
    .X(_1989_));
 sky130_fd_sc_hd__a221o_4 _2648_ (.A1(_1785_),
    .A2(_1985_),
    .B1(_1988_),
    .B2(_1923_),
    .C1(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__a31oi_2 _2649_ (.A1(_1973_),
    .A2(_1979_),
    .A3(_1982_),
    .B1(_1990_),
    .Y(_0076_));
 sky130_fd_sc_hd__mux4_1 _2650_ (.A0(\registers[17][1] ),
    .A1(\registers[19][1] ),
    .A2(\registers[21][1] ),
    .A3(\registers[23][1] ),
    .S0(_1801_),
    .S1(_1871_),
    .X(_1991_));
 sky130_fd_sc_hd__mux2i_1 _2651_ (.A0(\registers[18][1] ),
    .A1(\registers[22][1] ),
    .S(_1829_),
    .Y(_1992_));
 sky130_fd_sc_hd__mux2i_1 _2652_ (.A0(\registers[16][1] ),
    .A1(\registers[20][1] ),
    .S(_1943_),
    .Y(_1993_));
 sky130_fd_sc_hd__a221oi_2 _2653_ (.A1(_1828_),
    .A2(_1992_),
    .B1(_1993_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_1994_));
 sky130_fd_sc_hd__o21ai_1 _2654_ (.A1(_1800_),
    .A2(_1991_),
    .B1(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__mux4_1 _2655_ (.A0(\registers[24][1] ),
    .A1(\registers[26][1] ),
    .A2(\registers[28][1] ),
    .A3(\registers[30][1] ),
    .S0(_1962_),
    .S1(_1877_),
    .X(_1996_));
 sky130_fd_sc_hd__mux4_1 _2656_ (.A0(\registers[25][1] ),
    .A1(\registers[27][1] ),
    .A2(\registers[29][1] ),
    .A3(\registers[31][1] ),
    .S0(_1839_),
    .S1(_1879_),
    .X(_1997_));
 sky130_fd_sc_hd__a22oi_4 _2657_ (.A1(_1836_),
    .A2(_1996_),
    .B1(_1997_),
    .B2(_1812_),
    .Y(_1998_));
 sky130_fd_sc_hd__mux4_1 _2658_ (.A0(\registers[8][1] ),
    .A1(\registers[9][1] ),
    .A2(\registers[10][1] ),
    .A3(\registers[11][1] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_1999_));
 sky130_fd_sc_hd__buf_6 _2659_ (.A(_1753_),
    .X(_2000_));
 sky130_fd_sc_hd__mux4_1 _2660_ (.A0(\registers[12][1] ),
    .A1(\registers[13][1] ),
    .A2(\registers[14][1] ),
    .A3(\registers[15][1] ),
    .S0(_1862_),
    .S1(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__mux2i_2 _2661_ (.A0(_1999_),
    .A1(_2001_),
    .S(_1845_),
    .Y(_2002_));
 sky130_fd_sc_hd__mux4_1 _2662_ (.A0(\registers[1][1] ),
    .A1(\registers[3][1] ),
    .A2(\registers[5][1] ),
    .A3(\registers[7][1] ),
    .S0(_1865_),
    .S1(_1885_),
    .X(_2003_));
 sky130_fd_sc_hd__mux4_1 _2663_ (.A0(\registers[0][1] ),
    .A1(\registers[2][1] ),
    .A2(\registers[4][1] ),
    .A3(\registers[6][1] ),
    .S0(_1848_),
    .S1(_1867_),
    .X(_2004_));
 sky130_fd_sc_hd__mux2i_1 _2664_ (.A0(_2003_),
    .A1(_2004_),
    .S(_1938_),
    .Y(_2005_));
 sky130_fd_sc_hd__a221o_4 _2665_ (.A1(_1785_),
    .A2(_2002_),
    .B1(_2005_),
    .B2(_1923_),
    .C1(_1989_),
    .X(_2006_));
 sky130_fd_sc_hd__a31oi_4 _2666_ (.A1(_1973_),
    .A2(_1995_),
    .A3(_1998_),
    .B1(_2006_),
    .Y(_0077_));
 sky130_fd_sc_hd__mux4_1 _2667_ (.A0(\registers[17][20] ),
    .A1(\registers[19][20] ),
    .A2(\registers[21][20] ),
    .A3(\registers[23][20] ),
    .S0(_1801_),
    .S1(_1871_),
    .X(_2007_));
 sky130_fd_sc_hd__mux2i_1 _2668_ (.A0(\registers[18][20] ),
    .A1(\registers[22][20] ),
    .S(_1829_),
    .Y(_2008_));
 sky130_fd_sc_hd__mux2i_1 _2669_ (.A0(\registers[16][20] ),
    .A1(\registers[20][20] ),
    .S(_1943_),
    .Y(_2009_));
 sky130_fd_sc_hd__a221oi_2 _2670_ (.A1(_1828_),
    .A2(_2008_),
    .B1(_2009_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_2010_));
 sky130_fd_sc_hd__o21ai_1 _2671_ (.A1(_1800_),
    .A2(_2007_),
    .B1(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__mux4_1 _2672_ (.A0(\registers[24][20] ),
    .A1(\registers[26][20] ),
    .A2(\registers[28][20] ),
    .A3(\registers[30][20] ),
    .S0(_1962_),
    .S1(_1877_),
    .X(_2012_));
 sky130_fd_sc_hd__buf_8 _2673_ (.A(_1763_),
    .X(_2013_));
 sky130_fd_sc_hd__mux4_1 _2674_ (.A0(\registers[25][20] ),
    .A1(\registers[27][20] ),
    .A2(\registers[29][20] ),
    .A3(\registers[31][20] ),
    .S0(_2013_),
    .S1(_1879_),
    .X(_2014_));
 sky130_fd_sc_hd__a22oi_4 _2675_ (.A1(_1836_),
    .A2(_2012_),
    .B1(_2014_),
    .B2(_1812_),
    .Y(_2015_));
 sky130_fd_sc_hd__mux4_1 _2676_ (.A0(\registers[0][20] ),
    .A1(\registers[1][20] ),
    .A2(\registers[2][20] ),
    .A3(\registers[3][20] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_2016_));
 sky130_fd_sc_hd__mux4_1 _2677_ (.A0(\registers[4][20] ),
    .A1(\registers[5][20] ),
    .A2(\registers[6][20] ),
    .A3(\registers[7][20] ),
    .S0(_1862_),
    .S1(_2000_),
    .X(_2017_));
 sky130_fd_sc_hd__buf_8 _2678_ (.A(_1819_),
    .X(_2018_));
 sky130_fd_sc_hd__mux2i_1 _2679_ (.A0(_2016_),
    .A1(_2017_),
    .S(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__mux4_1 _2680_ (.A0(\registers[9][20] ),
    .A1(\registers[11][20] ),
    .A2(\registers[13][20] ),
    .A3(\registers[15][20] ),
    .S0(_1865_),
    .S1(_1885_),
    .X(_2020_));
 sky130_fd_sc_hd__buf_6 _2681_ (.A(_1752_),
    .X(_2021_));
 sky130_fd_sc_hd__mux4_1 _2682_ (.A0(\registers[8][20] ),
    .A1(\registers[10][20] ),
    .A2(\registers[12][20] ),
    .A3(\registers[14][20] ),
    .S0(_2021_),
    .S1(_1867_),
    .X(_2022_));
 sky130_fd_sc_hd__mux2i_4 _2683_ (.A0(_2020_),
    .A1(_2022_),
    .S(_1938_),
    .Y(_2023_));
 sky130_fd_sc_hd__a221o_2 _2684_ (.A1(_1793_),
    .A2(_2019_),
    .B1(_2023_),
    .B2(_1825_),
    .C1(_1989_),
    .X(_2024_));
 sky130_fd_sc_hd__a31oi_4 _2685_ (.A1(_1973_),
    .A2(_2011_),
    .A3(_2015_),
    .B1(_2024_),
    .Y(_0078_));
 sky130_fd_sc_hd__mux4_1 _2686_ (.A0(\registers[17][21] ),
    .A1(\registers[19][21] ),
    .A2(\registers[21][21] ),
    .A3(\registers[23][21] ),
    .S0(_1801_),
    .S1(_1871_),
    .X(_2025_));
 sky130_fd_sc_hd__mux2i_1 _2687_ (.A0(\registers[18][21] ),
    .A1(\registers[22][21] ),
    .S(_1829_),
    .Y(_2026_));
 sky130_fd_sc_hd__mux2i_1 _2688_ (.A0(\registers[16][21] ),
    .A1(\registers[20][21] ),
    .S(_1943_),
    .Y(_2027_));
 sky130_fd_sc_hd__a221oi_2 _2689_ (.A1(_1828_),
    .A2(_2026_),
    .B1(_2027_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_2028_));
 sky130_fd_sc_hd__o21ai_1 _2690_ (.A1(_1800_),
    .A2(_2025_),
    .B1(_2028_),
    .Y(_2029_));
 sky130_fd_sc_hd__mux4_1 _2691_ (.A0(\registers[24][21] ),
    .A1(\registers[26][21] ),
    .A2(\registers[28][21] ),
    .A3(\registers[30][21] ),
    .S0(_1962_),
    .S1(_1877_),
    .X(_2030_));
 sky130_fd_sc_hd__mux4_1 _2692_ (.A0(\registers[25][21] ),
    .A1(\registers[27][21] ),
    .A2(\registers[29][21] ),
    .A3(\registers[31][21] ),
    .S0(_2013_),
    .S1(_1879_),
    .X(_2031_));
 sky130_fd_sc_hd__a22oi_4 _2693_ (.A1(_1836_),
    .A2(_2030_),
    .B1(_2031_),
    .B2(_1812_),
    .Y(_2032_));
 sky130_fd_sc_hd__mux4_1 _2694_ (.A0(\registers[0][21] ),
    .A1(\registers[1][21] ),
    .A2(\registers[2][21] ),
    .A3(\registers[3][21] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_2033_));
 sky130_fd_sc_hd__buf_6 _2695_ (.A(_1747_),
    .X(_2034_));
 sky130_fd_sc_hd__mux4_1 _2696_ (.A0(\registers[4][21] ),
    .A1(\registers[5][21] ),
    .A2(\registers[6][21] ),
    .A3(\registers[7][21] ),
    .S0(_2034_),
    .S1(_2000_),
    .X(_2035_));
 sky130_fd_sc_hd__mux2i_2 _2697_ (.A0(_2033_),
    .A1(_2035_),
    .S(_2018_),
    .Y(_2036_));
 sky130_fd_sc_hd__buf_6 _2698_ (.A(_1752_),
    .X(_2037_));
 sky130_fd_sc_hd__mux4_1 _2699_ (.A0(\registers[9][21] ),
    .A1(\registers[11][21] ),
    .A2(\registers[13][21] ),
    .A3(\registers[15][21] ),
    .S0(_2037_),
    .S1(_1885_),
    .X(_2038_));
 sky130_fd_sc_hd__buf_4 _2700_ (.A(_1755_),
    .X(_2039_));
 sky130_fd_sc_hd__mux4_1 _2701_ (.A0(\registers[8][21] ),
    .A1(\registers[10][21] ),
    .A2(\registers[12][21] ),
    .A3(\registers[14][21] ),
    .S0(_2021_),
    .S1(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__mux2i_4 _2702_ (.A0(_2038_),
    .A1(_2040_),
    .S(_1938_),
    .Y(_2041_));
 sky130_fd_sc_hd__a221o_4 _2703_ (.A1(_1793_),
    .A2(_2036_),
    .B1(_2041_),
    .B2(_1825_),
    .C1(_1989_),
    .X(_2042_));
 sky130_fd_sc_hd__a31oi_4 _2704_ (.A1(_1973_),
    .A2(_2029_),
    .A3(_2032_),
    .B1(_2042_),
    .Y(_0079_));
 sky130_fd_sc_hd__mux4_1 _2705_ (.A0(\registers[25][22] ),
    .A1(\registers[27][22] ),
    .A2(\registers[29][22] ),
    .A3(\registers[31][22] ),
    .S0(_1754_),
    .S1(_1757_),
    .X(_2043_));
 sky130_fd_sc_hd__mux2i_1 _2706_ (.A0(\registers[24][22] ),
    .A1(\registers[28][22] ),
    .S(_1840_),
    .Y(_2044_));
 sky130_fd_sc_hd__nand2_1 _2707_ (.A(_1766_),
    .B(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__mux2i_1 _2708_ (.A0(\registers[26][22] ),
    .A1(\registers[30][22] ),
    .S(_1760_),
    .Y(_2046_));
 sky130_fd_sc_hd__nand2_1 _2709_ (.A(_1770_),
    .B(_2046_),
    .Y(_2047_));
 sky130_fd_sc_hd__o2111ai_4 _2710_ (.A1(_1751_),
    .A2(_2043_),
    .B1(_2045_),
    .C1(_2047_),
    .D1(_1773_),
    .Y(_2048_));
 sky130_fd_sc_hd__buf_6 _2711_ (.A(_1819_),
    .X(_2049_));
 sky130_fd_sc_hd__mux4_1 _2712_ (.A0(\registers[16][22] ),
    .A1(\registers[18][22] ),
    .A2(\registers[20][22] ),
    .A3(\registers[22][22] ),
    .S0(_1962_),
    .S1(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__buf_6 _2713_ (.A(_1759_),
    .X(_2051_));
 sky130_fd_sc_hd__mux4_1 _2714_ (.A0(\registers[17][22] ),
    .A1(\registers[19][22] ),
    .A2(\registers[21][22] ),
    .A3(\registers[23][22] ),
    .S0(_2013_),
    .S1(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__a22oi_1 _2715_ (.A1(_1778_),
    .A2(_2050_),
    .B1(_2052_),
    .B2(_1779_),
    .Y(_2053_));
 sky130_fd_sc_hd__buf_6 _2716_ (.A(_1792_),
    .X(_2054_));
 sky130_fd_sc_hd__mux4_1 _2717_ (.A0(\registers[0][22] ),
    .A1(\registers[1][22] ),
    .A2(\registers[2][22] ),
    .A3(\registers[3][22] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_2055_));
 sky130_fd_sc_hd__mux4_1 _2718_ (.A0(\registers[4][22] ),
    .A1(\registers[5][22] ),
    .A2(\registers[6][22] ),
    .A3(\registers[7][22] ),
    .S0(_2034_),
    .S1(_2000_),
    .X(_2056_));
 sky130_fd_sc_hd__mux2i_1 _2719_ (.A0(_2055_),
    .A1(_2056_),
    .S(_2018_),
    .Y(_2057_));
 sky130_fd_sc_hd__buf_6 _2720_ (.A(_1756_),
    .X(_2058_));
 sky130_fd_sc_hd__mux4_1 _2721_ (.A0(\registers[9][22] ),
    .A1(\registers[11][22] ),
    .A2(\registers[13][22] ),
    .A3(\registers[15][22] ),
    .S0(_2037_),
    .S1(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__mux4_1 _2722_ (.A0(\registers[8][22] ),
    .A1(\registers[10][22] ),
    .A2(\registers[12][22] ),
    .A3(\registers[14][22] ),
    .S0(_2021_),
    .S1(_2039_),
    .X(_2060_));
 sky130_fd_sc_hd__mux2i_2 _2723_ (.A0(_2059_),
    .A1(_2060_),
    .S(_1938_),
    .Y(_2061_));
 sky130_fd_sc_hd__buf_6 _2724_ (.A(_1784_),
    .X(_2062_));
 sky130_fd_sc_hd__a221o_4 _2725_ (.A1(_2054_),
    .A2(_2057_),
    .B1(_2061_),
    .B2(_2062_),
    .C1(_1989_),
    .X(_2063_));
 sky130_fd_sc_hd__a31oi_2 _2726_ (.A1(_1973_),
    .A2(_2048_),
    .A3(_2053_),
    .B1(_2063_),
    .Y(_0080_));
 sky130_fd_sc_hd__buf_4 _2727_ (.A(_1748_),
    .X(_2064_));
 sky130_fd_sc_hd__buf_4 _2728_ (.A(_1763_),
    .X(_2065_));
 sky130_fd_sc_hd__mux4_1 _2729_ (.A0(\registers[17][23] ),
    .A1(\registers[19][23] ),
    .A2(\registers[21][23] ),
    .A3(\registers[23][23] ),
    .S0(_2065_),
    .S1(_1871_),
    .X(_2066_));
 sky130_fd_sc_hd__mux2i_2 _2730_ (.A0(\registers[18][23] ),
    .A1(\registers[22][23] ),
    .S(_1829_),
    .Y(_2067_));
 sky130_fd_sc_hd__mux2i_2 _2731_ (.A0(\registers[16][23] ),
    .A1(\registers[20][23] ),
    .S(_1943_),
    .Y(_2068_));
 sky130_fd_sc_hd__a221oi_4 _2732_ (.A1(_1828_),
    .A2(_2067_),
    .B1(_2068_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_2069_));
 sky130_fd_sc_hd__o21ai_1 _2733_ (.A1(_2064_),
    .A2(_2066_),
    .B1(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__mux4_1 _2734_ (.A0(\registers[24][23] ),
    .A1(\registers[26][23] ),
    .A2(\registers[28][23] ),
    .A3(\registers[30][23] ),
    .S0(_1962_),
    .S1(_2049_),
    .X(_2071_));
 sky130_fd_sc_hd__mux4_1 _2735_ (.A0(\registers[25][23] ),
    .A1(\registers[27][23] ),
    .A2(\registers[29][23] ),
    .A3(\registers[31][23] ),
    .S0(_2013_),
    .S1(_2051_),
    .X(_2072_));
 sky130_fd_sc_hd__buf_8 _2736_ (.A(_1811_),
    .X(_2073_));
 sky130_fd_sc_hd__a22oi_4 _2737_ (.A1(_1836_),
    .A2(_2071_),
    .B1(_2072_),
    .B2(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__buf_6 _2738_ (.A(_1747_),
    .X(_2075_));
 sky130_fd_sc_hd__buf_6 _2739_ (.A(_1763_),
    .X(_2076_));
 sky130_fd_sc_hd__mux4_1 _2740_ (.A0(\registers[0][23] ),
    .A1(\registers[1][23] ),
    .A2(\registers[2][23] ),
    .A3(\registers[3][23] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__mux4_1 _2741_ (.A0(\registers[4][23] ),
    .A1(\registers[5][23] ),
    .A2(\registers[6][23] ),
    .A3(\registers[7][23] ),
    .S0(_2034_),
    .S1(_2000_),
    .X(_2078_));
 sky130_fd_sc_hd__mux2i_1 _2742_ (.A0(_2077_),
    .A1(_2078_),
    .S(_2018_),
    .Y(_2079_));
 sky130_fd_sc_hd__mux4_1 _2743_ (.A0(\registers[9][23] ),
    .A1(\registers[11][23] ),
    .A2(\registers[13][23] ),
    .A3(\registers[15][23] ),
    .S0(_2037_),
    .S1(_2058_),
    .X(_2080_));
 sky130_fd_sc_hd__mux4_1 _2744_ (.A0(\registers[8][23] ),
    .A1(\registers[10][23] ),
    .A2(\registers[12][23] ),
    .A3(\registers[14][23] ),
    .S0(_2021_),
    .S1(_2039_),
    .X(_2081_));
 sky130_fd_sc_hd__mux2i_2 _2745_ (.A0(_2080_),
    .A1(_2081_),
    .S(_1938_),
    .Y(_2082_));
 sky130_fd_sc_hd__a221o_4 _2746_ (.A1(_2054_),
    .A2(_2079_),
    .B1(_2082_),
    .B2(_2062_),
    .C1(_1989_),
    .X(_2083_));
 sky130_fd_sc_hd__a31oi_4 _2747_ (.A1(_1973_),
    .A2(_2070_),
    .A3(_2074_),
    .B1(_2083_),
    .Y(_0081_));
 sky130_fd_sc_hd__mux4_1 _2748_ (.A0(\registers[25][24] ),
    .A1(\registers[27][24] ),
    .A2(\registers[29][24] ),
    .A3(\registers[31][24] ),
    .S0(_1754_),
    .S1(_1757_),
    .X(_2084_));
 sky130_fd_sc_hd__mux2i_1 _2749_ (.A0(\registers[24][24] ),
    .A1(\registers[28][24] ),
    .S(_1840_),
    .Y(_2085_));
 sky130_fd_sc_hd__nand2_1 _2750_ (.A(_1766_),
    .B(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__mux2i_1 _2751_ (.A0(\registers[26][24] ),
    .A1(\registers[30][24] ),
    .S(_1760_),
    .Y(_2087_));
 sky130_fd_sc_hd__nand2_1 _2752_ (.A(_1770_),
    .B(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__o2111ai_4 _2753_ (.A1(_1751_),
    .A2(_2084_),
    .B1(_2086_),
    .C1(_2088_),
    .D1(_1773_),
    .Y(_2089_));
 sky130_fd_sc_hd__mux4_2 _2754_ (.A0(\registers[16][24] ),
    .A1(\registers[18][24] ),
    .A2(\registers[20][24] ),
    .A3(\registers[22][24] ),
    .S0(_1962_),
    .S1(_2049_),
    .X(_2090_));
 sky130_fd_sc_hd__mux4_1 _2755_ (.A0(\registers[17][24] ),
    .A1(\registers[19][24] ),
    .A2(\registers[21][24] ),
    .A3(\registers[23][24] ),
    .S0(_2013_),
    .S1(_2051_),
    .X(_2091_));
 sky130_fd_sc_hd__a22oi_2 _2756_ (.A1(_1778_),
    .A2(_2090_),
    .B1(_2091_),
    .B2(_1779_),
    .Y(_2092_));
 sky130_fd_sc_hd__mux4_1 _2757_ (.A0(\registers[0][24] ),
    .A1(\registers[1][24] ),
    .A2(\registers[2][24] ),
    .A3(\registers[3][24] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2093_));
 sky130_fd_sc_hd__mux4_1 _2758_ (.A0(\registers[4][24] ),
    .A1(\registers[5][24] ),
    .A2(\registers[6][24] ),
    .A3(\registers[7][24] ),
    .S0(_2034_),
    .S1(_2000_),
    .X(_2094_));
 sky130_fd_sc_hd__mux2i_1 _2759_ (.A0(_2093_),
    .A1(_2094_),
    .S(_2018_),
    .Y(_2095_));
 sky130_fd_sc_hd__mux4_1 _2760_ (.A0(\registers[9][24] ),
    .A1(\registers[11][24] ),
    .A2(\registers[13][24] ),
    .A3(\registers[15][24] ),
    .S0(_2037_),
    .S1(_2058_),
    .X(_2096_));
 sky130_fd_sc_hd__mux4_1 _2761_ (.A0(\registers[8][24] ),
    .A1(\registers[10][24] ),
    .A2(\registers[12][24] ),
    .A3(\registers[14][24] ),
    .S0(_2021_),
    .S1(_2039_),
    .X(_2097_));
 sky130_fd_sc_hd__mux2i_4 _2762_ (.A0(_2096_),
    .A1(_2097_),
    .S(_1938_),
    .Y(_2098_));
 sky130_fd_sc_hd__a221o_4 _2763_ (.A1(_2054_),
    .A2(_2095_),
    .B1(_2098_),
    .B2(_2062_),
    .C1(_1989_),
    .X(_2099_));
 sky130_fd_sc_hd__a31oi_4 _2764_ (.A1(_1973_),
    .A2(_2089_),
    .A3(_2092_),
    .B1(_2099_),
    .Y(_0082_));
 sky130_fd_sc_hd__mux4_1 _2765_ (.A0(\registers[17][25] ),
    .A1(\registers[19][25] ),
    .A2(\registers[21][25] ),
    .A3(\registers[23][25] ),
    .S0(_2065_),
    .S1(_1871_),
    .X(_2100_));
 sky130_fd_sc_hd__buf_4 _2766_ (.A(_1769_),
    .X(_2101_));
 sky130_fd_sc_hd__buf_6 _2767_ (.A(_1756_),
    .X(_2102_));
 sky130_fd_sc_hd__mux2i_1 _2768_ (.A0(\registers[18][25] ),
    .A1(\registers[22][25] ),
    .S(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__mux2i_1 _2769_ (.A0(\registers[16][25] ),
    .A1(\registers[20][25] ),
    .S(_1943_),
    .Y(_2104_));
 sky130_fd_sc_hd__buf_6 _2770_ (.A(_1765_),
    .X(_2105_));
 sky130_fd_sc_hd__buf_4 _2771_ (.A(_1772_),
    .X(_2106_));
 sky130_fd_sc_hd__a221oi_2 _2772_ (.A1(_2101_),
    .A2(_2103_),
    .B1(_2104_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__o21ai_1 _2773_ (.A1(_2064_),
    .A2(_2100_),
    .B1(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__buf_8 _2774_ (.A(_1809_),
    .X(_2109_));
 sky130_fd_sc_hd__mux4_1 _2775_ (.A0(\registers[24][25] ),
    .A1(\registers[26][25] ),
    .A2(\registers[28][25] ),
    .A3(\registers[30][25] ),
    .S0(_1962_),
    .S1(_2049_),
    .X(_2110_));
 sky130_fd_sc_hd__mux4_1 _2776_ (.A0(\registers[25][25] ),
    .A1(\registers[27][25] ),
    .A2(\registers[29][25] ),
    .A3(\registers[31][25] ),
    .S0(_2013_),
    .S1(_2051_),
    .X(_2111_));
 sky130_fd_sc_hd__a22oi_4 _2777_ (.A1(_2109_),
    .A2(_2110_),
    .B1(_2111_),
    .B2(_2073_),
    .Y(_2112_));
 sky130_fd_sc_hd__mux4_1 _2778_ (.A0(\registers[8][25] ),
    .A1(\registers[9][25] ),
    .A2(\registers[10][25] ),
    .A3(\registers[11][25] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2113_));
 sky130_fd_sc_hd__mux4_1 _2779_ (.A0(\registers[12][25] ),
    .A1(\registers[13][25] ),
    .A2(\registers[14][25] ),
    .A3(\registers[15][25] ),
    .S0(_2034_),
    .S1(_2000_),
    .X(_2114_));
 sky130_fd_sc_hd__mux2i_2 _2780_ (.A0(_2113_),
    .A1(_2114_),
    .S(_2018_),
    .Y(_2115_));
 sky130_fd_sc_hd__mux4_1 _2781_ (.A0(\registers[1][25] ),
    .A1(\registers[3][25] ),
    .A2(\registers[5][25] ),
    .A3(\registers[7][25] ),
    .S0(_2037_),
    .S1(_2058_),
    .X(_2116_));
 sky130_fd_sc_hd__mux4_1 _2782_ (.A0(\registers[0][25] ),
    .A1(\registers[2][25] ),
    .A2(\registers[4][25] ),
    .A3(\registers[6][25] ),
    .S0(_2021_),
    .S1(_2039_),
    .X(_2117_));
 sky130_fd_sc_hd__buf_8 _2783_ (.A(_1749_),
    .X(_2118_));
 sky130_fd_sc_hd__mux2i_1 _2784_ (.A0(_2116_),
    .A1(_2117_),
    .S(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__a221o_4 _2785_ (.A1(_1785_),
    .A2(_2115_),
    .B1(_2119_),
    .B2(_1923_),
    .C1(_1989_),
    .X(_2120_));
 sky130_fd_sc_hd__a31oi_4 _2786_ (.A1(_1973_),
    .A2(_2108_),
    .A3(_2112_),
    .B1(_2120_),
    .Y(_0083_));
 sky130_fd_sc_hd__buf_4 _2787_ (.A(_1759_),
    .X(_2121_));
 sky130_fd_sc_hd__mux4_1 _2788_ (.A0(\registers[17][26] ),
    .A1(\registers[19][26] ),
    .A2(\registers[21][26] ),
    .A3(\registers[23][26] ),
    .S0(_2065_),
    .S1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__mux2i_1 _2789_ (.A0(\registers[18][26] ),
    .A1(\registers[22][26] ),
    .S(_2102_),
    .Y(_2123_));
 sky130_fd_sc_hd__mux2i_1 _2790_ (.A0(\registers[16][26] ),
    .A1(\registers[20][26] ),
    .S(_1943_),
    .Y(_2124_));
 sky130_fd_sc_hd__a221oi_2 _2791_ (.A1(_2101_),
    .A2(_2123_),
    .B1(_2124_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2125_));
 sky130_fd_sc_hd__o21ai_1 _2792_ (.A1(_2064_),
    .A2(_2122_),
    .B1(_2125_),
    .Y(_2126_));
 sky130_fd_sc_hd__mux4_1 _2793_ (.A0(\registers[24][26] ),
    .A1(\registers[26][26] ),
    .A2(\registers[28][26] ),
    .A3(\registers[30][26] ),
    .S0(_1962_),
    .S1(_2049_),
    .X(_2127_));
 sky130_fd_sc_hd__mux4_1 _2794_ (.A0(\registers[25][26] ),
    .A1(\registers[27][26] ),
    .A2(\registers[29][26] ),
    .A3(\registers[31][26] ),
    .S0(_2013_),
    .S1(_2051_),
    .X(_2128_));
 sky130_fd_sc_hd__a22oi_4 _2795_ (.A1(_2109_),
    .A2(_2127_),
    .B1(_2128_),
    .B2(_2073_),
    .Y(_2129_));
 sky130_fd_sc_hd__mux4_1 _2796_ (.A0(\registers[0][26] ),
    .A1(\registers[1][26] ),
    .A2(\registers[2][26] ),
    .A3(\registers[3][26] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2130_));
 sky130_fd_sc_hd__mux4_1 _2797_ (.A0(\registers[4][26] ),
    .A1(\registers[5][26] ),
    .A2(\registers[6][26] ),
    .A3(\registers[7][26] ),
    .S0(_2034_),
    .S1(_2000_),
    .X(_2131_));
 sky130_fd_sc_hd__mux2i_1 _2798_ (.A0(_2130_),
    .A1(_2131_),
    .S(_2018_),
    .Y(_2132_));
 sky130_fd_sc_hd__mux4_1 _2799_ (.A0(\registers[9][26] ),
    .A1(\registers[11][26] ),
    .A2(\registers[13][26] ),
    .A3(\registers[15][26] ),
    .S0(_2037_),
    .S1(_2058_),
    .X(_2133_));
 sky130_fd_sc_hd__mux4_1 _2800_ (.A0(\registers[8][26] ),
    .A1(\registers[10][26] ),
    .A2(\registers[12][26] ),
    .A3(\registers[14][26] ),
    .S0(_2021_),
    .S1(_2039_),
    .X(_2134_));
 sky130_fd_sc_hd__mux2i_4 _2801_ (.A0(_2133_),
    .A1(_2134_),
    .S(_2118_),
    .Y(_2135_));
 sky130_fd_sc_hd__a221o_2 _2802_ (.A1(_2054_),
    .A2(_2132_),
    .B1(_2135_),
    .B2(_2062_),
    .C1(_1989_),
    .X(_2136_));
 sky130_fd_sc_hd__a31oi_4 _2803_ (.A1(_1973_),
    .A2(_2126_),
    .A3(_2129_),
    .B1(_2136_),
    .Y(_0084_));
 sky130_fd_sc_hd__mux4_1 _2804_ (.A0(\registers[17][27] ),
    .A1(\registers[19][27] ),
    .A2(\registers[21][27] ),
    .A3(\registers[23][27] ),
    .S0(_2065_),
    .S1(_2121_),
    .X(_2137_));
 sky130_fd_sc_hd__mux2i_1 _2805_ (.A0(\registers[18][27] ),
    .A1(\registers[22][27] ),
    .S(_2102_),
    .Y(_2138_));
 sky130_fd_sc_hd__mux2i_1 _2806_ (.A0(\registers[16][27] ),
    .A1(\registers[20][27] ),
    .S(_1943_),
    .Y(_2139_));
 sky130_fd_sc_hd__a221oi_2 _2807_ (.A1(_2101_),
    .A2(_2138_),
    .B1(_2139_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2140_));
 sky130_fd_sc_hd__o21ai_1 _2808_ (.A1(_2064_),
    .A2(_2137_),
    .B1(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__buf_6 _2809_ (.A(_1753_),
    .X(_2142_));
 sky130_fd_sc_hd__mux4_1 _2810_ (.A0(\registers[24][27] ),
    .A1(\registers[26][27] ),
    .A2(\registers[28][27] ),
    .A3(\registers[30][27] ),
    .S0(_2142_),
    .S1(_2049_),
    .X(_2143_));
 sky130_fd_sc_hd__mux4_1 _2811_ (.A0(\registers[25][27] ),
    .A1(\registers[27][27] ),
    .A2(\registers[29][27] ),
    .A3(\registers[31][27] ),
    .S0(_2013_),
    .S1(_2051_),
    .X(_2144_));
 sky130_fd_sc_hd__a22oi_4 _2812_ (.A1(_2109_),
    .A2(_2143_),
    .B1(_2144_),
    .B2(_2073_),
    .Y(_2145_));
 sky130_fd_sc_hd__mux4_1 _2813_ (.A0(\registers[8][27] ),
    .A1(\registers[9][27] ),
    .A2(\registers[10][27] ),
    .A3(\registers[11][27] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2146_));
 sky130_fd_sc_hd__mux4_1 _2814_ (.A0(\registers[12][27] ),
    .A1(\registers[13][27] ),
    .A2(\registers[14][27] ),
    .A3(\registers[15][27] ),
    .S0(_2034_),
    .S1(_2000_),
    .X(_2147_));
 sky130_fd_sc_hd__mux2i_2 _2815_ (.A0(_2146_),
    .A1(_2147_),
    .S(_2018_),
    .Y(_2148_));
 sky130_fd_sc_hd__mux4_1 _2816_ (.A0(\registers[1][27] ),
    .A1(\registers[3][27] ),
    .A2(\registers[5][27] ),
    .A3(\registers[7][27] ),
    .S0(_2037_),
    .S1(_2058_),
    .X(_2149_));
 sky130_fd_sc_hd__mux4_1 _2817_ (.A0(\registers[0][27] ),
    .A1(\registers[2][27] ),
    .A2(\registers[4][27] ),
    .A3(\registers[6][27] ),
    .S0(_2021_),
    .S1(_2039_),
    .X(_2150_));
 sky130_fd_sc_hd__mux2i_1 _2818_ (.A0(_2149_),
    .A1(_2150_),
    .S(_2118_),
    .Y(_2151_));
 sky130_fd_sc_hd__a221o_4 _2819_ (.A1(_1785_),
    .A2(_2148_),
    .B1(_2151_),
    .B2(_1923_),
    .C1(_1989_),
    .X(_2152_));
 sky130_fd_sc_hd__a31oi_4 _2820_ (.A1(_1973_),
    .A2(_2141_),
    .A3(_2145_),
    .B1(_2152_),
    .Y(_0085_));
 sky130_fd_sc_hd__buf_4 _2821_ (.A(_1745_),
    .X(_2153_));
 sky130_fd_sc_hd__mux4_1 _2822_ (.A0(\registers[17][28] ),
    .A1(\registers[19][28] ),
    .A2(\registers[21][28] ),
    .A3(\registers[23][28] ),
    .S0(_2065_),
    .S1(_2121_),
    .X(_2154_));
 sky130_fd_sc_hd__mux2i_1 _2823_ (.A0(\registers[18][28] ),
    .A1(\registers[22][28] ),
    .S(_2102_),
    .Y(_2155_));
 sky130_fd_sc_hd__mux2i_1 _2824_ (.A0(\registers[16][28] ),
    .A1(\registers[20][28] ),
    .S(_1943_),
    .Y(_2156_));
 sky130_fd_sc_hd__a221oi_1 _2825_ (.A1(_2101_),
    .A2(_2155_),
    .B1(_2156_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2157_));
 sky130_fd_sc_hd__o21ai_0 _2826_ (.A1(_2064_),
    .A2(_2154_),
    .B1(_2157_),
    .Y(_2158_));
 sky130_fd_sc_hd__mux4_1 _2827_ (.A0(\registers[24][28] ),
    .A1(\registers[26][28] ),
    .A2(\registers[28][28] ),
    .A3(\registers[30][28] ),
    .S0(_2142_),
    .S1(_2049_),
    .X(_2159_));
 sky130_fd_sc_hd__mux4_1 _2828_ (.A0(\registers[25][28] ),
    .A1(\registers[27][28] ),
    .A2(\registers[29][28] ),
    .A3(\registers[31][28] ),
    .S0(_2013_),
    .S1(_2051_),
    .X(_2160_));
 sky130_fd_sc_hd__a22oi_4 _2829_ (.A1(_2109_),
    .A2(_2159_),
    .B1(_2160_),
    .B2(_2073_),
    .Y(_2161_));
 sky130_fd_sc_hd__mux4_1 _2830_ (.A0(\registers[0][28] ),
    .A1(\registers[1][28] ),
    .A2(\registers[2][28] ),
    .A3(\registers[3][28] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2162_));
 sky130_fd_sc_hd__mux4_1 _2831_ (.A0(\registers[4][28] ),
    .A1(\registers[5][28] ),
    .A2(\registers[6][28] ),
    .A3(\registers[7][28] ),
    .S0(_2034_),
    .S1(_2000_),
    .X(_2163_));
 sky130_fd_sc_hd__mux2i_1 _2832_ (.A0(_2162_),
    .A1(_2163_),
    .S(_2018_),
    .Y(_2164_));
 sky130_fd_sc_hd__mux4_1 _2833_ (.A0(\registers[9][28] ),
    .A1(\registers[11][28] ),
    .A2(\registers[13][28] ),
    .A3(\registers[15][28] ),
    .S0(_2037_),
    .S1(_2058_),
    .X(_2165_));
 sky130_fd_sc_hd__mux4_1 _2834_ (.A0(\registers[8][28] ),
    .A1(\registers[10][28] ),
    .A2(\registers[12][28] ),
    .A3(\registers[14][28] ),
    .S0(_2021_),
    .S1(_2039_),
    .X(_2166_));
 sky130_fd_sc_hd__mux2i_2 _2835_ (.A0(_2165_),
    .A1(_2166_),
    .S(_2118_),
    .Y(_2167_));
 sky130_fd_sc_hd__buf_4 _2836_ (.A(_1797_),
    .X(_2168_));
 sky130_fd_sc_hd__a221o_2 _2837_ (.A1(_2054_),
    .A2(_2164_),
    .B1(_2167_),
    .B2(_2062_),
    .C1(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__a31oi_2 _2838_ (.A1(_2153_),
    .A2(_2158_),
    .A3(_2161_),
    .B1(_2169_),
    .Y(_0086_));
 sky130_fd_sc_hd__mux4_1 _2839_ (.A0(\registers[25][29] ),
    .A1(\registers[27][29] ),
    .A2(\registers[29][29] ),
    .A3(\registers[31][29] ),
    .S0(_1754_),
    .S1(_1757_),
    .X(_2170_));
 sky130_fd_sc_hd__mux2i_1 _2840_ (.A0(\registers[24][29] ),
    .A1(\registers[28][29] ),
    .S(_1840_),
    .Y(_2171_));
 sky130_fd_sc_hd__nand2_1 _2841_ (.A(_1766_),
    .B(_2171_),
    .Y(_2172_));
 sky130_fd_sc_hd__mux2i_1 _2842_ (.A0(\registers[26][29] ),
    .A1(\registers[30][29] ),
    .S(_1760_),
    .Y(_2173_));
 sky130_fd_sc_hd__nand2_1 _2843_ (.A(_1770_),
    .B(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__o2111ai_4 _2844_ (.A1(_1751_),
    .A2(_2170_),
    .B1(_2172_),
    .C1(_2174_),
    .D1(_1773_),
    .Y(_2175_));
 sky130_fd_sc_hd__mux4_1 _2845_ (.A0(\registers[16][29] ),
    .A1(\registers[18][29] ),
    .A2(\registers[20][29] ),
    .A3(\registers[22][29] ),
    .S0(_2142_),
    .S1(_2049_),
    .X(_2176_));
 sky130_fd_sc_hd__mux4_1 _2846_ (.A0(\registers[17][29] ),
    .A1(\registers[19][29] ),
    .A2(\registers[21][29] ),
    .A3(\registers[23][29] ),
    .S0(_2013_),
    .S1(_2051_),
    .X(_2177_));
 sky130_fd_sc_hd__a22oi_1 _2847_ (.A1(_1778_),
    .A2(_2176_),
    .B1(_2177_),
    .B2(_1779_),
    .Y(_2178_));
 sky130_fd_sc_hd__mux4_1 _2848_ (.A0(\registers[8][29] ),
    .A1(\registers[9][29] ),
    .A2(\registers[10][29] ),
    .A3(\registers[11][29] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2179_));
 sky130_fd_sc_hd__buf_6 _2849_ (.A(_1753_),
    .X(_2180_));
 sky130_fd_sc_hd__mux4_1 _2850_ (.A0(\registers[12][29] ),
    .A1(\registers[13][29] ),
    .A2(\registers[14][29] ),
    .A3(\registers[15][29] ),
    .S0(_2034_),
    .S1(_2180_),
    .X(_2181_));
 sky130_fd_sc_hd__mux2i_2 _2851_ (.A0(_2179_),
    .A1(_2181_),
    .S(_2018_),
    .Y(_2182_));
 sky130_fd_sc_hd__mux4_1 _2852_ (.A0(\registers[1][29] ),
    .A1(\registers[3][29] ),
    .A2(\registers[5][29] ),
    .A3(\registers[7][29] ),
    .S0(_2037_),
    .S1(_2058_),
    .X(_2183_));
 sky130_fd_sc_hd__mux4_1 _2853_ (.A0(\registers[0][29] ),
    .A1(\registers[2][29] ),
    .A2(\registers[4][29] ),
    .A3(\registers[6][29] ),
    .S0(_2021_),
    .S1(_2039_),
    .X(_2184_));
 sky130_fd_sc_hd__mux2i_1 _2854_ (.A0(_2183_),
    .A1(_2184_),
    .S(_2118_),
    .Y(_2185_));
 sky130_fd_sc_hd__a221o_2 _2855_ (.A1(_1785_),
    .A2(_2182_),
    .B1(_2185_),
    .B2(_1923_),
    .C1(_2168_),
    .X(_2186_));
 sky130_fd_sc_hd__a31oi_2 _2856_ (.A1(_2153_),
    .A2(_2175_),
    .A3(_2178_),
    .B1(_2186_),
    .Y(_0087_));
 sky130_fd_sc_hd__mux4_1 _2857_ (.A0(\registers[17][2] ),
    .A1(\registers[19][2] ),
    .A2(\registers[21][2] ),
    .A3(\registers[23][2] ),
    .S0(_2065_),
    .S1(_2121_),
    .X(_2187_));
 sky130_fd_sc_hd__mux2i_1 _2858_ (.A0(\registers[18][2] ),
    .A1(\registers[22][2] ),
    .S(_2102_),
    .Y(_2188_));
 sky130_fd_sc_hd__mux2i_1 _2859_ (.A0(\registers[16][2] ),
    .A1(\registers[20][2] ),
    .S(_1837_),
    .Y(_2189_));
 sky130_fd_sc_hd__a221oi_1 _2860_ (.A1(_2101_),
    .A2(_2188_),
    .B1(_2189_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2190_));
 sky130_fd_sc_hd__o21ai_0 _2861_ (.A1(_2064_),
    .A2(_2187_),
    .B1(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__mux4_1 _2862_ (.A0(\registers[24][2] ),
    .A1(\registers[26][2] ),
    .A2(\registers[28][2] ),
    .A3(\registers[30][2] ),
    .S0(_2142_),
    .S1(_2049_),
    .X(_2192_));
 sky130_fd_sc_hd__buf_6 _2863_ (.A(_1763_),
    .X(_2193_));
 sky130_fd_sc_hd__mux4_1 _2864_ (.A0(\registers[25][2] ),
    .A1(\registers[27][2] ),
    .A2(\registers[29][2] ),
    .A3(\registers[31][2] ),
    .S0(_2193_),
    .S1(_2051_),
    .X(_2194_));
 sky130_fd_sc_hd__a22oi_4 _2865_ (.A1(_2109_),
    .A2(_2192_),
    .B1(_2194_),
    .B2(_2073_),
    .Y(_2195_));
 sky130_fd_sc_hd__mux4_1 _2866_ (.A0(\registers[8][2] ),
    .A1(\registers[9][2] ),
    .A2(\registers[10][2] ),
    .A3(\registers[11][2] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2196_));
 sky130_fd_sc_hd__mux4_1 _2867_ (.A0(\registers[12][2] ),
    .A1(\registers[13][2] ),
    .A2(\registers[14][2] ),
    .A3(\registers[15][2] ),
    .S0(_2034_),
    .S1(_2180_),
    .X(_2197_));
 sky130_fd_sc_hd__buf_8 _2868_ (.A(_1819_),
    .X(_2198_));
 sky130_fd_sc_hd__mux2i_2 _2869_ (.A0(_2196_),
    .A1(_2197_),
    .S(_2198_),
    .Y(_2199_));
 sky130_fd_sc_hd__mux4_1 _2870_ (.A0(\registers[1][2] ),
    .A1(\registers[3][2] ),
    .A2(\registers[5][2] ),
    .A3(\registers[7][2] ),
    .S0(_2037_),
    .S1(_2058_),
    .X(_2200_));
 sky130_fd_sc_hd__buf_8 _2871_ (.A(_1752_),
    .X(_2201_));
 sky130_fd_sc_hd__mux4_1 _2872_ (.A0(\registers[0][2] ),
    .A1(\registers[2][2] ),
    .A2(\registers[4][2] ),
    .A3(\registers[6][2] ),
    .S0(_2201_),
    .S1(_2039_),
    .X(_2202_));
 sky130_fd_sc_hd__mux2i_1 _2873_ (.A0(_2200_),
    .A1(_2202_),
    .S(_2118_),
    .Y(_2203_));
 sky130_fd_sc_hd__a221o_2 _2874_ (.A1(_1785_),
    .A2(_2199_),
    .B1(_2203_),
    .B2(_1923_),
    .C1(_2168_),
    .X(_2204_));
 sky130_fd_sc_hd__a31oi_1 _2875_ (.A1(_2153_),
    .A2(_2191_),
    .A3(_2195_),
    .B1(_2204_),
    .Y(_0088_));
 sky130_fd_sc_hd__mux4_1 _2876_ (.A0(\registers[17][30] ),
    .A1(\registers[19][30] ),
    .A2(\registers[21][30] ),
    .A3(\registers[23][30] ),
    .S0(_2065_),
    .S1(_2121_),
    .X(_2205_));
 sky130_fd_sc_hd__mux2i_2 _2877_ (.A0(\registers[18][30] ),
    .A1(\registers[22][30] ),
    .S(_2102_),
    .Y(_2206_));
 sky130_fd_sc_hd__mux2i_1 _2878_ (.A0(\registers[16][30] ),
    .A1(\registers[20][30] ),
    .S(_1837_),
    .Y(_2207_));
 sky130_fd_sc_hd__a221oi_2 _2879_ (.A1(_2101_),
    .A2(_2206_),
    .B1(_2207_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2208_));
 sky130_fd_sc_hd__o21ai_0 _2880_ (.A1(_2064_),
    .A2(_2205_),
    .B1(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__mux4_1 _2881_ (.A0(\registers[24][30] ),
    .A1(\registers[26][30] ),
    .A2(\registers[28][30] ),
    .A3(\registers[30][30] ),
    .S0(_2142_),
    .S1(_2049_),
    .X(_2210_));
 sky130_fd_sc_hd__mux4_1 _2882_ (.A0(\registers[25][30] ),
    .A1(\registers[27][30] ),
    .A2(\registers[29][30] ),
    .A3(\registers[31][30] ),
    .S0(_2193_),
    .S1(_2051_),
    .X(_2211_));
 sky130_fd_sc_hd__a22oi_2 _2883_ (.A1(_2109_),
    .A2(_2210_),
    .B1(_2211_),
    .B2(_2073_),
    .Y(_2212_));
 sky130_fd_sc_hd__mux4_1 _2884_ (.A0(\registers[0][30] ),
    .A1(\registers[1][30] ),
    .A2(\registers[2][30] ),
    .A3(\registers[3][30] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2213_));
 sky130_fd_sc_hd__mux4_1 _2885_ (.A0(\registers[4][30] ),
    .A1(\registers[5][30] ),
    .A2(\registers[6][30] ),
    .A3(\registers[7][30] ),
    .S0(_1899_),
    .S1(_2180_),
    .X(_2214_));
 sky130_fd_sc_hd__mux2i_1 _2886_ (.A0(_2213_),
    .A1(_2214_),
    .S(_2198_),
    .Y(_2215_));
 sky130_fd_sc_hd__mux4_1 _2887_ (.A0(\registers[9][30] ),
    .A1(\registers[11][30] ),
    .A2(\registers[13][30] ),
    .A3(\registers[15][30] ),
    .S0(_1821_),
    .S1(_2058_),
    .X(_2216_));
 sky130_fd_sc_hd__mux4_1 _2888_ (.A0(\registers[8][30] ),
    .A1(\registers[10][30] ),
    .A2(\registers[12][30] ),
    .A3(\registers[14][30] ),
    .S0(_2201_),
    .S1(_1789_),
    .X(_2217_));
 sky130_fd_sc_hd__mux2i_2 _2889_ (.A0(_2216_),
    .A1(_2217_),
    .S(_2118_),
    .Y(_2218_));
 sky130_fd_sc_hd__a221o_2 _2890_ (.A1(_2054_),
    .A2(_2215_),
    .B1(_2218_),
    .B2(_2062_),
    .C1(_2168_),
    .X(_2219_));
 sky130_fd_sc_hd__a31oi_1 _2891_ (.A1(_2153_),
    .A2(_2209_),
    .A3(_2212_),
    .B1(_2219_),
    .Y(_0089_));
 sky130_fd_sc_hd__mux4_1 _2892_ (.A0(\registers[17][31] ),
    .A1(\registers[19][31] ),
    .A2(\registers[21][31] ),
    .A3(\registers[23][31] ),
    .S0(_2065_),
    .S1(_2121_),
    .X(_2220_));
 sky130_fd_sc_hd__mux2i_2 _2893_ (.A0(\registers[18][31] ),
    .A1(\registers[22][31] ),
    .S(_2102_),
    .Y(_2221_));
 sky130_fd_sc_hd__mux2i_1 _2894_ (.A0(\registers[16][31] ),
    .A1(\registers[20][31] ),
    .S(_1837_),
    .Y(_2222_));
 sky130_fd_sc_hd__a221oi_2 _2895_ (.A1(_2101_),
    .A2(_2221_),
    .B1(_2222_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2223_));
 sky130_fd_sc_hd__o21ai_0 _2896_ (.A1(_2064_),
    .A2(_2220_),
    .B1(_2223_),
    .Y(_2224_));
 sky130_fd_sc_hd__mux4_1 _2897_ (.A0(\registers[24][31] ),
    .A1(\registers[26][31] ),
    .A2(\registers[28][31] ),
    .A3(\registers[30][31] ),
    .S0(_2142_),
    .S1(_1790_),
    .X(_2225_));
 sky130_fd_sc_hd__mux4_1 _2898_ (.A0(\registers[25][31] ),
    .A1(\registers[27][31] ),
    .A2(\registers[29][31] ),
    .A3(\registers[31][31] ),
    .S0(_2193_),
    .S1(_1802_),
    .X(_2226_));
 sky130_fd_sc_hd__a22oi_2 _2899_ (.A1(_2109_),
    .A2(_2225_),
    .B1(_2226_),
    .B2(_2073_),
    .Y(_2227_));
 sky130_fd_sc_hd__mux4_1 _2900_ (.A0(\registers[0][31] ),
    .A1(\registers[1][31] ),
    .A2(\registers[2][31] ),
    .A3(\registers[3][31] ),
    .S0(_2075_),
    .S1(_2076_),
    .X(_2228_));
 sky130_fd_sc_hd__mux4_1 _2901_ (.A0(\registers[4][31] ),
    .A1(\registers[5][31] ),
    .A2(\registers[6][31] ),
    .A3(\registers[7][31] ),
    .S0(_1899_),
    .S1(_2180_),
    .X(_2229_));
 sky130_fd_sc_hd__mux2i_1 _2902_ (.A0(_2228_),
    .A1(_2229_),
    .S(_2198_),
    .Y(_2230_));
 sky130_fd_sc_hd__mux4_1 _2903_ (.A0(\registers[9][31] ),
    .A1(\registers[11][31] ),
    .A2(\registers[13][31] ),
    .A3(\registers[15][31] ),
    .S0(_1821_),
    .S1(_1822_),
    .X(_2231_));
 sky130_fd_sc_hd__mux4_1 _2904_ (.A0(\registers[8][31] ),
    .A1(\registers[10][31] ),
    .A2(\registers[12][31] ),
    .A3(\registers[14][31] ),
    .S0(_2201_),
    .S1(_1789_),
    .X(_2232_));
 sky130_fd_sc_hd__mux2i_2 _2905_ (.A0(_2231_),
    .A1(_2232_),
    .S(_2118_),
    .Y(_2233_));
 sky130_fd_sc_hd__a221o_2 _2906_ (.A1(_2054_),
    .A2(_2230_),
    .B1(_2233_),
    .B2(_2062_),
    .C1(_2168_),
    .X(_2234_));
 sky130_fd_sc_hd__a31oi_1 _2907_ (.A1(_2153_),
    .A2(_2224_),
    .A3(_2227_),
    .B1(_2234_),
    .Y(_0090_));
 sky130_fd_sc_hd__mux4_1 _2908_ (.A0(\registers[25][3] ),
    .A1(\registers[27][3] ),
    .A2(\registers[29][3] ),
    .A3(\registers[31][3] ),
    .S0(_1763_),
    .S1(_1757_),
    .X(_2235_));
 sky130_fd_sc_hd__mux2i_1 _2909_ (.A0(\registers[24][3] ),
    .A1(\registers[28][3] ),
    .S(_1840_),
    .Y(_2236_));
 sky130_fd_sc_hd__nand2_1 _2910_ (.A(_1766_),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__mux2i_1 _2911_ (.A0(\registers[26][3] ),
    .A1(\registers[30][3] ),
    .S(_1760_),
    .Y(_2238_));
 sky130_fd_sc_hd__nand2_1 _2912_ (.A(_1770_),
    .B(_2238_),
    .Y(_2239_));
 sky130_fd_sc_hd__o2111ai_4 _2913_ (.A1(_1750_),
    .A2(_2235_),
    .B1(_2237_),
    .C1(_2239_),
    .D1(_1773_),
    .Y(_2240_));
 sky130_fd_sc_hd__mux4_1 _2914_ (.A0(\registers[16][3] ),
    .A1(\registers[18][3] ),
    .A2(\registers[20][3] ),
    .A3(\registers[22][3] ),
    .S0(_2142_),
    .S1(_1790_),
    .X(_2241_));
 sky130_fd_sc_hd__mux4_1 _2915_ (.A0(\registers[17][3] ),
    .A1(\registers[19][3] ),
    .A2(\registers[21][3] ),
    .A3(\registers[23][3] ),
    .S0(_2193_),
    .S1(_1802_),
    .X(_2242_));
 sky130_fd_sc_hd__a22oi_1 _2916_ (.A1(_1778_),
    .A2(_2241_),
    .B1(_2242_),
    .B2(_1779_),
    .Y(_2243_));
 sky130_fd_sc_hd__mux4_1 _2917_ (.A0(\registers[0][3] ),
    .A1(\registers[1][3] ),
    .A2(\registers[2][3] ),
    .A3(\registers[3][3] ),
    .S0(_1787_),
    .S1(_1775_),
    .X(_2244_));
 sky130_fd_sc_hd__mux4_1 _2918_ (.A0(\registers[4][3] ),
    .A1(\registers[5][3] ),
    .A2(\registers[6][3] ),
    .A3(\registers[7][3] ),
    .S0(_1899_),
    .S1(_2180_),
    .X(_2245_));
 sky130_fd_sc_hd__mux2i_1 _2919_ (.A0(_2244_),
    .A1(_2245_),
    .S(_2198_),
    .Y(_2246_));
 sky130_fd_sc_hd__mux4_1 _2920_ (.A0(\registers[9][3] ),
    .A1(\registers[11][3] ),
    .A2(\registers[13][3] ),
    .A3(\registers[15][3] ),
    .S0(_1821_),
    .S1(_1822_),
    .X(_2247_));
 sky130_fd_sc_hd__mux4_1 _2921_ (.A0(\registers[8][3] ),
    .A1(\registers[10][3] ),
    .A2(\registers[12][3] ),
    .A3(\registers[14][3] ),
    .S0(_2201_),
    .S1(_1789_),
    .X(_2248_));
 sky130_fd_sc_hd__mux2i_4 _2922_ (.A0(_2247_),
    .A1(_2248_),
    .S(_2118_),
    .Y(_2249_));
 sky130_fd_sc_hd__a221o_2 _2923_ (.A1(_2054_),
    .A2(_2246_),
    .B1(_2249_),
    .B2(_2062_),
    .C1(_2168_),
    .X(_2250_));
 sky130_fd_sc_hd__a31oi_2 _2924_ (.A1(_2153_),
    .A2(_2240_),
    .A3(_2243_),
    .B1(_2250_),
    .Y(_0091_));
 sky130_fd_sc_hd__mux4_1 _2925_ (.A0(\registers[17][4] ),
    .A1(\registers[19][4] ),
    .A2(\registers[21][4] ),
    .A3(\registers[23][4] ),
    .S0(_2065_),
    .S1(_2121_),
    .X(_2251_));
 sky130_fd_sc_hd__mux2i_1 _2926_ (.A0(\registers[18][4] ),
    .A1(\registers[22][4] ),
    .S(_2102_),
    .Y(_2252_));
 sky130_fd_sc_hd__mux2i_1 _2927_ (.A0(\registers[16][4] ),
    .A1(\registers[20][4] ),
    .S(_1837_),
    .Y(_2253_));
 sky130_fd_sc_hd__a221oi_1 _2928_ (.A1(_2101_),
    .A2(_2252_),
    .B1(_2253_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2254_));
 sky130_fd_sc_hd__o21ai_0 _2929_ (.A1(_2064_),
    .A2(_2251_),
    .B1(_2254_),
    .Y(_2255_));
 sky130_fd_sc_hd__mux4_1 _2930_ (.A0(\registers[24][4] ),
    .A1(\registers[26][4] ),
    .A2(\registers[28][4] ),
    .A3(\registers[30][4] ),
    .S0(_2142_),
    .S1(_1790_),
    .X(_2256_));
 sky130_fd_sc_hd__mux4_1 _2931_ (.A0(\registers[25][4] ),
    .A1(\registers[27][4] ),
    .A2(\registers[29][4] ),
    .A3(\registers[31][4] ),
    .S0(_2193_),
    .S1(_1802_),
    .X(_2257_));
 sky130_fd_sc_hd__a22oi_2 _2932_ (.A1(_2109_),
    .A2(_2256_),
    .B1(_2257_),
    .B2(_2073_),
    .Y(_2258_));
 sky130_fd_sc_hd__mux4_1 _2933_ (.A0(\registers[0][4] ),
    .A1(\registers[1][4] ),
    .A2(\registers[2][4] ),
    .A3(\registers[3][4] ),
    .S0(_1787_),
    .S1(_1775_),
    .X(_2259_));
 sky130_fd_sc_hd__mux4_1 _2934_ (.A0(\registers[4][4] ),
    .A1(\registers[5][4] ),
    .A2(\registers[6][4] ),
    .A3(\registers[7][4] ),
    .S0(_1899_),
    .S1(_2180_),
    .X(_2260_));
 sky130_fd_sc_hd__mux2i_1 _2935_ (.A0(_2259_),
    .A1(_2260_),
    .S(_2198_),
    .Y(_2261_));
 sky130_fd_sc_hd__mux4_1 _2936_ (.A0(\registers[9][4] ),
    .A1(\registers[11][4] ),
    .A2(\registers[13][4] ),
    .A3(\registers[15][4] ),
    .S0(_1821_),
    .S1(_1822_),
    .X(_2262_));
 sky130_fd_sc_hd__mux4_1 _2937_ (.A0(\registers[8][4] ),
    .A1(\registers[10][4] ),
    .A2(\registers[12][4] ),
    .A3(\registers[14][4] ),
    .S0(_2201_),
    .S1(_1789_),
    .X(_2263_));
 sky130_fd_sc_hd__mux2i_2 _2938_ (.A0(_2262_),
    .A1(_2263_),
    .S(_2118_),
    .Y(_2264_));
 sky130_fd_sc_hd__a221o_1 _2939_ (.A1(_2054_),
    .A2(_2261_),
    .B1(_2264_),
    .B2(_2062_),
    .C1(_2168_),
    .X(_2265_));
 sky130_fd_sc_hd__a31oi_1 _2940_ (.A1(_2153_),
    .A2(_2255_),
    .A3(_2258_),
    .B1(_2265_),
    .Y(_0092_));
 sky130_fd_sc_hd__mux4_1 _2941_ (.A0(\registers[25][5] ),
    .A1(\registers[27][5] ),
    .A2(\registers[29][5] ),
    .A3(\registers[31][5] ),
    .S0(_1763_),
    .S1(_1757_),
    .X(_2266_));
 sky130_fd_sc_hd__mux2i_1 _2942_ (.A0(\registers[24][5] ),
    .A1(\registers[28][5] ),
    .S(_1840_),
    .Y(_2267_));
 sky130_fd_sc_hd__nand2_1 _2943_ (.A(_1766_),
    .B(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__mux2i_1 _2944_ (.A0(\registers[26][5] ),
    .A1(\registers[30][5] ),
    .S(_1760_),
    .Y(_2269_));
 sky130_fd_sc_hd__nand2_1 _2945_ (.A(_1770_),
    .B(_2269_),
    .Y(_2270_));
 sky130_fd_sc_hd__o2111ai_4 _2946_ (.A1(_1750_),
    .A2(_2266_),
    .B1(_2268_),
    .C1(_2270_),
    .D1(_1773_),
    .Y(_2271_));
 sky130_fd_sc_hd__mux4_1 _2947_ (.A0(\registers[16][5] ),
    .A1(\registers[18][5] ),
    .A2(\registers[20][5] ),
    .A3(\registers[22][5] ),
    .S0(_2142_),
    .S1(_1790_),
    .X(_2272_));
 sky130_fd_sc_hd__mux4_1 _2948_ (.A0(\registers[17][5] ),
    .A1(\registers[19][5] ),
    .A2(\registers[21][5] ),
    .A3(\registers[23][5] ),
    .S0(_2193_),
    .S1(_1802_),
    .X(_2273_));
 sky130_fd_sc_hd__a22oi_1 _2949_ (.A1(_1778_),
    .A2(_2272_),
    .B1(_2273_),
    .B2(_1779_),
    .Y(_2274_));
 sky130_fd_sc_hd__mux4_1 _2950_ (.A0(\registers[0][5] ),
    .A1(\registers[1][5] ),
    .A2(\registers[2][5] ),
    .A3(\registers[3][5] ),
    .S0(_1787_),
    .S1(_1775_),
    .X(_2275_));
 sky130_fd_sc_hd__mux4_1 _2951_ (.A0(\registers[4][5] ),
    .A1(\registers[5][5] ),
    .A2(\registers[6][5] ),
    .A3(\registers[7][5] ),
    .S0(_1899_),
    .S1(_2180_),
    .X(_2276_));
 sky130_fd_sc_hd__mux2i_1 _2952_ (.A0(_2275_),
    .A1(_2276_),
    .S(_2198_),
    .Y(_2277_));
 sky130_fd_sc_hd__mux4_1 _2953_ (.A0(\registers[9][5] ),
    .A1(\registers[11][5] ),
    .A2(\registers[13][5] ),
    .A3(\registers[15][5] ),
    .S0(_1821_),
    .S1(_1822_),
    .X(_2278_));
 sky130_fd_sc_hd__mux4_1 _2954_ (.A0(\registers[8][5] ),
    .A1(\registers[10][5] ),
    .A2(\registers[12][5] ),
    .A3(\registers[14][5] ),
    .S0(_2201_),
    .S1(_1789_),
    .X(_2279_));
 sky130_fd_sc_hd__mux2i_2 _2955_ (.A0(_2278_),
    .A1(_2279_),
    .S(_1749_),
    .Y(_2280_));
 sky130_fd_sc_hd__a221o_2 _2956_ (.A1(_2054_),
    .A2(_2277_),
    .B1(_2280_),
    .B2(_2062_),
    .C1(_2168_),
    .X(_2281_));
 sky130_fd_sc_hd__a31oi_2 _2957_ (.A1(_2153_),
    .A2(_2271_),
    .A3(_2274_),
    .B1(_2281_),
    .Y(_0093_));
 sky130_fd_sc_hd__mux4_1 _2958_ (.A0(\registers[17][6] ),
    .A1(\registers[19][6] ),
    .A2(\registers[21][6] ),
    .A3(\registers[23][6] ),
    .S0(_2065_),
    .S1(_2121_),
    .X(_2282_));
 sky130_fd_sc_hd__mux2i_1 _2959_ (.A0(\registers[18][6] ),
    .A1(\registers[22][6] ),
    .S(_2102_),
    .Y(_2283_));
 sky130_fd_sc_hd__mux2i_1 _2960_ (.A0(\registers[16][6] ),
    .A1(\registers[20][6] ),
    .S(_1837_),
    .Y(_2284_));
 sky130_fd_sc_hd__a221oi_1 _2961_ (.A1(_2101_),
    .A2(_2283_),
    .B1(_2284_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2285_));
 sky130_fd_sc_hd__o21ai_0 _2962_ (.A1(_2064_),
    .A2(_2282_),
    .B1(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__mux4_1 _2963_ (.A0(\registers[24][6] ),
    .A1(\registers[26][6] ),
    .A2(\registers[28][6] ),
    .A3(\registers[30][6] ),
    .S0(_2142_),
    .S1(_1790_),
    .X(_2287_));
 sky130_fd_sc_hd__mux4_1 _2964_ (.A0(\registers[25][6] ),
    .A1(\registers[27][6] ),
    .A2(\registers[29][6] ),
    .A3(\registers[31][6] ),
    .S0(_2193_),
    .S1(_1802_),
    .X(_2288_));
 sky130_fd_sc_hd__a22oi_2 _2965_ (.A1(_2109_),
    .A2(_2287_),
    .B1(_2288_),
    .B2(_2073_),
    .Y(_2289_));
 sky130_fd_sc_hd__mux4_1 _2966_ (.A0(\registers[8][6] ),
    .A1(\registers[9][6] ),
    .A2(\registers[10][6] ),
    .A3(\registers[11][6] ),
    .S0(_1787_),
    .S1(_1775_),
    .X(_2290_));
 sky130_fd_sc_hd__mux4_1 _2967_ (.A0(\registers[12][6] ),
    .A1(\registers[13][6] ),
    .A2(\registers[14][6] ),
    .A3(\registers[15][6] ),
    .S0(_1899_),
    .S1(_2180_),
    .X(_2291_));
 sky130_fd_sc_hd__mux2i_1 _2968_ (.A0(_2290_),
    .A1(_2291_),
    .S(_2198_),
    .Y(_2292_));
 sky130_fd_sc_hd__mux4_1 _2969_ (.A0(\registers[1][6] ),
    .A1(\registers[3][6] ),
    .A2(\registers[5][6] ),
    .A3(\registers[7][6] ),
    .S0(_1821_),
    .S1(_1822_),
    .X(_2293_));
 sky130_fd_sc_hd__mux4_1 _2970_ (.A0(\registers[0][6] ),
    .A1(\registers[2][6] ),
    .A2(\registers[4][6] ),
    .A3(\registers[6][6] ),
    .S0(_2201_),
    .S1(_1789_),
    .X(_2294_));
 sky130_fd_sc_hd__mux2i_1 _2971_ (.A0(_2293_),
    .A1(_2294_),
    .S(_1749_),
    .Y(_2295_));
 sky130_fd_sc_hd__a221o_1 _2972_ (.A1(_1785_),
    .A2(_2292_),
    .B1(_2295_),
    .B2(_1792_),
    .C1(_2168_),
    .X(_2296_));
 sky130_fd_sc_hd__a31oi_1 _2973_ (.A1(_2153_),
    .A2(_2286_),
    .A3(_2289_),
    .B1(_2296_),
    .Y(_0094_));
 sky130_fd_sc_hd__mux4_1 _2974_ (.A0(\registers[17][7] ),
    .A1(\registers[19][7] ),
    .A2(\registers[21][7] ),
    .A3(\registers[23][7] ),
    .S0(_1780_),
    .S1(_2121_),
    .X(_2297_));
 sky130_fd_sc_hd__mux2i_1 _2975_ (.A0(\registers[18][7] ),
    .A1(\registers[22][7] ),
    .S(_2102_),
    .Y(_2298_));
 sky130_fd_sc_hd__mux2i_1 _2976_ (.A0(\registers[16][7] ),
    .A1(\registers[20][7] ),
    .S(_1837_),
    .Y(_2299_));
 sky130_fd_sc_hd__a221oi_1 _2977_ (.A1(_2101_),
    .A2(_2298_),
    .B1(_2299_),
    .B2(_2105_),
    .C1(_2106_),
    .Y(_2300_));
 sky130_fd_sc_hd__o21ai_1 _2978_ (.A1(_1751_),
    .A2(_2297_),
    .B1(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hd__mux4_1 _2979_ (.A0(\registers[24][7] ),
    .A1(\registers[26][7] ),
    .A2(\registers[28][7] ),
    .A3(\registers[30][7] ),
    .S0(_1754_),
    .S1(_1790_),
    .X(_2302_));
 sky130_fd_sc_hd__mux4_1 _2980_ (.A0(\registers[25][7] ),
    .A1(\registers[27][7] ),
    .A2(\registers[29][7] ),
    .A3(\registers[31][7] ),
    .S0(_2193_),
    .S1(_1802_),
    .X(_2303_));
 sky130_fd_sc_hd__a22oi_4 _2981_ (.A1(_2109_),
    .A2(_2302_),
    .B1(_2303_),
    .B2(_1811_),
    .Y(_2304_));
 sky130_fd_sc_hd__mux4_1 _2982_ (.A0(\registers[0][7] ),
    .A1(\registers[1][7] ),
    .A2(\registers[2][7] ),
    .A3(\registers[3][7] ),
    .S0(_1787_),
    .S1(_1775_),
    .X(_2305_));
 sky130_fd_sc_hd__mux4_1 _2983_ (.A0(\registers[4][7] ),
    .A1(\registers[5][7] ),
    .A2(\registers[6][7] ),
    .A3(\registers[7][7] ),
    .S0(_1899_),
    .S1(_2180_),
    .X(_2306_));
 sky130_fd_sc_hd__mux2i_1 _2984_ (.A0(_2305_),
    .A1(_2306_),
    .S(_2198_),
    .Y(_2307_));
 sky130_fd_sc_hd__mux4_1 _2985_ (.A0(\registers[9][7] ),
    .A1(\registers[11][7] ),
    .A2(\registers[13][7] ),
    .A3(\registers[15][7] ),
    .S0(_1821_),
    .S1(_1822_),
    .X(_2308_));
 sky130_fd_sc_hd__mux4_1 _2986_ (.A0(\registers[8][7] ),
    .A1(\registers[10][7] ),
    .A2(\registers[12][7] ),
    .A3(\registers[14][7] ),
    .S0(_2201_),
    .S1(_1789_),
    .X(_2309_));
 sky130_fd_sc_hd__mux2i_1 _2987_ (.A0(_2308_),
    .A1(_2309_),
    .S(_1749_),
    .Y(_2310_));
 sky130_fd_sc_hd__a221o_2 _2988_ (.A1(_1923_),
    .A2(_2307_),
    .B1(_2310_),
    .B2(_1784_),
    .C1(_2168_),
    .X(_2311_));
 sky130_fd_sc_hd__a31oi_4 _2989_ (.A1(_2153_),
    .A2(_2301_),
    .A3(_2304_),
    .B1(_2311_),
    .Y(_0095_));
 sky130_fd_sc_hd__mux4_1 _2990_ (.A0(\registers[17][8] ),
    .A1(\registers[19][8] ),
    .A2(\registers[21][8] ),
    .A3(\registers[23][8] ),
    .S0(_1780_),
    .S1(_2121_),
    .X(_2312_));
 sky130_fd_sc_hd__mux2i_1 _2991_ (.A0(\registers[18][8] ),
    .A1(\registers[22][8] ),
    .S(_1759_),
    .Y(_2313_));
 sky130_fd_sc_hd__mux2i_1 _2992_ (.A0(\registers[16][8] ),
    .A1(\registers[20][8] ),
    .S(_1837_),
    .Y(_2314_));
 sky130_fd_sc_hd__a221oi_1 _2993_ (.A1(_1769_),
    .A2(_2313_),
    .B1(_2314_),
    .B2(_1765_),
    .C1(_1772_),
    .Y(_2315_));
 sky130_fd_sc_hd__o21ai_1 _2994_ (.A1(_1751_),
    .A2(_2312_),
    .B1(_2315_),
    .Y(_2316_));
 sky130_fd_sc_hd__mux4_1 _2995_ (.A0(\registers[24][8] ),
    .A1(\registers[26][8] ),
    .A2(\registers[28][8] ),
    .A3(\registers[30][8] ),
    .S0(_1754_),
    .S1(_1790_),
    .X(_2317_));
 sky130_fd_sc_hd__mux4_1 _2996_ (.A0(\registers[25][8] ),
    .A1(\registers[27][8] ),
    .A2(\registers[29][8] ),
    .A3(\registers[31][8] ),
    .S0(_2193_),
    .S1(_1802_),
    .X(_2318_));
 sky130_fd_sc_hd__a22oi_4 _2997_ (.A1(_1809_),
    .A2(_2317_),
    .B1(_2318_),
    .B2(_1811_),
    .Y(_2319_));
 sky130_fd_sc_hd__mux4_1 _2998_ (.A0(\registers[8][8] ),
    .A1(\registers[9][8] ),
    .A2(\registers[10][8] ),
    .A3(\registers[11][8] ),
    .S0(_1787_),
    .S1(_1775_),
    .X(_2320_));
 sky130_fd_sc_hd__mux4_1 _2999_ (.A0(\registers[12][8] ),
    .A1(\registers[13][8] ),
    .A2(\registers[14][8] ),
    .A3(\registers[15][8] ),
    .S0(_1899_),
    .S1(_2180_),
    .X(_2321_));
 sky130_fd_sc_hd__mux2i_1 _3000_ (.A0(_2320_),
    .A1(_2321_),
    .S(_2198_),
    .Y(_2322_));
 sky130_fd_sc_hd__mux4_1 _3001_ (.A0(\registers[1][8] ),
    .A1(\registers[3][8] ),
    .A2(\registers[5][8] ),
    .A3(\registers[7][8] ),
    .S0(_1821_),
    .S1(_1822_),
    .X(_2323_));
 sky130_fd_sc_hd__mux4_1 _3002_ (.A0(\registers[0][8] ),
    .A1(\registers[2][8] ),
    .A2(\registers[4][8] ),
    .A3(\registers[6][8] ),
    .S0(_2201_),
    .S1(_1789_),
    .X(_2324_));
 sky130_fd_sc_hd__mux2i_1 _3003_ (.A0(_2323_),
    .A1(_2324_),
    .S(_1749_),
    .Y(_2325_));
 sky130_fd_sc_hd__a221o_2 _3004_ (.A1(_1825_),
    .A2(_2322_),
    .B1(_2325_),
    .B2(_1792_),
    .C1(_1797_),
    .X(_2326_));
 sky130_fd_sc_hd__a31oi_4 _3005_ (.A1(_1745_),
    .A2(_2316_),
    .A3(_2319_),
    .B1(_2326_),
    .Y(_0096_));
 sky130_fd_sc_hd__mux4_1 _3006_ (.A0(\registers[17][9] ),
    .A1(\registers[19][9] ),
    .A2(\registers[21][9] ),
    .A3(\registers[23][9] ),
    .S0(_1780_),
    .S1(_1776_),
    .X(_2327_));
 sky130_fd_sc_hd__mux2i_1 _3007_ (.A0(\registers[18][9] ),
    .A1(\registers[22][9] ),
    .S(_1759_),
    .Y(_2328_));
 sky130_fd_sc_hd__mux2i_1 _3008_ (.A0(\registers[16][9] ),
    .A1(\registers[20][9] ),
    .S(_1837_),
    .Y(_2329_));
 sky130_fd_sc_hd__a221oi_1 _3009_ (.A1(_1769_),
    .A2(_2328_),
    .B1(_2329_),
    .B2(_1765_),
    .C1(_1772_),
    .Y(_2330_));
 sky130_fd_sc_hd__o21ai_1 _3010_ (.A1(_1751_),
    .A2(_2327_),
    .B1(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__mux4_1 _3011_ (.A0(\registers[24][9] ),
    .A1(\registers[26][9] ),
    .A2(\registers[28][9] ),
    .A3(\registers[30][9] ),
    .S0(_1754_),
    .S1(_1790_),
    .X(_2332_));
 sky130_fd_sc_hd__mux4_1 _3012_ (.A0(\registers[25][9] ),
    .A1(\registers[27][9] ),
    .A2(\registers[29][9] ),
    .A3(\registers[31][9] ),
    .S0(_2193_),
    .S1(_1802_),
    .X(_2333_));
 sky130_fd_sc_hd__a22oi_4 _3013_ (.A1(_1809_),
    .A2(_2332_),
    .B1(_2333_),
    .B2(_1811_),
    .Y(_2334_));
 sky130_fd_sc_hd__mux4_1 _3014_ (.A0(\registers[0][9] ),
    .A1(\registers[1][9] ),
    .A2(\registers[2][9] ),
    .A3(\registers[3][9] ),
    .S0(_1787_),
    .S1(_1775_),
    .X(_2335_));
 sky130_fd_sc_hd__mux4_1 _3015_ (.A0(\registers[4][9] ),
    .A1(\registers[5][9] ),
    .A2(\registers[6][9] ),
    .A3(\registers[7][9] ),
    .S0(_1899_),
    .S1(_1764_),
    .X(_2336_));
 sky130_fd_sc_hd__mux2i_1 _3016_ (.A0(_2335_),
    .A1(_2336_),
    .S(_2198_),
    .Y(_2337_));
 sky130_fd_sc_hd__mux4_1 _3017_ (.A0(\registers[9][9] ),
    .A1(\registers[11][9] ),
    .A2(\registers[13][9] ),
    .A3(\registers[15][9] ),
    .S0(_1821_),
    .S1(_1822_),
    .X(_2338_));
 sky130_fd_sc_hd__mux4_1 _3018_ (.A0(\registers[8][9] ),
    .A1(\registers[10][9] ),
    .A2(\registers[12][9] ),
    .A3(\registers[14][9] ),
    .S0(_2201_),
    .S1(_1789_),
    .X(_2339_));
 sky130_fd_sc_hd__mux2i_1 _3019_ (.A0(_2338_),
    .A1(_2339_),
    .S(_1749_),
    .Y(_2340_));
 sky130_fd_sc_hd__a221o_2 _3020_ (.A1(_1923_),
    .A2(_2337_),
    .B1(_2340_),
    .B2(_1784_),
    .C1(_1797_),
    .X(_2341_));
 sky130_fd_sc_hd__a31oi_4 _3021_ (.A1(_1745_),
    .A2(_2331_),
    .A3(_2334_),
    .B1(_2341_),
    .Y(_0097_));
 sky130_fd_sc_hd__buf_2 _3022_ (.A(net11),
    .X(_2342_));
 sky130_fd_sc_hd__nor2_4 _3023_ (.A(_1124_),
    .B(_1128_),
    .Y(_2343_));
 sky130_fd_sc_hd__clkbuf_4 _3024_ (.A(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__and2_0 _3025_ (.A(_2342_),
    .B(_2344_),
    .X(_0098_));
 sky130_fd_sc_hd__buf_2 _3026_ (.A(net12),
    .X(_2345_));
 sky130_fd_sc_hd__and2_0 _3027_ (.A(_2345_),
    .B(_2344_),
    .X(_0099_));
 sky130_fd_sc_hd__buf_2 _3028_ (.A(net13),
    .X(_2346_));
 sky130_fd_sc_hd__and2_0 _3029_ (.A(_2346_),
    .B(_2344_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_4 _3030_ (.A(net14),
    .X(_2347_));
 sky130_fd_sc_hd__and2_0 _3031_ (.A(_2347_),
    .B(_2344_),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_4 _3032_ (.A(net15),
    .X(_2348_));
 sky130_fd_sc_hd__and2_0 _3033_ (.A(_2348_),
    .B(_2344_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_4 _3034_ (.A(net16),
    .X(_2349_));
 sky130_fd_sc_hd__and2_0 _3035_ (.A(_2349_),
    .B(_2344_),
    .X(_0103_));
 sky130_fd_sc_hd__buf_4 _3036_ (.A(net17),
    .X(_2350_));
 sky130_fd_sc_hd__and2_0 _3037_ (.A(_2350_),
    .B(_2344_),
    .X(_0104_));
 sky130_fd_sc_hd__buf_4 _3038_ (.A(net18),
    .X(_2351_));
 sky130_fd_sc_hd__and2_0 _3039_ (.A(_2351_),
    .B(_2344_),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_4 _3040_ (.A(net19),
    .X(_2352_));
 sky130_fd_sc_hd__and2_0 _3041_ (.A(_2352_),
    .B(_2344_),
    .X(_0106_));
 sky130_fd_sc_hd__buf_4 _3042_ (.A(net20),
    .X(_2353_));
 sky130_fd_sc_hd__and2_0 _3043_ (.A(_2353_),
    .B(_2344_),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_4 _3044_ (.A(net21),
    .X(_2354_));
 sky130_fd_sc_hd__buf_4 _3045_ (.A(_2343_),
    .X(_2355_));
 sky130_fd_sc_hd__and2_0 _3046_ (.A(_2354_),
    .B(_2355_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_4 _3047_ (.A(net22),
    .X(_2356_));
 sky130_fd_sc_hd__and2_0 _3048_ (.A(_2356_),
    .B(_2355_),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_4 _3049_ (.A(net23),
    .X(_2357_));
 sky130_fd_sc_hd__and2_0 _3050_ (.A(_2357_),
    .B(_2355_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_4 _3051_ (.A(net24),
    .X(_2358_));
 sky130_fd_sc_hd__and2_0 _3052_ (.A(_2358_),
    .B(_2355_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_4 _3053_ (.A(net25),
    .X(_2359_));
 sky130_fd_sc_hd__and2_0 _3054_ (.A(_2359_),
    .B(_2355_),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_4 _3055_ (.A(net26),
    .X(_2360_));
 sky130_fd_sc_hd__and2_0 _3056_ (.A(_2360_),
    .B(_2355_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_4 _3057_ (.A(net27),
    .X(_2361_));
 sky130_fd_sc_hd__and2_0 _3058_ (.A(_2361_),
    .B(_2355_),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_4 _3059_ (.A(net28),
    .X(_2362_));
 sky130_fd_sc_hd__and2_0 _3060_ (.A(_2362_),
    .B(_2355_),
    .X(_0115_));
 sky130_fd_sc_hd__clkbuf_4 _3061_ (.A(net29),
    .X(_2363_));
 sky130_fd_sc_hd__and2_0 _3062_ (.A(_2363_),
    .B(_2355_),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_4 _3063_ (.A(net30),
    .X(_2364_));
 sky130_fd_sc_hd__and2_0 _3064_ (.A(_2364_),
    .B(_2355_),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_4 _3065_ (.A(net31),
    .X(_2365_));
 sky130_fd_sc_hd__buf_4 _3066_ (.A(_2343_),
    .X(_2366_));
 sky130_fd_sc_hd__and2_0 _3067_ (.A(_2365_),
    .B(_2366_),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_4 _3068_ (.A(net32),
    .X(_2367_));
 sky130_fd_sc_hd__and2_0 _3069_ (.A(_2367_),
    .B(_2366_),
    .X(_0119_));
 sky130_fd_sc_hd__buf_4 _3070_ (.A(net33),
    .X(_2368_));
 sky130_fd_sc_hd__and2_0 _3071_ (.A(_2368_),
    .B(_2366_),
    .X(_0120_));
 sky130_fd_sc_hd__buf_4 _3072_ (.A(net34),
    .X(_2369_));
 sky130_fd_sc_hd__and2_0 _3073_ (.A(_2369_),
    .B(_2366_),
    .X(_0121_));
 sky130_fd_sc_hd__clkbuf_4 _3074_ (.A(net35),
    .X(_2370_));
 sky130_fd_sc_hd__and2_0 _3075_ (.A(_2370_),
    .B(_2366_),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_4 _3076_ (.A(net36),
    .X(_2371_));
 sky130_fd_sc_hd__and2_0 _3077_ (.A(_2371_),
    .B(_2366_),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_4 _3078_ (.A(net37),
    .X(_2372_));
 sky130_fd_sc_hd__and2_0 _3079_ (.A(_2372_),
    .B(_2366_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_4 _3080_ (.A(net38),
    .X(_2373_));
 sky130_fd_sc_hd__and2_0 _3081_ (.A(_2373_),
    .B(_2366_),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_4 _3082_ (.A(net39),
    .X(_2374_));
 sky130_fd_sc_hd__and2_0 _3083_ (.A(_2374_),
    .B(_2366_),
    .X(_0126_));
 sky130_fd_sc_hd__buf_2 _3084_ (.A(net40),
    .X(_2375_));
 sky130_fd_sc_hd__and2_0 _3085_ (.A(_2375_),
    .B(_2366_),
    .X(_0127_));
 sky130_fd_sc_hd__buf_2 _3086_ (.A(net41),
    .X(_2376_));
 sky130_fd_sc_hd__and2_0 _3087_ (.A(_2376_),
    .B(_2343_),
    .X(_0128_));
 sky130_fd_sc_hd__buf_2 _3088_ (.A(net42),
    .X(_2377_));
 sky130_fd_sc_hd__and2_0 _3089_ (.A(_2377_),
    .B(_2343_),
    .X(_0129_));
 sky130_fd_sc_hd__nor2_4 _3090_ (.A(_1131_),
    .B(_1133_),
    .Y(_2378_));
 sky130_fd_sc_hd__buf_4 _3091_ (.A(_2378_),
    .X(_2379_));
 sky130_fd_sc_hd__and2_0 _3092_ (.A(_2342_),
    .B(_2379_),
    .X(_0130_));
 sky130_fd_sc_hd__and2_0 _3093_ (.A(_2345_),
    .B(_2379_),
    .X(_0131_));
 sky130_fd_sc_hd__and2_0 _3094_ (.A(_2346_),
    .B(_2379_),
    .X(_0132_));
 sky130_fd_sc_hd__and2_0 _3095_ (.A(_2347_),
    .B(_2379_),
    .X(_0133_));
 sky130_fd_sc_hd__and2_0 _3096_ (.A(_2348_),
    .B(_2379_),
    .X(_0134_));
 sky130_fd_sc_hd__and2_0 _3097_ (.A(_2349_),
    .B(_2379_),
    .X(_0135_));
 sky130_fd_sc_hd__and2_0 _3098_ (.A(_2350_),
    .B(_2379_),
    .X(_0136_));
 sky130_fd_sc_hd__and2_0 _3099_ (.A(_2351_),
    .B(_2379_),
    .X(_0137_));
 sky130_fd_sc_hd__and2_0 _3100_ (.A(_2352_),
    .B(_2379_),
    .X(_0138_));
 sky130_fd_sc_hd__and2_0 _3101_ (.A(_2353_),
    .B(_2379_),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_4 _3102_ (.A(_2378_),
    .X(_2380_));
 sky130_fd_sc_hd__and2_0 _3103_ (.A(_2354_),
    .B(_2380_),
    .X(_0140_));
 sky130_fd_sc_hd__and2_0 _3104_ (.A(_2356_),
    .B(_2380_),
    .X(_0141_));
 sky130_fd_sc_hd__and2_0 _3105_ (.A(_2357_),
    .B(_2380_),
    .X(_0142_));
 sky130_fd_sc_hd__and2_0 _3106_ (.A(_2358_),
    .B(_2380_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_0 _3107_ (.A(_2359_),
    .B(_2380_),
    .X(_0144_));
 sky130_fd_sc_hd__and2_0 _3108_ (.A(_2360_),
    .B(_2380_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_0 _3109_ (.A(_2361_),
    .B(_2380_),
    .X(_0146_));
 sky130_fd_sc_hd__and2_0 _3110_ (.A(_2362_),
    .B(_2380_),
    .X(_0147_));
 sky130_fd_sc_hd__and2_0 _3111_ (.A(_2363_),
    .B(_2380_),
    .X(_0148_));
 sky130_fd_sc_hd__and2_0 _3112_ (.A(_2364_),
    .B(_2380_),
    .X(_0149_));
 sky130_fd_sc_hd__buf_4 _3113_ (.A(_2378_),
    .X(_2381_));
 sky130_fd_sc_hd__and2_0 _3114_ (.A(_2365_),
    .B(_2381_),
    .X(_0150_));
 sky130_fd_sc_hd__and2_0 _3115_ (.A(_2367_),
    .B(_2381_),
    .X(_0151_));
 sky130_fd_sc_hd__and2_0 _3116_ (.A(_2368_),
    .B(_2381_),
    .X(_0152_));
 sky130_fd_sc_hd__and2_0 _3117_ (.A(_2369_),
    .B(_2381_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_0 _3118_ (.A(_2370_),
    .B(_2381_),
    .X(_0154_));
 sky130_fd_sc_hd__and2_0 _3119_ (.A(_2371_),
    .B(_2381_),
    .X(_0155_));
 sky130_fd_sc_hd__and2_0 _3120_ (.A(_2372_),
    .B(_2381_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_0 _3121_ (.A(_2373_),
    .B(_2381_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_0 _3122_ (.A(_2374_),
    .B(_2381_),
    .X(_0158_));
 sky130_fd_sc_hd__and2_0 _3123_ (.A(_2375_),
    .B(_2381_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_0 _3124_ (.A(_2376_),
    .B(_2378_),
    .X(_0160_));
 sky130_fd_sc_hd__and2_0 _3125_ (.A(_2377_),
    .B(_2378_),
    .X(_0161_));
 sky130_fd_sc_hd__nor2_4 _3126_ (.A(_1131_),
    .B(_1135_),
    .Y(_2382_));
 sky130_fd_sc_hd__clkbuf_8 _3127_ (.A(_2382_),
    .X(_2383_));
 sky130_fd_sc_hd__and2_0 _3128_ (.A(_2342_),
    .B(_2383_),
    .X(_0162_));
 sky130_fd_sc_hd__and2_0 _3129_ (.A(_2345_),
    .B(_2383_),
    .X(_0163_));
 sky130_fd_sc_hd__and2_0 _3130_ (.A(_2346_),
    .B(_2383_),
    .X(_0164_));
 sky130_fd_sc_hd__and2_0 _3131_ (.A(_2347_),
    .B(_2383_),
    .X(_0165_));
 sky130_fd_sc_hd__and2_0 _3132_ (.A(_2348_),
    .B(_2383_),
    .X(_0166_));
 sky130_fd_sc_hd__and2_0 _3133_ (.A(_2349_),
    .B(_2383_),
    .X(_0167_));
 sky130_fd_sc_hd__and2_0 _3134_ (.A(_2350_),
    .B(_2383_),
    .X(_0168_));
 sky130_fd_sc_hd__and2_0 _3135_ (.A(_2351_),
    .B(_2383_),
    .X(_0169_));
 sky130_fd_sc_hd__and2_0 _3136_ (.A(_2352_),
    .B(_2383_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_0 _3137_ (.A(_2353_),
    .B(_2383_),
    .X(_0171_));
 sky130_fd_sc_hd__buf_2 _3138_ (.A(_2382_),
    .X(_2384_));
 sky130_fd_sc_hd__and2_0 _3139_ (.A(_2354_),
    .B(_2384_),
    .X(_0172_));
 sky130_fd_sc_hd__and2_0 _3140_ (.A(_2356_),
    .B(_2384_),
    .X(_0173_));
 sky130_fd_sc_hd__and2_0 _3141_ (.A(_2357_),
    .B(_2384_),
    .X(_0174_));
 sky130_fd_sc_hd__and2_0 _3142_ (.A(_2358_),
    .B(_2384_),
    .X(_0175_));
 sky130_fd_sc_hd__and2_0 _3143_ (.A(_2359_),
    .B(_2384_),
    .X(_0176_));
 sky130_fd_sc_hd__and2_0 _3144_ (.A(_2360_),
    .B(_2384_),
    .X(_0177_));
 sky130_fd_sc_hd__and2_0 _3145_ (.A(_2361_),
    .B(_2384_),
    .X(_0178_));
 sky130_fd_sc_hd__and2_0 _3146_ (.A(_2362_),
    .B(_2384_),
    .X(_0179_));
 sky130_fd_sc_hd__and2_0 _3147_ (.A(_2363_),
    .B(_2384_),
    .X(_0180_));
 sky130_fd_sc_hd__and2_0 _3148_ (.A(_2364_),
    .B(_2384_),
    .X(_0181_));
 sky130_fd_sc_hd__buf_4 _3149_ (.A(_2382_),
    .X(_2385_));
 sky130_fd_sc_hd__and2_0 _3150_ (.A(_2365_),
    .B(_2385_),
    .X(_0182_));
 sky130_fd_sc_hd__and2_0 _3151_ (.A(_2367_),
    .B(_2385_),
    .X(_0183_));
 sky130_fd_sc_hd__and2_0 _3152_ (.A(_2368_),
    .B(_2385_),
    .X(_0184_));
 sky130_fd_sc_hd__and2_0 _3153_ (.A(_2369_),
    .B(_2385_),
    .X(_0185_));
 sky130_fd_sc_hd__and2_0 _3154_ (.A(_2370_),
    .B(_2385_),
    .X(_0186_));
 sky130_fd_sc_hd__and2_0 _3155_ (.A(_2371_),
    .B(_2385_),
    .X(_0187_));
 sky130_fd_sc_hd__and2_0 _3156_ (.A(_2372_),
    .B(_2385_),
    .X(_0188_));
 sky130_fd_sc_hd__and2_0 _3157_ (.A(_2373_),
    .B(_2385_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_0 _3158_ (.A(_2374_),
    .B(_2385_),
    .X(_0190_));
 sky130_fd_sc_hd__and2_0 _3159_ (.A(_2375_),
    .B(_2385_),
    .X(_0191_));
 sky130_fd_sc_hd__and2_0 _3160_ (.A(_2376_),
    .B(_2382_),
    .X(_0192_));
 sky130_fd_sc_hd__and2_0 _3161_ (.A(_2377_),
    .B(_2382_),
    .X(_0193_));
 sky130_fd_sc_hd__nor2_8 _3162_ (.A(_1128_),
    .B(_1136_),
    .Y(_2386_));
 sky130_fd_sc_hd__buf_4 _3163_ (.A(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__and2_0 _3164_ (.A(_2342_),
    .B(_2387_),
    .X(_0194_));
 sky130_fd_sc_hd__and2_0 _3165_ (.A(_2345_),
    .B(_2387_),
    .X(_0195_));
 sky130_fd_sc_hd__and2_0 _3166_ (.A(_2346_),
    .B(_2387_),
    .X(_0196_));
 sky130_fd_sc_hd__and2_0 _3167_ (.A(_2347_),
    .B(_2387_),
    .X(_0197_));
 sky130_fd_sc_hd__and2_0 _3168_ (.A(_2348_),
    .B(_2387_),
    .X(_0198_));
 sky130_fd_sc_hd__and2_0 _3169_ (.A(_2349_),
    .B(_2387_),
    .X(_0199_));
 sky130_fd_sc_hd__and2_0 _3170_ (.A(_2350_),
    .B(_2387_),
    .X(_0200_));
 sky130_fd_sc_hd__and2_0 _3171_ (.A(_2351_),
    .B(_2387_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_0 _3172_ (.A(_2352_),
    .B(_2387_),
    .X(_0202_));
 sky130_fd_sc_hd__and2_0 _3173_ (.A(_2353_),
    .B(_2387_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_4 _3174_ (.A(_2386_),
    .X(_2388_));
 sky130_fd_sc_hd__and2_0 _3175_ (.A(_2354_),
    .B(_2388_),
    .X(_0204_));
 sky130_fd_sc_hd__and2_0 _3176_ (.A(_2356_),
    .B(_2388_),
    .X(_0205_));
 sky130_fd_sc_hd__and2_0 _3177_ (.A(_2357_),
    .B(_2388_),
    .X(_0206_));
 sky130_fd_sc_hd__and2_0 _3178_ (.A(_2358_),
    .B(_2388_),
    .X(_0207_));
 sky130_fd_sc_hd__and2_0 _3179_ (.A(_2359_),
    .B(_2388_),
    .X(_0208_));
 sky130_fd_sc_hd__and2_0 _3180_ (.A(_2360_),
    .B(_2388_),
    .X(_0209_));
 sky130_fd_sc_hd__and2_0 _3181_ (.A(_2361_),
    .B(_2388_),
    .X(_0210_));
 sky130_fd_sc_hd__and2_0 _3182_ (.A(_2362_),
    .B(_2388_),
    .X(_0211_));
 sky130_fd_sc_hd__and2_0 _3183_ (.A(_2363_),
    .B(_2388_),
    .X(_0212_));
 sky130_fd_sc_hd__and2_0 _3184_ (.A(_2364_),
    .B(_2388_),
    .X(_0213_));
 sky130_fd_sc_hd__buf_4 _3185_ (.A(_2386_),
    .X(_2389_));
 sky130_fd_sc_hd__and2_0 _3186_ (.A(_2365_),
    .B(_2389_),
    .X(_0214_));
 sky130_fd_sc_hd__and2_0 _3187_ (.A(_2367_),
    .B(_2389_),
    .X(_0215_));
 sky130_fd_sc_hd__and2_0 _3188_ (.A(_2368_),
    .B(_2389_),
    .X(_0216_));
 sky130_fd_sc_hd__and2_0 _3189_ (.A(_2369_),
    .B(_2389_),
    .X(_0217_));
 sky130_fd_sc_hd__and2_0 _3190_ (.A(_2370_),
    .B(_2389_),
    .X(_0218_));
 sky130_fd_sc_hd__and2_0 _3191_ (.A(_2371_),
    .B(_2389_),
    .X(_0219_));
 sky130_fd_sc_hd__and2_0 _3192_ (.A(_2372_),
    .B(_2389_),
    .X(_0220_));
 sky130_fd_sc_hd__and2_0 _3193_ (.A(_2373_),
    .B(_2389_),
    .X(_0221_));
 sky130_fd_sc_hd__and2_0 _3194_ (.A(_2374_),
    .B(_2389_),
    .X(_0222_));
 sky130_fd_sc_hd__and2_0 _3195_ (.A(_2375_),
    .B(_2389_),
    .X(_0223_));
 sky130_fd_sc_hd__and2_0 _3196_ (.A(_2376_),
    .B(_2386_),
    .X(_0224_));
 sky130_fd_sc_hd__and2_0 _3197_ (.A(_2377_),
    .B(_2386_),
    .X(_0225_));
 sky130_fd_sc_hd__nor2_8 _3198_ (.A(_1136_),
    .B(_1138_),
    .Y(_2390_));
 sky130_fd_sc_hd__buf_4 _3199_ (.A(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__and2_0 _3200_ (.A(_2342_),
    .B(_2391_),
    .X(_0226_));
 sky130_fd_sc_hd__and2_0 _3201_ (.A(_2345_),
    .B(_2391_),
    .X(_0227_));
 sky130_fd_sc_hd__and2_0 _3202_ (.A(_2346_),
    .B(_2391_),
    .X(_0228_));
 sky130_fd_sc_hd__and2_0 _3203_ (.A(_2347_),
    .B(_2391_),
    .X(_0229_));
 sky130_fd_sc_hd__and2_0 _3204_ (.A(_2348_),
    .B(_2391_),
    .X(_0230_));
 sky130_fd_sc_hd__and2_0 _3205_ (.A(_2349_),
    .B(_2391_),
    .X(_0231_));
 sky130_fd_sc_hd__and2_0 _3206_ (.A(_2350_),
    .B(_2391_),
    .X(_0232_));
 sky130_fd_sc_hd__and2_0 _3207_ (.A(_2351_),
    .B(_2391_),
    .X(_0233_));
 sky130_fd_sc_hd__and2_0 _3208_ (.A(_2352_),
    .B(_2391_),
    .X(_0234_));
 sky130_fd_sc_hd__and2_0 _3209_ (.A(_2353_),
    .B(_2391_),
    .X(_0235_));
 sky130_fd_sc_hd__buf_2 _3210_ (.A(_2390_),
    .X(_2392_));
 sky130_fd_sc_hd__and2_0 _3211_ (.A(_2354_),
    .B(_2392_),
    .X(_0236_));
 sky130_fd_sc_hd__and2_0 _3212_ (.A(_2356_),
    .B(_2392_),
    .X(_0237_));
 sky130_fd_sc_hd__and2_0 _3213_ (.A(_2357_),
    .B(_2392_),
    .X(_0238_));
 sky130_fd_sc_hd__and2_0 _3214_ (.A(_2358_),
    .B(_2392_),
    .X(_0239_));
 sky130_fd_sc_hd__and2_0 _3215_ (.A(_2359_),
    .B(_2392_),
    .X(_0240_));
 sky130_fd_sc_hd__and2_0 _3216_ (.A(_2360_),
    .B(_2392_),
    .X(_0241_));
 sky130_fd_sc_hd__and2_0 _3217_ (.A(_2361_),
    .B(_2392_),
    .X(_0242_));
 sky130_fd_sc_hd__and2_0 _3218_ (.A(_2362_),
    .B(_2392_),
    .X(_0243_));
 sky130_fd_sc_hd__and2_0 _3219_ (.A(_2363_),
    .B(_2392_),
    .X(_0244_));
 sky130_fd_sc_hd__and2_0 _3220_ (.A(_2364_),
    .B(_2392_),
    .X(_0245_));
 sky130_fd_sc_hd__buf_4 _3221_ (.A(_2390_),
    .X(_2393_));
 sky130_fd_sc_hd__and2_0 _3222_ (.A(_2365_),
    .B(_2393_),
    .X(_0246_));
 sky130_fd_sc_hd__and2_0 _3223_ (.A(_2367_),
    .B(_2393_),
    .X(_0247_));
 sky130_fd_sc_hd__and2_0 _3224_ (.A(_2368_),
    .B(_2393_),
    .X(_0248_));
 sky130_fd_sc_hd__and2_0 _3225_ (.A(_2369_),
    .B(_2393_),
    .X(_0249_));
 sky130_fd_sc_hd__and2_0 _3226_ (.A(_2370_),
    .B(_2393_),
    .X(_0250_));
 sky130_fd_sc_hd__and2_0 _3227_ (.A(_2371_),
    .B(_2393_),
    .X(_0251_));
 sky130_fd_sc_hd__and2_0 _3228_ (.A(_2372_),
    .B(_2393_),
    .X(_0252_));
 sky130_fd_sc_hd__and2_0 _3229_ (.A(_2373_),
    .B(_2393_),
    .X(_0253_));
 sky130_fd_sc_hd__and2_0 _3230_ (.A(_2374_),
    .B(_2393_),
    .X(_0254_));
 sky130_fd_sc_hd__and2_0 _3231_ (.A(_2375_),
    .B(_2393_),
    .X(_0255_));
 sky130_fd_sc_hd__and2_0 _3232_ (.A(_2376_),
    .B(_2390_),
    .X(_0256_));
 sky130_fd_sc_hd__and2_0 _3233_ (.A(_2377_),
    .B(_2390_),
    .X(_0257_));
 sky130_fd_sc_hd__nor2_8 _3234_ (.A(_1132_),
    .B(_1136_),
    .Y(_2394_));
 sky130_fd_sc_hd__buf_4 _3235_ (.A(_2394_),
    .X(_2395_));
 sky130_fd_sc_hd__and2_0 _3236_ (.A(_2342_),
    .B(_2395_),
    .X(_0258_));
 sky130_fd_sc_hd__and2_0 _3237_ (.A(_2345_),
    .B(_2395_),
    .X(_0259_));
 sky130_fd_sc_hd__and2_0 _3238_ (.A(_2346_),
    .B(_2395_),
    .X(_0260_));
 sky130_fd_sc_hd__and2_0 _3239_ (.A(_2347_),
    .B(_2395_),
    .X(_0261_));
 sky130_fd_sc_hd__and2_0 _3240_ (.A(_2348_),
    .B(_2395_),
    .X(_0262_));
 sky130_fd_sc_hd__and2_0 _3241_ (.A(_2349_),
    .B(_2395_),
    .X(_0263_));
 sky130_fd_sc_hd__and2_0 _3242_ (.A(_2350_),
    .B(_2395_),
    .X(_0264_));
 sky130_fd_sc_hd__and2_0 _3243_ (.A(_2351_),
    .B(_2395_),
    .X(_0265_));
 sky130_fd_sc_hd__and2_0 _3244_ (.A(_2352_),
    .B(_2395_),
    .X(_0266_));
 sky130_fd_sc_hd__and2_0 _3245_ (.A(_2353_),
    .B(_2395_),
    .X(_0267_));
 sky130_fd_sc_hd__buf_2 _3246_ (.A(_2394_),
    .X(_2396_));
 sky130_fd_sc_hd__and2_0 _3247_ (.A(_2354_),
    .B(_2396_),
    .X(_0268_));
 sky130_fd_sc_hd__and2_0 _3248_ (.A(_2356_),
    .B(_2396_),
    .X(_0269_));
 sky130_fd_sc_hd__and2_0 _3249_ (.A(_2357_),
    .B(_2396_),
    .X(_0270_));
 sky130_fd_sc_hd__and2_0 _3250_ (.A(_2358_),
    .B(_2396_),
    .X(_0271_));
 sky130_fd_sc_hd__and2_0 _3251_ (.A(_2359_),
    .B(_2396_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_0 _3252_ (.A(_2360_),
    .B(_2396_),
    .X(_0273_));
 sky130_fd_sc_hd__and2_0 _3253_ (.A(_2361_),
    .B(_2396_),
    .X(_0274_));
 sky130_fd_sc_hd__and2_0 _3254_ (.A(_2362_),
    .B(_2396_),
    .X(_0275_));
 sky130_fd_sc_hd__and2_0 _3255_ (.A(_2363_),
    .B(_2396_),
    .X(_0276_));
 sky130_fd_sc_hd__and2_0 _3256_ (.A(_2364_),
    .B(_2396_),
    .X(_0277_));
 sky130_fd_sc_hd__clkbuf_8 _3257_ (.A(_2394_),
    .X(_2397_));
 sky130_fd_sc_hd__and2_0 _3258_ (.A(_2365_),
    .B(_2397_),
    .X(_0278_));
 sky130_fd_sc_hd__and2_0 _3259_ (.A(_2367_),
    .B(_2397_),
    .X(_0279_));
 sky130_fd_sc_hd__and2_0 _3260_ (.A(_2368_),
    .B(_2397_),
    .X(_0280_));
 sky130_fd_sc_hd__and2_0 _3261_ (.A(_2369_),
    .B(_2397_),
    .X(_0281_));
 sky130_fd_sc_hd__and2_0 _3262_ (.A(_2370_),
    .B(_2397_),
    .X(_0282_));
 sky130_fd_sc_hd__and2_0 _3263_ (.A(_2371_),
    .B(_2397_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_0 _3264_ (.A(_2372_),
    .B(_2397_),
    .X(_0284_));
 sky130_fd_sc_hd__and2_0 _3265_ (.A(_2373_),
    .B(_2397_),
    .X(_0285_));
 sky130_fd_sc_hd__and2_0 _3266_ (.A(_2374_),
    .B(_2397_),
    .X(_0286_));
 sky130_fd_sc_hd__and2_0 _3267_ (.A(_2375_),
    .B(_2397_),
    .X(_0287_));
 sky130_fd_sc_hd__and2_0 _3268_ (.A(_2376_),
    .B(_2394_),
    .X(_0288_));
 sky130_fd_sc_hd__and2_0 _3269_ (.A(_2377_),
    .B(_2394_),
    .X(_0289_));
 sky130_fd_sc_hd__nor2_8 _3270_ (.A(_1134_),
    .B(_1136_),
    .Y(_2398_));
 sky130_fd_sc_hd__buf_4 _3271_ (.A(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__and2_0 _3272_ (.A(_2342_),
    .B(_2399_),
    .X(_0290_));
 sky130_fd_sc_hd__and2_0 _3273_ (.A(_2345_),
    .B(_2399_),
    .X(_0291_));
 sky130_fd_sc_hd__and2_0 _3274_ (.A(_2346_),
    .B(_2399_),
    .X(_0292_));
 sky130_fd_sc_hd__and2_0 _3275_ (.A(_2347_),
    .B(_2399_),
    .X(_0293_));
 sky130_fd_sc_hd__and2_0 _3276_ (.A(_2348_),
    .B(_2399_),
    .X(_0294_));
 sky130_fd_sc_hd__and2_0 _3277_ (.A(_2349_),
    .B(_2399_),
    .X(_0295_));
 sky130_fd_sc_hd__and2_0 _3278_ (.A(_2350_),
    .B(_2399_),
    .X(_0296_));
 sky130_fd_sc_hd__and2_0 _3279_ (.A(_2351_),
    .B(_2399_),
    .X(_0297_));
 sky130_fd_sc_hd__and2_0 _3280_ (.A(_2352_),
    .B(_2399_),
    .X(_0298_));
 sky130_fd_sc_hd__and2_0 _3281_ (.A(_2353_),
    .B(_2399_),
    .X(_0299_));
 sky130_fd_sc_hd__buf_2 _3282_ (.A(_2398_),
    .X(_2400_));
 sky130_fd_sc_hd__and2_0 _3283_ (.A(_2354_),
    .B(_2400_),
    .X(_0300_));
 sky130_fd_sc_hd__and2_0 _3284_ (.A(_2356_),
    .B(_2400_),
    .X(_0301_));
 sky130_fd_sc_hd__and2_0 _3285_ (.A(_2357_),
    .B(_2400_),
    .X(_0302_));
 sky130_fd_sc_hd__and2_0 _3286_ (.A(_2358_),
    .B(_2400_),
    .X(_0303_));
 sky130_fd_sc_hd__and2_0 _3287_ (.A(_2359_),
    .B(_2400_),
    .X(_0304_));
 sky130_fd_sc_hd__and2_0 _3288_ (.A(_2360_),
    .B(_2400_),
    .X(_0305_));
 sky130_fd_sc_hd__and2_0 _3289_ (.A(_2361_),
    .B(_2400_),
    .X(_0306_));
 sky130_fd_sc_hd__and2_0 _3290_ (.A(_2362_),
    .B(_2400_),
    .X(_0307_));
 sky130_fd_sc_hd__and2_0 _3291_ (.A(_2363_),
    .B(_2400_),
    .X(_0308_));
 sky130_fd_sc_hd__and2_0 _3292_ (.A(_2364_),
    .B(_2400_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_4 _3293_ (.A(_2398_),
    .X(_2401_));
 sky130_fd_sc_hd__and2_0 _3294_ (.A(_2365_),
    .B(_2401_),
    .X(_0310_));
 sky130_fd_sc_hd__and2_0 _3295_ (.A(_2367_),
    .B(_2401_),
    .X(_0311_));
 sky130_fd_sc_hd__and2_0 _3296_ (.A(_2368_),
    .B(_2401_),
    .X(_0312_));
 sky130_fd_sc_hd__and2_0 _3297_ (.A(_2369_),
    .B(_2401_),
    .X(_0313_));
 sky130_fd_sc_hd__and2_0 _3298_ (.A(_2370_),
    .B(_2401_),
    .X(_0314_));
 sky130_fd_sc_hd__and2_0 _3299_ (.A(_2371_),
    .B(_2401_),
    .X(_0315_));
 sky130_fd_sc_hd__and2_0 _3300_ (.A(_2372_),
    .B(_2401_),
    .X(_0316_));
 sky130_fd_sc_hd__and2_0 _3301_ (.A(_2373_),
    .B(_2401_),
    .X(_0317_));
 sky130_fd_sc_hd__and2_0 _3302_ (.A(_2374_),
    .B(_2401_),
    .X(_0318_));
 sky130_fd_sc_hd__and2_0 _3303_ (.A(_2375_),
    .B(_2401_),
    .X(_0319_));
 sky130_fd_sc_hd__and2_0 _3304_ (.A(_2376_),
    .B(_2398_),
    .X(_0320_));
 sky130_fd_sc_hd__and2_0 _3305_ (.A(_2377_),
    .B(_2398_),
    .X(_0321_));
 sky130_fd_sc_hd__nor2_4 _3306_ (.A(_1127_),
    .B(_1140_),
    .Y(_2402_));
 sky130_fd_sc_hd__buf_2 _3307_ (.A(_2402_),
    .X(_2403_));
 sky130_fd_sc_hd__and2_0 _3308_ (.A(_2342_),
    .B(_2403_),
    .X(_0322_));
 sky130_fd_sc_hd__and2_0 _3309_ (.A(_2345_),
    .B(_2403_),
    .X(_0323_));
 sky130_fd_sc_hd__and2_0 _3310_ (.A(_2346_),
    .B(_2403_),
    .X(_0324_));
 sky130_fd_sc_hd__and2_0 _3311_ (.A(_2347_),
    .B(_2403_),
    .X(_0325_));
 sky130_fd_sc_hd__and2_0 _3312_ (.A(_2348_),
    .B(_2403_),
    .X(_0326_));
 sky130_fd_sc_hd__and2_0 _3313_ (.A(_2349_),
    .B(_2403_),
    .X(_0327_));
 sky130_fd_sc_hd__and2_0 _3314_ (.A(_2350_),
    .B(_2403_),
    .X(_0328_));
 sky130_fd_sc_hd__and2_0 _3315_ (.A(_2351_),
    .B(_2403_),
    .X(_0329_));
 sky130_fd_sc_hd__and2_0 _3316_ (.A(_2352_),
    .B(_2403_),
    .X(_0330_));
 sky130_fd_sc_hd__and2_0 _3317_ (.A(_2353_),
    .B(_2403_),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_4 _3318_ (.A(_2402_),
    .X(_2404_));
 sky130_fd_sc_hd__and2_0 _3319_ (.A(_2354_),
    .B(_2404_),
    .X(_0332_));
 sky130_fd_sc_hd__and2_0 _3320_ (.A(_2356_),
    .B(_2404_),
    .X(_0333_));
 sky130_fd_sc_hd__and2_0 _3321_ (.A(_2357_),
    .B(_2404_),
    .X(_0334_));
 sky130_fd_sc_hd__and2_0 _3322_ (.A(_2358_),
    .B(_2404_),
    .X(_0335_));
 sky130_fd_sc_hd__and2_0 _3323_ (.A(_2359_),
    .B(_2404_),
    .X(_0336_));
 sky130_fd_sc_hd__and2_0 _3324_ (.A(_2360_),
    .B(_2404_),
    .X(_0337_));
 sky130_fd_sc_hd__and2_0 _3325_ (.A(_2361_),
    .B(_2404_),
    .X(_0338_));
 sky130_fd_sc_hd__and2_0 _3326_ (.A(_2362_),
    .B(_2404_),
    .X(_0339_));
 sky130_fd_sc_hd__and2_0 _3327_ (.A(_2363_),
    .B(_2404_),
    .X(_0340_));
 sky130_fd_sc_hd__and2_0 _3328_ (.A(_2364_),
    .B(_2404_),
    .X(_0341_));
 sky130_fd_sc_hd__buf_2 _3329_ (.A(_2402_),
    .X(_2405_));
 sky130_fd_sc_hd__and2_0 _3330_ (.A(_2365_),
    .B(_2405_),
    .X(_0342_));
 sky130_fd_sc_hd__and2_0 _3331_ (.A(_2367_),
    .B(_2405_),
    .X(_0343_));
 sky130_fd_sc_hd__and2_0 _3332_ (.A(_2368_),
    .B(_2405_),
    .X(_0344_));
 sky130_fd_sc_hd__and2_0 _3333_ (.A(_2369_),
    .B(_2405_),
    .X(_0345_));
 sky130_fd_sc_hd__and2_0 _3334_ (.A(_2370_),
    .B(_2405_),
    .X(_0346_));
 sky130_fd_sc_hd__and2_0 _3335_ (.A(_2371_),
    .B(_2405_),
    .X(_0347_));
 sky130_fd_sc_hd__and2_0 _3336_ (.A(_2372_),
    .B(_2405_),
    .X(_0348_));
 sky130_fd_sc_hd__and2_0 _3337_ (.A(_2373_),
    .B(_2405_),
    .X(_0349_));
 sky130_fd_sc_hd__and2_0 _3338_ (.A(_2374_),
    .B(_2405_),
    .X(_0350_));
 sky130_fd_sc_hd__and2_0 _3339_ (.A(_2375_),
    .B(_2405_),
    .X(_0351_));
 sky130_fd_sc_hd__and2_0 _3340_ (.A(_2376_),
    .B(_2402_),
    .X(_0352_));
 sky130_fd_sc_hd__and2_0 _3341_ (.A(_2377_),
    .B(_2402_),
    .X(_0353_));
 sky130_fd_sc_hd__nor2_2 _3342_ (.A(_1137_),
    .B(_1140_),
    .Y(_2406_));
 sky130_fd_sc_hd__buf_2 _3343_ (.A(_2406_),
    .X(_2407_));
 sky130_fd_sc_hd__and2_0 _3344_ (.A(_2342_),
    .B(_2407_),
    .X(_0354_));
 sky130_fd_sc_hd__and2_0 _3345_ (.A(_2345_),
    .B(_2407_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_0 _3346_ (.A(_2346_),
    .B(_2407_),
    .X(_0356_));
 sky130_fd_sc_hd__and2_0 _3347_ (.A(_2347_),
    .B(_2407_),
    .X(_0357_));
 sky130_fd_sc_hd__and2_0 _3348_ (.A(_2348_),
    .B(_2407_),
    .X(_0358_));
 sky130_fd_sc_hd__and2_0 _3349_ (.A(_2349_),
    .B(_2407_),
    .X(_0359_));
 sky130_fd_sc_hd__and2_0 _3350_ (.A(_2350_),
    .B(_2407_),
    .X(_0360_));
 sky130_fd_sc_hd__and2_0 _3351_ (.A(_2351_),
    .B(_2407_),
    .X(_0361_));
 sky130_fd_sc_hd__and2_0 _3352_ (.A(_2352_),
    .B(_2407_),
    .X(_0362_));
 sky130_fd_sc_hd__and2_0 _3353_ (.A(_2353_),
    .B(_2407_),
    .X(_0363_));
 sky130_fd_sc_hd__buf_2 _3354_ (.A(_2406_),
    .X(_2408_));
 sky130_fd_sc_hd__and2_0 _3355_ (.A(_2354_),
    .B(_2408_),
    .X(_0364_));
 sky130_fd_sc_hd__and2_0 _3356_ (.A(_2356_),
    .B(_2408_),
    .X(_0365_));
 sky130_fd_sc_hd__and2_0 _3357_ (.A(_2357_),
    .B(_2408_),
    .X(_0366_));
 sky130_fd_sc_hd__and2_0 _3358_ (.A(_2358_),
    .B(_2408_),
    .X(_0367_));
 sky130_fd_sc_hd__and2_0 _3359_ (.A(_2359_),
    .B(_2408_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_0 _3360_ (.A(_2360_),
    .B(_2408_),
    .X(_0369_));
 sky130_fd_sc_hd__and2_0 _3361_ (.A(_2361_),
    .B(_2408_),
    .X(_0370_));
 sky130_fd_sc_hd__and2_0 _3362_ (.A(_2362_),
    .B(_2408_),
    .X(_0371_));
 sky130_fd_sc_hd__and2_0 _3363_ (.A(_2363_),
    .B(_2408_),
    .X(_0372_));
 sky130_fd_sc_hd__and2_0 _3364_ (.A(_2364_),
    .B(_2408_),
    .X(_0373_));
 sky130_fd_sc_hd__buf_2 _3365_ (.A(_2406_),
    .X(_2409_));
 sky130_fd_sc_hd__and2_0 _3366_ (.A(_2365_),
    .B(_2409_),
    .X(_0374_));
 sky130_fd_sc_hd__and2_0 _3367_ (.A(_2367_),
    .B(_2409_),
    .X(_0375_));
 sky130_fd_sc_hd__and2_0 _3368_ (.A(_2368_),
    .B(_2409_),
    .X(_0376_));
 sky130_fd_sc_hd__and2_0 _3369_ (.A(_2369_),
    .B(_2409_),
    .X(_0377_));
 sky130_fd_sc_hd__and2_0 _3370_ (.A(_2370_),
    .B(_2409_),
    .X(_0378_));
 sky130_fd_sc_hd__and2_0 _3371_ (.A(_2371_),
    .B(_2409_),
    .X(_0379_));
 sky130_fd_sc_hd__and2_0 _3372_ (.A(_2372_),
    .B(_2409_),
    .X(_0380_));
 sky130_fd_sc_hd__and2_0 _3373_ (.A(_2373_),
    .B(_2409_),
    .X(_0381_));
 sky130_fd_sc_hd__and2_0 _3374_ (.A(_2374_),
    .B(_2409_),
    .X(_0382_));
 sky130_fd_sc_hd__and2_0 _3375_ (.A(_2375_),
    .B(_2409_),
    .X(_0383_));
 sky130_fd_sc_hd__and2_0 _3376_ (.A(_2376_),
    .B(_2406_),
    .X(_0384_));
 sky130_fd_sc_hd__and2_0 _3377_ (.A(_2377_),
    .B(_2406_),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_4 _3378_ (.A(_1132_),
    .B(_1140_),
    .Y(_2410_));
 sky130_fd_sc_hd__clkbuf_4 _3379_ (.A(_2410_),
    .X(_2411_));
 sky130_fd_sc_hd__and2_0 _3380_ (.A(_2342_),
    .B(_2411_),
    .X(_0386_));
 sky130_fd_sc_hd__and2_0 _3381_ (.A(_2345_),
    .B(_2411_),
    .X(_0387_));
 sky130_fd_sc_hd__and2_0 _3382_ (.A(_2346_),
    .B(_2411_),
    .X(_0388_));
 sky130_fd_sc_hd__and2_0 _3383_ (.A(_2347_),
    .B(_2411_),
    .X(_0389_));
 sky130_fd_sc_hd__and2_0 _3384_ (.A(_2348_),
    .B(_2411_),
    .X(_0390_));
 sky130_fd_sc_hd__and2_0 _3385_ (.A(_2349_),
    .B(_2411_),
    .X(_0391_));
 sky130_fd_sc_hd__and2_0 _3386_ (.A(_2350_),
    .B(_2411_),
    .X(_0392_));
 sky130_fd_sc_hd__and2_0 _3387_ (.A(_2351_),
    .B(_2411_),
    .X(_0393_));
 sky130_fd_sc_hd__and2_0 _3388_ (.A(_2352_),
    .B(_2411_),
    .X(_0394_));
 sky130_fd_sc_hd__and2_0 _3389_ (.A(_2353_),
    .B(_2411_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_4 _3390_ (.A(_2410_),
    .X(_2412_));
 sky130_fd_sc_hd__and2_0 _3391_ (.A(_2354_),
    .B(_2412_),
    .X(_0396_));
 sky130_fd_sc_hd__and2_0 _3392_ (.A(_2356_),
    .B(_2412_),
    .X(_0397_));
 sky130_fd_sc_hd__and2_0 _3393_ (.A(_2357_),
    .B(_2412_),
    .X(_0398_));
 sky130_fd_sc_hd__and2_0 _3394_ (.A(_2358_),
    .B(_2412_),
    .X(_0399_));
 sky130_fd_sc_hd__and2_0 _3395_ (.A(_2359_),
    .B(_2412_),
    .X(_0400_));
 sky130_fd_sc_hd__and2_0 _3396_ (.A(_2360_),
    .B(_2412_),
    .X(_0401_));
 sky130_fd_sc_hd__and2_0 _3397_ (.A(_2361_),
    .B(_2412_),
    .X(_0402_));
 sky130_fd_sc_hd__and2_0 _3398_ (.A(_2362_),
    .B(_2412_),
    .X(_0403_));
 sky130_fd_sc_hd__and2_0 _3399_ (.A(_2363_),
    .B(_2412_),
    .X(_0404_));
 sky130_fd_sc_hd__and2_0 _3400_ (.A(_2364_),
    .B(_2412_),
    .X(_0405_));
 sky130_fd_sc_hd__buf_2 _3401_ (.A(_2410_),
    .X(_2413_));
 sky130_fd_sc_hd__and2_0 _3402_ (.A(_2365_),
    .B(_2413_),
    .X(_0406_));
 sky130_fd_sc_hd__and2_0 _3403_ (.A(_2367_),
    .B(_2413_),
    .X(_0407_));
 sky130_fd_sc_hd__and2_0 _3404_ (.A(_2368_),
    .B(_2413_),
    .X(_0408_));
 sky130_fd_sc_hd__and2_0 _3405_ (.A(_2369_),
    .B(_2413_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_0 _3406_ (.A(_2370_),
    .B(_2413_),
    .X(_0410_));
 sky130_fd_sc_hd__and2_0 _3407_ (.A(_2371_),
    .B(_2413_),
    .X(_0411_));
 sky130_fd_sc_hd__and2_0 _3408_ (.A(_2372_),
    .B(_2413_),
    .X(_0412_));
 sky130_fd_sc_hd__and2_0 _3409_ (.A(_2373_),
    .B(_2413_),
    .X(_0413_));
 sky130_fd_sc_hd__and2_0 _3410_ (.A(_2374_),
    .B(_2413_),
    .X(_0414_));
 sky130_fd_sc_hd__and2_0 _3411_ (.A(_2375_),
    .B(_2413_),
    .X(_0415_));
 sky130_fd_sc_hd__and2_0 _3412_ (.A(_2376_),
    .B(_2410_),
    .X(_0416_));
 sky130_fd_sc_hd__and2_0 _3413_ (.A(_2377_),
    .B(_2410_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_4 _3414_ (.A(net11),
    .X(_2414_));
 sky130_fd_sc_hd__nor2_4 _3415_ (.A(_1134_),
    .B(_1140_),
    .Y(_2415_));
 sky130_fd_sc_hd__clkbuf_4 _3416_ (.A(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__and2_0 _3417_ (.A(_2414_),
    .B(_2416_),
    .X(_0418_));
 sky130_fd_sc_hd__buf_2 _3418_ (.A(net12),
    .X(_2417_));
 sky130_fd_sc_hd__and2_0 _3419_ (.A(_2417_),
    .B(_2416_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_4 _3420_ (.A(net13),
    .X(_2418_));
 sky130_fd_sc_hd__and2_0 _3421_ (.A(_2418_),
    .B(_2416_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_4 _3422_ (.A(net14),
    .X(_2419_));
 sky130_fd_sc_hd__and2_0 _3423_ (.A(_2419_),
    .B(_2416_),
    .X(_0421_));
 sky130_fd_sc_hd__buf_4 _3424_ (.A(net15),
    .X(_2420_));
 sky130_fd_sc_hd__and2_0 _3425_ (.A(_2420_),
    .B(_2416_),
    .X(_0422_));
 sky130_fd_sc_hd__buf_4 _3426_ (.A(net16),
    .X(_2421_));
 sky130_fd_sc_hd__and2_0 _3427_ (.A(_2421_),
    .B(_2416_),
    .X(_0423_));
 sky130_fd_sc_hd__buf_4 _3428_ (.A(net17),
    .X(_2422_));
 sky130_fd_sc_hd__and2_0 _3429_ (.A(_2422_),
    .B(_2416_),
    .X(_0424_));
 sky130_fd_sc_hd__buf_4 _3430_ (.A(net18),
    .X(_2423_));
 sky130_fd_sc_hd__and2_0 _3431_ (.A(_2423_),
    .B(_2416_),
    .X(_0425_));
 sky130_fd_sc_hd__buf_4 _3432_ (.A(net19),
    .X(_2424_));
 sky130_fd_sc_hd__and2_0 _3433_ (.A(_2424_),
    .B(_2416_),
    .X(_0426_));
 sky130_fd_sc_hd__buf_4 _3434_ (.A(net20),
    .X(_2425_));
 sky130_fd_sc_hd__and2_0 _3435_ (.A(_2425_),
    .B(_2416_),
    .X(_0427_));
 sky130_fd_sc_hd__buf_4 _3436_ (.A(net21),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_4 _3437_ (.A(_2415_),
    .X(_2427_));
 sky130_fd_sc_hd__and2_0 _3438_ (.A(_2426_),
    .B(_2427_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_4 _3439_ (.A(net22),
    .X(_2428_));
 sky130_fd_sc_hd__and2_0 _3440_ (.A(_2428_),
    .B(_2427_),
    .X(_0429_));
 sky130_fd_sc_hd__buf_4 _3441_ (.A(net23),
    .X(_2429_));
 sky130_fd_sc_hd__and2_0 _3442_ (.A(_2429_),
    .B(_2427_),
    .X(_0430_));
 sky130_fd_sc_hd__buf_4 _3443_ (.A(net24),
    .X(_2430_));
 sky130_fd_sc_hd__and2_0 _3444_ (.A(_2430_),
    .B(_2427_),
    .X(_0431_));
 sky130_fd_sc_hd__buf_4 _3445_ (.A(net25),
    .X(_2431_));
 sky130_fd_sc_hd__and2_0 _3446_ (.A(_2431_),
    .B(_2427_),
    .X(_0432_));
 sky130_fd_sc_hd__buf_4 _3447_ (.A(net26),
    .X(_2432_));
 sky130_fd_sc_hd__and2_0 _3448_ (.A(_2432_),
    .B(_2427_),
    .X(_0433_));
 sky130_fd_sc_hd__buf_4 _3449_ (.A(net27),
    .X(_2433_));
 sky130_fd_sc_hd__and2_0 _3450_ (.A(_2433_),
    .B(_2427_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_4 _3451_ (.A(net28),
    .X(_2434_));
 sky130_fd_sc_hd__and2_0 _3452_ (.A(_2434_),
    .B(_2427_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_4 _3453_ (.A(net29),
    .X(_2435_));
 sky130_fd_sc_hd__and2_0 _3454_ (.A(_2435_),
    .B(_2427_),
    .X(_0436_));
 sky130_fd_sc_hd__buf_4 _3455_ (.A(net30),
    .X(_2436_));
 sky130_fd_sc_hd__and2_0 _3456_ (.A(_2436_),
    .B(_2427_),
    .X(_0437_));
 sky130_fd_sc_hd__buf_4 _3457_ (.A(net31),
    .X(_2437_));
 sky130_fd_sc_hd__buf_2 _3458_ (.A(_2415_),
    .X(_2438_));
 sky130_fd_sc_hd__and2_0 _3459_ (.A(_2437_),
    .B(_2438_),
    .X(_0438_));
 sky130_fd_sc_hd__buf_4 _3460_ (.A(net32),
    .X(_2439_));
 sky130_fd_sc_hd__and2_0 _3461_ (.A(_2439_),
    .B(_2438_),
    .X(_0439_));
 sky130_fd_sc_hd__buf_6 _3462_ (.A(net33),
    .X(_2440_));
 sky130_fd_sc_hd__and2_0 _3463_ (.A(_2440_),
    .B(_2438_),
    .X(_0440_));
 sky130_fd_sc_hd__buf_6 _3464_ (.A(net34),
    .X(_2441_));
 sky130_fd_sc_hd__and2_0 _3465_ (.A(_2441_),
    .B(_2438_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_8 _3466_ (.A(net35),
    .X(_2442_));
 sky130_fd_sc_hd__and2_0 _3467_ (.A(_2442_),
    .B(_2438_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_4 _3468_ (.A(net36),
    .X(_2443_));
 sky130_fd_sc_hd__and2_0 _3469_ (.A(_2443_),
    .B(_2438_),
    .X(_0443_));
 sky130_fd_sc_hd__buf_4 _3470_ (.A(net37),
    .X(_2444_));
 sky130_fd_sc_hd__and2_0 _3471_ (.A(_2444_),
    .B(_2438_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_4 _3472_ (.A(net38),
    .X(_2445_));
 sky130_fd_sc_hd__and2_0 _3473_ (.A(_2445_),
    .B(_2438_),
    .X(_0445_));
 sky130_fd_sc_hd__buf_4 _3474_ (.A(net39),
    .X(_2446_));
 sky130_fd_sc_hd__and2_0 _3475_ (.A(_2446_),
    .B(_2438_),
    .X(_0446_));
 sky130_fd_sc_hd__buf_2 _3476_ (.A(net40),
    .X(_2447_));
 sky130_fd_sc_hd__and2_0 _3477_ (.A(_2447_),
    .B(_2438_),
    .X(_0447_));
 sky130_fd_sc_hd__buf_2 _3478_ (.A(net41),
    .X(_2448_));
 sky130_fd_sc_hd__and2_0 _3479_ (.A(_2448_),
    .B(_2415_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_4 _3480_ (.A(net42),
    .X(_2449_));
 sky130_fd_sc_hd__and2_0 _3481_ (.A(_2449_),
    .B(_2415_),
    .X(_0449_));
 sky130_fd_sc_hd__nor2_4 _3482_ (.A(_1124_),
    .B(_1138_),
    .Y(_2450_));
 sky130_fd_sc_hd__buf_4 _3483_ (.A(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__and2_0 _3484_ (.A(_2414_),
    .B(_2451_),
    .X(_0450_));
 sky130_fd_sc_hd__and2_0 _3485_ (.A(_2417_),
    .B(_2451_),
    .X(_0451_));
 sky130_fd_sc_hd__and2_0 _3486_ (.A(_2418_),
    .B(_2451_),
    .X(_0452_));
 sky130_fd_sc_hd__and2_0 _3487_ (.A(_2419_),
    .B(_2451_),
    .X(_0453_));
 sky130_fd_sc_hd__and2_0 _3488_ (.A(_2420_),
    .B(_2451_),
    .X(_0454_));
 sky130_fd_sc_hd__and2_0 _3489_ (.A(_2421_),
    .B(_2451_),
    .X(_0455_));
 sky130_fd_sc_hd__and2_0 _3490_ (.A(_2422_),
    .B(_2451_),
    .X(_0456_));
 sky130_fd_sc_hd__and2_0 _3491_ (.A(_2423_),
    .B(_2451_),
    .X(_0457_));
 sky130_fd_sc_hd__and2_0 _3492_ (.A(_2424_),
    .B(_2451_),
    .X(_0458_));
 sky130_fd_sc_hd__and2_0 _3493_ (.A(_2425_),
    .B(_2451_),
    .X(_0459_));
 sky130_fd_sc_hd__buf_4 _3494_ (.A(_2450_),
    .X(_2452_));
 sky130_fd_sc_hd__and2_0 _3495_ (.A(_2426_),
    .B(_2452_),
    .X(_0460_));
 sky130_fd_sc_hd__and2_0 _3496_ (.A(_2428_),
    .B(_2452_),
    .X(_0461_));
 sky130_fd_sc_hd__and2_0 _3497_ (.A(_2429_),
    .B(_2452_),
    .X(_0462_));
 sky130_fd_sc_hd__and2_0 _3498_ (.A(_2430_),
    .B(_2452_),
    .X(_0463_));
 sky130_fd_sc_hd__and2_0 _3499_ (.A(_2431_),
    .B(_2452_),
    .X(_0464_));
 sky130_fd_sc_hd__and2_0 _3500_ (.A(_2432_),
    .B(_2452_),
    .X(_0465_));
 sky130_fd_sc_hd__and2_0 _3501_ (.A(_2433_),
    .B(_2452_),
    .X(_0466_));
 sky130_fd_sc_hd__and2_0 _3502_ (.A(_2434_),
    .B(_2452_),
    .X(_0467_));
 sky130_fd_sc_hd__and2_0 _3503_ (.A(_2435_),
    .B(_2452_),
    .X(_0468_));
 sky130_fd_sc_hd__and2_0 _3504_ (.A(_2436_),
    .B(_2452_),
    .X(_0469_));
 sky130_fd_sc_hd__buf_4 _3505_ (.A(_2450_),
    .X(_2453_));
 sky130_fd_sc_hd__and2_0 _3506_ (.A(_2437_),
    .B(_2453_),
    .X(_0470_));
 sky130_fd_sc_hd__and2_0 _3507_ (.A(_2439_),
    .B(_2453_),
    .X(_0471_));
 sky130_fd_sc_hd__and2_0 _3508_ (.A(_2440_),
    .B(_2453_),
    .X(_0472_));
 sky130_fd_sc_hd__and2_0 _3509_ (.A(_2441_),
    .B(_2453_),
    .X(_0473_));
 sky130_fd_sc_hd__and2_0 _3510_ (.A(_2442_),
    .B(_2453_),
    .X(_0474_));
 sky130_fd_sc_hd__and2_0 _3511_ (.A(_2443_),
    .B(_2453_),
    .X(_0475_));
 sky130_fd_sc_hd__and2_0 _3512_ (.A(_2444_),
    .B(_2453_),
    .X(_0476_));
 sky130_fd_sc_hd__and2_0 _3513_ (.A(_2445_),
    .B(_2453_),
    .X(_0477_));
 sky130_fd_sc_hd__and2_0 _3514_ (.A(_2446_),
    .B(_2453_),
    .X(_0478_));
 sky130_fd_sc_hd__and2_0 _3515_ (.A(_2447_),
    .B(_2453_),
    .X(_0479_));
 sky130_fd_sc_hd__and2_0 _3516_ (.A(_2448_),
    .B(_2450_),
    .X(_0480_));
 sky130_fd_sc_hd__and2_0 _3517_ (.A(_2449_),
    .B(_2450_),
    .X(_0481_));
 sky130_fd_sc_hd__nor2_4 _3518_ (.A(_1127_),
    .B(_1142_),
    .Y(_2454_));
 sky130_fd_sc_hd__buf_2 _3519_ (.A(_2454_),
    .X(_2455_));
 sky130_fd_sc_hd__and2_0 _3520_ (.A(_2414_),
    .B(_2455_),
    .X(_0482_));
 sky130_fd_sc_hd__and2_0 _3521_ (.A(_2417_),
    .B(_2455_),
    .X(_0483_));
 sky130_fd_sc_hd__and2_0 _3522_ (.A(_2418_),
    .B(_2455_),
    .X(_0484_));
 sky130_fd_sc_hd__and2_0 _3523_ (.A(_2419_),
    .B(_2455_),
    .X(_0485_));
 sky130_fd_sc_hd__and2_0 _3524_ (.A(_2420_),
    .B(_2455_),
    .X(_0486_));
 sky130_fd_sc_hd__and2_0 _3525_ (.A(_2421_),
    .B(_2455_),
    .X(_0487_));
 sky130_fd_sc_hd__and2_0 _3526_ (.A(_2422_),
    .B(_2455_),
    .X(_0488_));
 sky130_fd_sc_hd__and2_0 _3527_ (.A(_2423_),
    .B(_2455_),
    .X(_0489_));
 sky130_fd_sc_hd__and2_0 _3528_ (.A(_2424_),
    .B(_2455_),
    .X(_0490_));
 sky130_fd_sc_hd__and2_0 _3529_ (.A(_2425_),
    .B(_2455_),
    .X(_0491_));
 sky130_fd_sc_hd__buf_2 _3530_ (.A(_2454_),
    .X(_2456_));
 sky130_fd_sc_hd__and2_0 _3531_ (.A(_2426_),
    .B(_2456_),
    .X(_0492_));
 sky130_fd_sc_hd__and2_0 _3532_ (.A(_2428_),
    .B(_2456_),
    .X(_0493_));
 sky130_fd_sc_hd__and2_0 _3533_ (.A(_2429_),
    .B(_2456_),
    .X(_0494_));
 sky130_fd_sc_hd__and2_0 _3534_ (.A(_2430_),
    .B(_2456_),
    .X(_0495_));
 sky130_fd_sc_hd__and2_0 _3535_ (.A(_2431_),
    .B(_2456_),
    .X(_0496_));
 sky130_fd_sc_hd__and2_0 _3536_ (.A(_2432_),
    .B(_2456_),
    .X(_0497_));
 sky130_fd_sc_hd__and2_0 _3537_ (.A(_2433_),
    .B(_2456_),
    .X(_0498_));
 sky130_fd_sc_hd__and2_0 _3538_ (.A(_2434_),
    .B(_2456_),
    .X(_0499_));
 sky130_fd_sc_hd__and2_0 _3539_ (.A(_2435_),
    .B(_2456_),
    .X(_0500_));
 sky130_fd_sc_hd__and2_0 _3540_ (.A(_2436_),
    .B(_2456_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_2 _3541_ (.A(_2454_),
    .X(_2457_));
 sky130_fd_sc_hd__and2_0 _3542_ (.A(_2437_),
    .B(_2457_),
    .X(_0502_));
 sky130_fd_sc_hd__and2_0 _3543_ (.A(_2439_),
    .B(_2457_),
    .X(_0503_));
 sky130_fd_sc_hd__and2_0 _3544_ (.A(_2440_),
    .B(_2457_),
    .X(_0504_));
 sky130_fd_sc_hd__and2_0 _3545_ (.A(_2441_),
    .B(_2457_),
    .X(_0505_));
 sky130_fd_sc_hd__and2_0 _3546_ (.A(_2442_),
    .B(_2457_),
    .X(_0506_));
 sky130_fd_sc_hd__and2_0 _3547_ (.A(_2443_),
    .B(_2457_),
    .X(_0507_));
 sky130_fd_sc_hd__and2_0 _3548_ (.A(_2444_),
    .B(_2457_),
    .X(_0508_));
 sky130_fd_sc_hd__and2_0 _3549_ (.A(_2445_),
    .B(_2457_),
    .X(_0509_));
 sky130_fd_sc_hd__and2_0 _3550_ (.A(_2446_),
    .B(_2457_),
    .X(_0510_));
 sky130_fd_sc_hd__and2_0 _3551_ (.A(_2447_),
    .B(_2457_),
    .X(_0511_));
 sky130_fd_sc_hd__and2_0 _3552_ (.A(_2448_),
    .B(_2454_),
    .X(_0512_));
 sky130_fd_sc_hd__and2_0 _3553_ (.A(_2449_),
    .B(_2454_),
    .X(_0513_));
 sky130_fd_sc_hd__nor2_2 _3554_ (.A(_1137_),
    .B(_1142_),
    .Y(_2458_));
 sky130_fd_sc_hd__buf_2 _3555_ (.A(_2458_),
    .X(_2459_));
 sky130_fd_sc_hd__and2_0 _3556_ (.A(_2414_),
    .B(_2459_),
    .X(_0514_));
 sky130_fd_sc_hd__and2_0 _3557_ (.A(_2417_),
    .B(_2459_),
    .X(_0515_));
 sky130_fd_sc_hd__and2_0 _3558_ (.A(_2418_),
    .B(_2459_),
    .X(_0516_));
 sky130_fd_sc_hd__and2_0 _3559_ (.A(_2419_),
    .B(_2459_),
    .X(_0517_));
 sky130_fd_sc_hd__and2_0 _3560_ (.A(_2420_),
    .B(_2459_),
    .X(_0518_));
 sky130_fd_sc_hd__and2_0 _3561_ (.A(_2421_),
    .B(_2459_),
    .X(_0519_));
 sky130_fd_sc_hd__and2_0 _3562_ (.A(_2422_),
    .B(_2459_),
    .X(_0520_));
 sky130_fd_sc_hd__and2_0 _3563_ (.A(_2423_),
    .B(_2459_),
    .X(_0521_));
 sky130_fd_sc_hd__and2_0 _3564_ (.A(_2424_),
    .B(_2459_),
    .X(_0522_));
 sky130_fd_sc_hd__and2_0 _3565_ (.A(_2425_),
    .B(_2459_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_4 _3566_ (.A(_2458_),
    .X(_2460_));
 sky130_fd_sc_hd__and2_0 _3567_ (.A(_2426_),
    .B(_2460_),
    .X(_0524_));
 sky130_fd_sc_hd__and2_0 _3568_ (.A(_2428_),
    .B(_2460_),
    .X(_0525_));
 sky130_fd_sc_hd__and2_0 _3569_ (.A(_2429_),
    .B(_2460_),
    .X(_0526_));
 sky130_fd_sc_hd__and2_0 _3570_ (.A(_2430_),
    .B(_2460_),
    .X(_0527_));
 sky130_fd_sc_hd__and2_0 _3571_ (.A(_2431_),
    .B(_2460_),
    .X(_0528_));
 sky130_fd_sc_hd__and2_0 _3572_ (.A(_2432_),
    .B(_2460_),
    .X(_0529_));
 sky130_fd_sc_hd__and2_0 _3573_ (.A(_2433_),
    .B(_2460_),
    .X(_0530_));
 sky130_fd_sc_hd__and2_0 _3574_ (.A(_2434_),
    .B(_2460_),
    .X(_0531_));
 sky130_fd_sc_hd__and2_0 _3575_ (.A(_2435_),
    .B(_2460_),
    .X(_0532_));
 sky130_fd_sc_hd__and2_0 _3576_ (.A(_2436_),
    .B(_2460_),
    .X(_0533_));
 sky130_fd_sc_hd__buf_2 _3577_ (.A(_2458_),
    .X(_2461_));
 sky130_fd_sc_hd__and2_0 _3578_ (.A(_2437_),
    .B(_2461_),
    .X(_0534_));
 sky130_fd_sc_hd__and2_0 _3579_ (.A(_2439_),
    .B(_2461_),
    .X(_0535_));
 sky130_fd_sc_hd__and2_0 _3580_ (.A(_2440_),
    .B(_2461_),
    .X(_0536_));
 sky130_fd_sc_hd__and2_0 _3581_ (.A(_2441_),
    .B(_2461_),
    .X(_0537_));
 sky130_fd_sc_hd__and2_0 _3582_ (.A(_2442_),
    .B(_2461_),
    .X(_0538_));
 sky130_fd_sc_hd__and2_0 _3583_ (.A(_2443_),
    .B(_2461_),
    .X(_0539_));
 sky130_fd_sc_hd__and2_0 _3584_ (.A(_2444_),
    .B(_2461_),
    .X(_0540_));
 sky130_fd_sc_hd__and2_0 _3585_ (.A(_2445_),
    .B(_2461_),
    .X(_0541_));
 sky130_fd_sc_hd__and2_0 _3586_ (.A(_2446_),
    .B(_2461_),
    .X(_0542_));
 sky130_fd_sc_hd__and2_0 _3587_ (.A(_2447_),
    .B(_2461_),
    .X(_0543_));
 sky130_fd_sc_hd__and2_0 _3588_ (.A(_2448_),
    .B(_2458_),
    .X(_0544_));
 sky130_fd_sc_hd__and2_0 _3589_ (.A(_2449_),
    .B(_2458_),
    .X(_0545_));
 sky130_fd_sc_hd__nor2_4 _3590_ (.A(_1132_),
    .B(_1142_),
    .Y(_2462_));
 sky130_fd_sc_hd__clkbuf_4 _3591_ (.A(_2462_),
    .X(_2463_));
 sky130_fd_sc_hd__and2_0 _3592_ (.A(_2414_),
    .B(_2463_),
    .X(_0546_));
 sky130_fd_sc_hd__and2_0 _3593_ (.A(_2417_),
    .B(_2463_),
    .X(_0547_));
 sky130_fd_sc_hd__and2_0 _3594_ (.A(_2418_),
    .B(_2463_),
    .X(_0548_));
 sky130_fd_sc_hd__and2_0 _3595_ (.A(_2419_),
    .B(_2463_),
    .X(_0549_));
 sky130_fd_sc_hd__and2_0 _3596_ (.A(_2420_),
    .B(_2463_),
    .X(_0550_));
 sky130_fd_sc_hd__and2_0 _3597_ (.A(_2421_),
    .B(_2463_),
    .X(_0551_));
 sky130_fd_sc_hd__and2_0 _3598_ (.A(_2422_),
    .B(_2463_),
    .X(_0552_));
 sky130_fd_sc_hd__and2_0 _3599_ (.A(_2423_),
    .B(_2463_),
    .X(_0553_));
 sky130_fd_sc_hd__and2_0 _3600_ (.A(_2424_),
    .B(_2463_),
    .X(_0554_));
 sky130_fd_sc_hd__and2_0 _3601_ (.A(_2425_),
    .B(_2463_),
    .X(_0555_));
 sky130_fd_sc_hd__clkbuf_4 _3602_ (.A(_2462_),
    .X(_2464_));
 sky130_fd_sc_hd__and2_0 _3603_ (.A(_2426_),
    .B(_2464_),
    .X(_0556_));
 sky130_fd_sc_hd__and2_0 _3604_ (.A(_2428_),
    .B(_2464_),
    .X(_0557_));
 sky130_fd_sc_hd__and2_0 _3605_ (.A(_2429_),
    .B(_2464_),
    .X(_0558_));
 sky130_fd_sc_hd__and2_0 _3606_ (.A(_2430_),
    .B(_2464_),
    .X(_0559_));
 sky130_fd_sc_hd__and2_0 _3607_ (.A(_2431_),
    .B(_2464_),
    .X(_0560_));
 sky130_fd_sc_hd__and2_0 _3608_ (.A(_2432_),
    .B(_2464_),
    .X(_0561_));
 sky130_fd_sc_hd__and2_0 _3609_ (.A(_2433_),
    .B(_2464_),
    .X(_0562_));
 sky130_fd_sc_hd__and2_0 _3610_ (.A(_2434_),
    .B(_2464_),
    .X(_0563_));
 sky130_fd_sc_hd__and2_0 _3611_ (.A(_2435_),
    .B(_2464_),
    .X(_0564_));
 sky130_fd_sc_hd__and2_0 _3612_ (.A(_2436_),
    .B(_2464_),
    .X(_0565_));
 sky130_fd_sc_hd__buf_2 _3613_ (.A(_2462_),
    .X(_2465_));
 sky130_fd_sc_hd__and2_0 _3614_ (.A(_2437_),
    .B(_2465_),
    .X(_0566_));
 sky130_fd_sc_hd__and2_0 _3615_ (.A(_2439_),
    .B(_2465_),
    .X(_0567_));
 sky130_fd_sc_hd__and2_0 _3616_ (.A(_2440_),
    .B(_2465_),
    .X(_0568_));
 sky130_fd_sc_hd__and2_0 _3617_ (.A(_2441_),
    .B(_2465_),
    .X(_0569_));
 sky130_fd_sc_hd__and2_0 _3618_ (.A(_2442_),
    .B(_2465_),
    .X(_0570_));
 sky130_fd_sc_hd__and2_0 _3619_ (.A(_2443_),
    .B(_2465_),
    .X(_0571_));
 sky130_fd_sc_hd__and2_0 _3620_ (.A(_2444_),
    .B(_2465_),
    .X(_0572_));
 sky130_fd_sc_hd__and2_0 _3621_ (.A(_2445_),
    .B(_2465_),
    .X(_0573_));
 sky130_fd_sc_hd__and2_0 _3622_ (.A(_2446_),
    .B(_2465_),
    .X(_0574_));
 sky130_fd_sc_hd__and2_0 _3623_ (.A(_2447_),
    .B(_2465_),
    .X(_0575_));
 sky130_fd_sc_hd__and2_0 _3624_ (.A(_2448_),
    .B(_2462_),
    .X(_0576_));
 sky130_fd_sc_hd__and2_0 _3625_ (.A(_2449_),
    .B(_2462_),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_2 _3626_ (.A(_1134_),
    .B(_1142_),
    .Y(_2466_));
 sky130_fd_sc_hd__buf_2 _3627_ (.A(_2466_),
    .X(_2467_));
 sky130_fd_sc_hd__and2_0 _3628_ (.A(_2414_),
    .B(_2467_),
    .X(_0578_));
 sky130_fd_sc_hd__and2_0 _3629_ (.A(_2417_),
    .B(_2467_),
    .X(_0579_));
 sky130_fd_sc_hd__and2_0 _3630_ (.A(_2418_),
    .B(_2467_),
    .X(_0580_));
 sky130_fd_sc_hd__and2_0 _3631_ (.A(_2419_),
    .B(_2467_),
    .X(_0581_));
 sky130_fd_sc_hd__and2_0 _3632_ (.A(_2420_),
    .B(_2467_),
    .X(_0582_));
 sky130_fd_sc_hd__and2_0 _3633_ (.A(_2421_),
    .B(_2467_),
    .X(_0583_));
 sky130_fd_sc_hd__and2_0 _3634_ (.A(_2422_),
    .B(_2467_),
    .X(_0584_));
 sky130_fd_sc_hd__and2_0 _3635_ (.A(_2423_),
    .B(_2467_),
    .X(_0585_));
 sky130_fd_sc_hd__and2_0 _3636_ (.A(_2424_),
    .B(_2467_),
    .X(_0586_));
 sky130_fd_sc_hd__and2_0 _3637_ (.A(_2425_),
    .B(_2467_),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_4 _3638_ (.A(_2466_),
    .X(_2468_));
 sky130_fd_sc_hd__and2_0 _3639_ (.A(_2426_),
    .B(_2468_),
    .X(_0588_));
 sky130_fd_sc_hd__and2_0 _3640_ (.A(_2428_),
    .B(_2468_),
    .X(_0589_));
 sky130_fd_sc_hd__and2_0 _3641_ (.A(_2429_),
    .B(_2468_),
    .X(_0590_));
 sky130_fd_sc_hd__and2_0 _3642_ (.A(_2430_),
    .B(_2468_),
    .X(_0591_));
 sky130_fd_sc_hd__and2_0 _3643_ (.A(_2431_),
    .B(_2468_),
    .X(_0592_));
 sky130_fd_sc_hd__and2_0 _3644_ (.A(_2432_),
    .B(_2468_),
    .X(_0593_));
 sky130_fd_sc_hd__and2_0 _3645_ (.A(_2433_),
    .B(_2468_),
    .X(_0594_));
 sky130_fd_sc_hd__and2_0 _3646_ (.A(_2434_),
    .B(_2468_),
    .X(_0595_));
 sky130_fd_sc_hd__and2_0 _3647_ (.A(_2435_),
    .B(_2468_),
    .X(_0596_));
 sky130_fd_sc_hd__and2_0 _3648_ (.A(_2436_),
    .B(_2468_),
    .X(_0597_));
 sky130_fd_sc_hd__clkbuf_4 _3649_ (.A(_2466_),
    .X(_2469_));
 sky130_fd_sc_hd__and2_0 _3650_ (.A(_2437_),
    .B(_2469_),
    .X(_0598_));
 sky130_fd_sc_hd__and2_0 _3651_ (.A(_2439_),
    .B(_2469_),
    .X(_0599_));
 sky130_fd_sc_hd__and2_0 _3652_ (.A(_2440_),
    .B(_2469_),
    .X(_0600_));
 sky130_fd_sc_hd__and2_0 _3653_ (.A(_2441_),
    .B(_2469_),
    .X(_0601_));
 sky130_fd_sc_hd__and2_0 _3654_ (.A(_2442_),
    .B(_2469_),
    .X(_0602_));
 sky130_fd_sc_hd__and2_0 _3655_ (.A(_2443_),
    .B(_2469_),
    .X(_0603_));
 sky130_fd_sc_hd__and2_0 _3656_ (.A(_2444_),
    .B(_2469_),
    .X(_0604_));
 sky130_fd_sc_hd__and2_0 _3657_ (.A(_2445_),
    .B(_2469_),
    .X(_0605_));
 sky130_fd_sc_hd__and2_0 _3658_ (.A(_2446_),
    .B(_2469_),
    .X(_0606_));
 sky130_fd_sc_hd__and2_0 _3659_ (.A(_2447_),
    .B(_2469_),
    .X(_0607_));
 sky130_fd_sc_hd__and2_0 _3660_ (.A(_2448_),
    .B(_2466_),
    .X(_0608_));
 sky130_fd_sc_hd__and2_0 _3661_ (.A(_2449_),
    .B(_2466_),
    .X(_0609_));
 sky130_fd_sc_hd__nor2_4 _3662_ (.A(_1127_),
    .B(_1143_),
    .Y(_2470_));
 sky130_fd_sc_hd__clkbuf_4 _3663_ (.A(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__and2_0 _3664_ (.A(_2414_),
    .B(_2471_),
    .X(_0610_));
 sky130_fd_sc_hd__and2_0 _3665_ (.A(_2417_),
    .B(_2471_),
    .X(_0611_));
 sky130_fd_sc_hd__and2_0 _3666_ (.A(_2418_),
    .B(_2471_),
    .X(_0612_));
 sky130_fd_sc_hd__and2_0 _3667_ (.A(_2419_),
    .B(_2471_),
    .X(_0613_));
 sky130_fd_sc_hd__and2_0 _3668_ (.A(_2420_),
    .B(_2471_),
    .X(_0614_));
 sky130_fd_sc_hd__and2_0 _3669_ (.A(_2421_),
    .B(_2471_),
    .X(_0615_));
 sky130_fd_sc_hd__and2_0 _3670_ (.A(_2422_),
    .B(_2471_),
    .X(_0616_));
 sky130_fd_sc_hd__and2_0 _3671_ (.A(_2423_),
    .B(_2471_),
    .X(_0617_));
 sky130_fd_sc_hd__and2_0 _3672_ (.A(_2424_),
    .B(_2471_),
    .X(_0618_));
 sky130_fd_sc_hd__and2_0 _3673_ (.A(_2425_),
    .B(_2471_),
    .X(_0619_));
 sky130_fd_sc_hd__clkbuf_4 _3674_ (.A(_2470_),
    .X(_2472_));
 sky130_fd_sc_hd__and2_0 _3675_ (.A(_2426_),
    .B(_2472_),
    .X(_0620_));
 sky130_fd_sc_hd__and2_0 _3676_ (.A(_2428_),
    .B(_2472_),
    .X(_0621_));
 sky130_fd_sc_hd__and2_0 _3677_ (.A(_2429_),
    .B(_2472_),
    .X(_0622_));
 sky130_fd_sc_hd__and2_0 _3678_ (.A(_2430_),
    .B(_2472_),
    .X(_0623_));
 sky130_fd_sc_hd__and2_0 _3679_ (.A(_2431_),
    .B(_2472_),
    .X(_0624_));
 sky130_fd_sc_hd__and2_0 _3680_ (.A(_2432_),
    .B(_2472_),
    .X(_0625_));
 sky130_fd_sc_hd__and2_0 _3681_ (.A(_2433_),
    .B(_2472_),
    .X(_0626_));
 sky130_fd_sc_hd__and2_0 _3682_ (.A(_2434_),
    .B(_2472_),
    .X(_0627_));
 sky130_fd_sc_hd__and2_0 _3683_ (.A(_2435_),
    .B(_2472_),
    .X(_0628_));
 sky130_fd_sc_hd__and2_0 _3684_ (.A(_2436_),
    .B(_2472_),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_4 _3685_ (.A(_2470_),
    .X(_2473_));
 sky130_fd_sc_hd__and2_0 _3686_ (.A(_2437_),
    .B(_2473_),
    .X(_0630_));
 sky130_fd_sc_hd__and2_0 _3687_ (.A(_2439_),
    .B(_2473_),
    .X(_0631_));
 sky130_fd_sc_hd__and2_0 _3688_ (.A(_2440_),
    .B(_2473_),
    .X(_0632_));
 sky130_fd_sc_hd__and2_0 _3689_ (.A(_2441_),
    .B(_2473_),
    .X(_0633_));
 sky130_fd_sc_hd__and2_0 _3690_ (.A(_2442_),
    .B(_2473_),
    .X(_0634_));
 sky130_fd_sc_hd__and2_0 _3691_ (.A(_2443_),
    .B(_2473_),
    .X(_0635_));
 sky130_fd_sc_hd__and2_0 _3692_ (.A(_2444_),
    .B(_2473_),
    .X(_0636_));
 sky130_fd_sc_hd__and2_0 _3693_ (.A(_2445_),
    .B(_2473_),
    .X(_0637_));
 sky130_fd_sc_hd__and2_0 _3694_ (.A(_2446_),
    .B(_2473_),
    .X(_0638_));
 sky130_fd_sc_hd__and2_0 _3695_ (.A(_2447_),
    .B(_2473_),
    .X(_0639_));
 sky130_fd_sc_hd__and2_0 _3696_ (.A(_2448_),
    .B(_2470_),
    .X(_0640_));
 sky130_fd_sc_hd__and2_0 _3697_ (.A(_2449_),
    .B(_2470_),
    .X(_0641_));
 sky130_fd_sc_hd__nor2_4 _3698_ (.A(_1137_),
    .B(_1143_),
    .Y(_2474_));
 sky130_fd_sc_hd__buf_4 _3699_ (.A(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__and2_0 _3700_ (.A(_2414_),
    .B(_2475_),
    .X(_0642_));
 sky130_fd_sc_hd__and2_0 _3701_ (.A(_2417_),
    .B(_2475_),
    .X(_0643_));
 sky130_fd_sc_hd__and2_0 _3702_ (.A(_2418_),
    .B(_2475_),
    .X(_0644_));
 sky130_fd_sc_hd__and2_0 _3703_ (.A(_2419_),
    .B(_2475_),
    .X(_0645_));
 sky130_fd_sc_hd__and2_0 _3704_ (.A(_2420_),
    .B(_2475_),
    .X(_0646_));
 sky130_fd_sc_hd__and2_0 _3705_ (.A(_2421_),
    .B(_2475_),
    .X(_0647_));
 sky130_fd_sc_hd__and2_0 _3706_ (.A(_2422_),
    .B(_2475_),
    .X(_0648_));
 sky130_fd_sc_hd__and2_0 _3707_ (.A(_2423_),
    .B(_2475_),
    .X(_0649_));
 sky130_fd_sc_hd__and2_0 _3708_ (.A(_2424_),
    .B(_2475_),
    .X(_0650_));
 sky130_fd_sc_hd__and2_0 _3709_ (.A(_2425_),
    .B(_2475_),
    .X(_0651_));
 sky130_fd_sc_hd__buf_4 _3710_ (.A(_2474_),
    .X(_2476_));
 sky130_fd_sc_hd__and2_0 _3711_ (.A(_2426_),
    .B(_2476_),
    .X(_0652_));
 sky130_fd_sc_hd__and2_0 _3712_ (.A(_2428_),
    .B(_2476_),
    .X(_0653_));
 sky130_fd_sc_hd__and2_0 _3713_ (.A(_2429_),
    .B(_2476_),
    .X(_0654_));
 sky130_fd_sc_hd__and2_0 _3714_ (.A(_2430_),
    .B(_2476_),
    .X(_0655_));
 sky130_fd_sc_hd__and2_0 _3715_ (.A(_2431_),
    .B(_2476_),
    .X(_0656_));
 sky130_fd_sc_hd__and2_0 _3716_ (.A(_2432_),
    .B(_2476_),
    .X(_0657_));
 sky130_fd_sc_hd__and2_0 _3717_ (.A(_2433_),
    .B(_2476_),
    .X(_0658_));
 sky130_fd_sc_hd__and2_0 _3718_ (.A(_2434_),
    .B(_2476_),
    .X(_0659_));
 sky130_fd_sc_hd__and2_0 _3719_ (.A(_2435_),
    .B(_2476_),
    .X(_0660_));
 sky130_fd_sc_hd__and2_0 _3720_ (.A(_2436_),
    .B(_2476_),
    .X(_0661_));
 sky130_fd_sc_hd__buf_4 _3721_ (.A(_2474_),
    .X(_2477_));
 sky130_fd_sc_hd__and2_0 _3722_ (.A(_2437_),
    .B(_2477_),
    .X(_0662_));
 sky130_fd_sc_hd__and2_0 _3723_ (.A(_2439_),
    .B(_2477_),
    .X(_0663_));
 sky130_fd_sc_hd__and2_0 _3724_ (.A(_2440_),
    .B(_2477_),
    .X(_0664_));
 sky130_fd_sc_hd__and2_0 _3725_ (.A(_2441_),
    .B(_2477_),
    .X(_0665_));
 sky130_fd_sc_hd__and2_0 _3726_ (.A(_2442_),
    .B(_2477_),
    .X(_0666_));
 sky130_fd_sc_hd__and2_0 _3727_ (.A(_2443_),
    .B(_2477_),
    .X(_0667_));
 sky130_fd_sc_hd__and2_0 _3728_ (.A(_2444_),
    .B(_2477_),
    .X(_0668_));
 sky130_fd_sc_hd__and2_0 _3729_ (.A(_2445_),
    .B(_2477_),
    .X(_0669_));
 sky130_fd_sc_hd__and2_0 _3730_ (.A(_2446_),
    .B(_2477_),
    .X(_0670_));
 sky130_fd_sc_hd__and2_0 _3731_ (.A(_2447_),
    .B(_2477_),
    .X(_0671_));
 sky130_fd_sc_hd__and2_0 _3732_ (.A(_2448_),
    .B(_2474_),
    .X(_0672_));
 sky130_fd_sc_hd__and2_0 _3733_ (.A(_2449_),
    .B(_2474_),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_2 _3734_ (.A(_1132_),
    .B(_1143_),
    .Y(_2478_));
 sky130_fd_sc_hd__buf_4 _3735_ (.A(_2478_),
    .X(_2479_));
 sky130_fd_sc_hd__and2_0 _3736_ (.A(_2414_),
    .B(_2479_),
    .X(_0674_));
 sky130_fd_sc_hd__and2_0 _3737_ (.A(_2417_),
    .B(_2479_),
    .X(_0675_));
 sky130_fd_sc_hd__and2_0 _3738_ (.A(_2418_),
    .B(_2479_),
    .X(_0676_));
 sky130_fd_sc_hd__and2_0 _3739_ (.A(_2419_),
    .B(_2479_),
    .X(_0677_));
 sky130_fd_sc_hd__and2_0 _3740_ (.A(_2420_),
    .B(_2479_),
    .X(_0678_));
 sky130_fd_sc_hd__and2_0 _3741_ (.A(_2421_),
    .B(_2479_),
    .X(_0679_));
 sky130_fd_sc_hd__and2_0 _3742_ (.A(_2422_),
    .B(_2479_),
    .X(_0680_));
 sky130_fd_sc_hd__and2_0 _3743_ (.A(_2423_),
    .B(_2479_),
    .X(_0681_));
 sky130_fd_sc_hd__and2_0 _3744_ (.A(_2424_),
    .B(_2479_),
    .X(_0682_));
 sky130_fd_sc_hd__and2_0 _3745_ (.A(_2425_),
    .B(_2479_),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_4 _3746_ (.A(_2478_),
    .X(_2480_));
 sky130_fd_sc_hd__and2_0 _3747_ (.A(_2426_),
    .B(_2480_),
    .X(_0684_));
 sky130_fd_sc_hd__and2_0 _3748_ (.A(_2428_),
    .B(_2480_),
    .X(_0685_));
 sky130_fd_sc_hd__and2_0 _3749_ (.A(_2429_),
    .B(_2480_),
    .X(_0686_));
 sky130_fd_sc_hd__and2_0 _3750_ (.A(_2430_),
    .B(_2480_),
    .X(_0687_));
 sky130_fd_sc_hd__and2_0 _3751_ (.A(_2431_),
    .B(_2480_),
    .X(_0688_));
 sky130_fd_sc_hd__and2_0 _3752_ (.A(_2432_),
    .B(_2480_),
    .X(_0689_));
 sky130_fd_sc_hd__and2_0 _3753_ (.A(_2433_),
    .B(_2480_),
    .X(_0690_));
 sky130_fd_sc_hd__and2_0 _3754_ (.A(_2434_),
    .B(_2480_),
    .X(_0691_));
 sky130_fd_sc_hd__and2_0 _3755_ (.A(_2435_),
    .B(_2480_),
    .X(_0692_));
 sky130_fd_sc_hd__and2_0 _3756_ (.A(_2436_),
    .B(_2480_),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_4 _3757_ (.A(_2478_),
    .X(_2481_));
 sky130_fd_sc_hd__and2_0 _3758_ (.A(_2437_),
    .B(_2481_),
    .X(_0694_));
 sky130_fd_sc_hd__and2_0 _3759_ (.A(_2439_),
    .B(_2481_),
    .X(_0695_));
 sky130_fd_sc_hd__and2_0 _3760_ (.A(_2440_),
    .B(_2481_),
    .X(_0696_));
 sky130_fd_sc_hd__and2_0 _3761_ (.A(_2441_),
    .B(_2481_),
    .X(_0697_));
 sky130_fd_sc_hd__and2_0 _3762_ (.A(_2442_),
    .B(_2481_),
    .X(_0698_));
 sky130_fd_sc_hd__and2_0 _3763_ (.A(_2443_),
    .B(_2481_),
    .X(_0699_));
 sky130_fd_sc_hd__and2_0 _3764_ (.A(_2444_),
    .B(_2481_),
    .X(_0700_));
 sky130_fd_sc_hd__and2_0 _3765_ (.A(_2445_),
    .B(_2481_),
    .X(_0701_));
 sky130_fd_sc_hd__and2_0 _3766_ (.A(_2446_),
    .B(_2481_),
    .X(_0702_));
 sky130_fd_sc_hd__and2_0 _3767_ (.A(_2447_),
    .B(_2481_),
    .X(_0703_));
 sky130_fd_sc_hd__and2_0 _3768_ (.A(_2448_),
    .B(_2478_),
    .X(_0704_));
 sky130_fd_sc_hd__and2_0 _3769_ (.A(_2449_),
    .B(_2478_),
    .X(_0705_));
 sky130_fd_sc_hd__nor2_4 _3770_ (.A(_1134_),
    .B(_1143_),
    .Y(_2482_));
 sky130_fd_sc_hd__buf_4 _3771_ (.A(_2482_),
    .X(_2483_));
 sky130_fd_sc_hd__and2_0 _3772_ (.A(_2414_),
    .B(_2483_),
    .X(_0706_));
 sky130_fd_sc_hd__and2_0 _3773_ (.A(_2417_),
    .B(_2483_),
    .X(_0707_));
 sky130_fd_sc_hd__and2_0 _3774_ (.A(_2418_),
    .B(_2483_),
    .X(_0708_));
 sky130_fd_sc_hd__and2_0 _3775_ (.A(_2419_),
    .B(_2483_),
    .X(_0709_));
 sky130_fd_sc_hd__and2_0 _3776_ (.A(_2420_),
    .B(_2483_),
    .X(_0710_));
 sky130_fd_sc_hd__and2_0 _3777_ (.A(_2421_),
    .B(_2483_),
    .X(_0711_));
 sky130_fd_sc_hd__and2_0 _3778_ (.A(_2422_),
    .B(_2483_),
    .X(_0712_));
 sky130_fd_sc_hd__and2_0 _3779_ (.A(_2423_),
    .B(_2483_),
    .X(_0713_));
 sky130_fd_sc_hd__and2_0 _3780_ (.A(_2424_),
    .B(_2483_),
    .X(_0714_));
 sky130_fd_sc_hd__and2_0 _3781_ (.A(_2425_),
    .B(_2483_),
    .X(_0715_));
 sky130_fd_sc_hd__buf_4 _3782_ (.A(_2482_),
    .X(_2484_));
 sky130_fd_sc_hd__and2_0 _3783_ (.A(_2426_),
    .B(_2484_),
    .X(_0716_));
 sky130_fd_sc_hd__and2_0 _3784_ (.A(_2428_),
    .B(_2484_),
    .X(_0717_));
 sky130_fd_sc_hd__and2_0 _3785_ (.A(_2429_),
    .B(_2484_),
    .X(_0718_));
 sky130_fd_sc_hd__and2_0 _3786_ (.A(_2430_),
    .B(_2484_),
    .X(_0719_));
 sky130_fd_sc_hd__and2_0 _3787_ (.A(_2431_),
    .B(_2484_),
    .X(_0720_));
 sky130_fd_sc_hd__and2_0 _3788_ (.A(_2432_),
    .B(_2484_),
    .X(_0721_));
 sky130_fd_sc_hd__and2_0 _3789_ (.A(_2433_),
    .B(_2484_),
    .X(_0722_));
 sky130_fd_sc_hd__and2_0 _3790_ (.A(_2434_),
    .B(_2484_),
    .X(_0723_));
 sky130_fd_sc_hd__and2_0 _3791_ (.A(_2435_),
    .B(_2484_),
    .X(_0724_));
 sky130_fd_sc_hd__and2_0 _3792_ (.A(_2436_),
    .B(_2484_),
    .X(_0725_));
 sky130_fd_sc_hd__buf_4 _3793_ (.A(_2482_),
    .X(_2485_));
 sky130_fd_sc_hd__and2_0 _3794_ (.A(_2437_),
    .B(_2485_),
    .X(_0726_));
 sky130_fd_sc_hd__and2_0 _3795_ (.A(_2439_),
    .B(_2485_),
    .X(_0727_));
 sky130_fd_sc_hd__and2_0 _3796_ (.A(_2440_),
    .B(_2485_),
    .X(_0728_));
 sky130_fd_sc_hd__and2_0 _3797_ (.A(_2441_),
    .B(_2485_),
    .X(_0729_));
 sky130_fd_sc_hd__and2_0 _3798_ (.A(_2442_),
    .B(_2485_),
    .X(_0730_));
 sky130_fd_sc_hd__and2_0 _3799_ (.A(_2443_),
    .B(_2485_),
    .X(_0731_));
 sky130_fd_sc_hd__and2_0 _3800_ (.A(_2444_),
    .B(_2485_),
    .X(_0732_));
 sky130_fd_sc_hd__and2_0 _3801_ (.A(_2445_),
    .B(_2485_),
    .X(_0733_));
 sky130_fd_sc_hd__and2_0 _3802_ (.A(_2446_),
    .B(_2485_),
    .X(_0734_));
 sky130_fd_sc_hd__and2_0 _3803_ (.A(_2447_),
    .B(_2485_),
    .X(_0735_));
 sky130_fd_sc_hd__and2_0 _3804_ (.A(_2448_),
    .B(_2482_),
    .X(_0736_));
 sky130_fd_sc_hd__and2_0 _3805_ (.A(_2449_),
    .B(_2482_),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_4 _3806_ (.A(net11),
    .X(_2486_));
 sky130_fd_sc_hd__nor2_2 _3807_ (.A(_1127_),
    .B(_1144_),
    .Y(_2487_));
 sky130_fd_sc_hd__clkbuf_4 _3808_ (.A(_2487_),
    .X(_2488_));
 sky130_fd_sc_hd__and2_0 _3809_ (.A(_2486_),
    .B(_2488_),
    .X(_0738_));
 sky130_fd_sc_hd__buf_2 _3810_ (.A(net12),
    .X(_2489_));
 sky130_fd_sc_hd__and2_0 _3811_ (.A(_2489_),
    .B(_2488_),
    .X(_0739_));
 sky130_fd_sc_hd__clkbuf_4 _3812_ (.A(net13),
    .X(_2490_));
 sky130_fd_sc_hd__and2_0 _3813_ (.A(_2490_),
    .B(_2488_),
    .X(_0740_));
 sky130_fd_sc_hd__buf_4 _3814_ (.A(net14),
    .X(_2491_));
 sky130_fd_sc_hd__and2_0 _3815_ (.A(_2491_),
    .B(_2488_),
    .X(_0741_));
 sky130_fd_sc_hd__clkbuf_4 _3816_ (.A(net15),
    .X(_2492_));
 sky130_fd_sc_hd__and2_0 _3817_ (.A(_2492_),
    .B(_2488_),
    .X(_0742_));
 sky130_fd_sc_hd__buf_4 _3818_ (.A(net16),
    .X(_2493_));
 sky130_fd_sc_hd__and2_0 _3819_ (.A(_2493_),
    .B(_2488_),
    .X(_0743_));
 sky130_fd_sc_hd__buf_4 _3820_ (.A(net17),
    .X(_2494_));
 sky130_fd_sc_hd__and2_0 _3821_ (.A(_2494_),
    .B(_2488_),
    .X(_0744_));
 sky130_fd_sc_hd__clkbuf_4 _3822_ (.A(net18),
    .X(_2495_));
 sky130_fd_sc_hd__and2_0 _3823_ (.A(_2495_),
    .B(_2488_),
    .X(_0745_));
 sky130_fd_sc_hd__buf_4 _3824_ (.A(net19),
    .X(_2496_));
 sky130_fd_sc_hd__and2_0 _3825_ (.A(_2496_),
    .B(_2488_),
    .X(_0746_));
 sky130_fd_sc_hd__clkbuf_4 _3826_ (.A(net20),
    .X(_2497_));
 sky130_fd_sc_hd__and2_0 _3827_ (.A(_2497_),
    .B(_2488_),
    .X(_0747_));
 sky130_fd_sc_hd__buf_4 _3828_ (.A(net21),
    .X(_2498_));
 sky130_fd_sc_hd__clkbuf_4 _3829_ (.A(_2487_),
    .X(_2499_));
 sky130_fd_sc_hd__and2_0 _3830_ (.A(_2498_),
    .B(_2499_),
    .X(_0748_));
 sky130_fd_sc_hd__buf_4 _3831_ (.A(net22),
    .X(_2500_));
 sky130_fd_sc_hd__and2_0 _3832_ (.A(_2500_),
    .B(_2499_),
    .X(_0749_));
 sky130_fd_sc_hd__buf_4 _3833_ (.A(net23),
    .X(_2501_));
 sky130_fd_sc_hd__and2_0 _3834_ (.A(_2501_),
    .B(_2499_),
    .X(_0750_));
 sky130_fd_sc_hd__buf_4 _3835_ (.A(net24),
    .X(_2502_));
 sky130_fd_sc_hd__and2_0 _3836_ (.A(_2502_),
    .B(_2499_),
    .X(_0751_));
 sky130_fd_sc_hd__buf_4 _3837_ (.A(net25),
    .X(_2503_));
 sky130_fd_sc_hd__and2_0 _3838_ (.A(_2503_),
    .B(_2499_),
    .X(_0752_));
 sky130_fd_sc_hd__buf_4 _3839_ (.A(net26),
    .X(_2504_));
 sky130_fd_sc_hd__and2_0 _3840_ (.A(_2504_),
    .B(_2499_),
    .X(_0753_));
 sky130_fd_sc_hd__buf_4 _3841_ (.A(net27),
    .X(_2505_));
 sky130_fd_sc_hd__and2_0 _3842_ (.A(_2505_),
    .B(_2499_),
    .X(_0754_));
 sky130_fd_sc_hd__buf_4 _3843_ (.A(net28),
    .X(_2506_));
 sky130_fd_sc_hd__and2_0 _3844_ (.A(_2506_),
    .B(_2499_),
    .X(_0755_));
 sky130_fd_sc_hd__clkbuf_4 _3845_ (.A(net29),
    .X(_2507_));
 sky130_fd_sc_hd__and2_0 _3846_ (.A(_2507_),
    .B(_2499_),
    .X(_0756_));
 sky130_fd_sc_hd__buf_4 _3847_ (.A(net30),
    .X(_2508_));
 sky130_fd_sc_hd__and2_0 _3848_ (.A(_2508_),
    .B(_2499_),
    .X(_0757_));
 sky130_fd_sc_hd__buf_4 _3849_ (.A(net31),
    .X(_2509_));
 sky130_fd_sc_hd__clkbuf_4 _3850_ (.A(_2487_),
    .X(_2510_));
 sky130_fd_sc_hd__and2_0 _3851_ (.A(_2509_),
    .B(_2510_),
    .X(_0758_));
 sky130_fd_sc_hd__buf_4 _3852_ (.A(net32),
    .X(_2511_));
 sky130_fd_sc_hd__and2_0 _3853_ (.A(_2511_),
    .B(_2510_),
    .X(_0759_));
 sky130_fd_sc_hd__buf_4 _3854_ (.A(net33),
    .X(_2512_));
 sky130_fd_sc_hd__and2_0 _3855_ (.A(_2512_),
    .B(_2510_),
    .X(_0760_));
 sky130_fd_sc_hd__buf_4 _3856_ (.A(net34),
    .X(_2513_));
 sky130_fd_sc_hd__and2_0 _3857_ (.A(_2513_),
    .B(_2510_),
    .X(_0761_));
 sky130_fd_sc_hd__buf_4 _3858_ (.A(net35),
    .X(_2514_));
 sky130_fd_sc_hd__and2_0 _3859_ (.A(_2514_),
    .B(_2510_),
    .X(_0762_));
 sky130_fd_sc_hd__clkbuf_4 _3860_ (.A(net36),
    .X(_2515_));
 sky130_fd_sc_hd__and2_0 _3861_ (.A(_2515_),
    .B(_2510_),
    .X(_0763_));
 sky130_fd_sc_hd__buf_4 _3862_ (.A(net37),
    .X(_2516_));
 sky130_fd_sc_hd__and2_0 _3863_ (.A(_2516_),
    .B(_2510_),
    .X(_0764_));
 sky130_fd_sc_hd__clkbuf_4 _3864_ (.A(net38),
    .X(_2517_));
 sky130_fd_sc_hd__and2_0 _3865_ (.A(_2517_),
    .B(_2510_),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_4 _3866_ (.A(net39),
    .X(_2518_));
 sky130_fd_sc_hd__and2_0 _3867_ (.A(_2518_),
    .B(_2510_),
    .X(_0766_));
 sky130_fd_sc_hd__clkbuf_4 _3868_ (.A(net40),
    .X(_2519_));
 sky130_fd_sc_hd__and2_0 _3869_ (.A(_2519_),
    .B(_2510_),
    .X(_0767_));
 sky130_fd_sc_hd__clkbuf_4 _3870_ (.A(net41),
    .X(_2520_));
 sky130_fd_sc_hd__and2_0 _3871_ (.A(_2520_),
    .B(_2487_),
    .X(_0768_));
 sky130_fd_sc_hd__clkbuf_4 _3872_ (.A(net42),
    .X(_2521_));
 sky130_fd_sc_hd__and2_0 _3873_ (.A(_2521_),
    .B(_2487_),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_2 _3874_ (.A(_1137_),
    .B(_1144_),
    .Y(_2522_));
 sky130_fd_sc_hd__buf_4 _3875_ (.A(_2522_),
    .X(_2523_));
 sky130_fd_sc_hd__and2_0 _3876_ (.A(_2486_),
    .B(_2523_),
    .X(_0770_));
 sky130_fd_sc_hd__and2_0 _3877_ (.A(_2489_),
    .B(_2523_),
    .X(_0771_));
 sky130_fd_sc_hd__and2_0 _3878_ (.A(_2490_),
    .B(_2523_),
    .X(_0772_));
 sky130_fd_sc_hd__and2_0 _3879_ (.A(_2491_),
    .B(_2523_),
    .X(_0773_));
 sky130_fd_sc_hd__and2_0 _3880_ (.A(_2492_),
    .B(_2523_),
    .X(_0774_));
 sky130_fd_sc_hd__and2_0 _3881_ (.A(_2493_),
    .B(_2523_),
    .X(_0775_));
 sky130_fd_sc_hd__and2_0 _3882_ (.A(_2494_),
    .B(_2523_),
    .X(_0776_));
 sky130_fd_sc_hd__and2_0 _3883_ (.A(_2495_),
    .B(_2523_),
    .X(_0777_));
 sky130_fd_sc_hd__and2_0 _3884_ (.A(_2496_),
    .B(_2523_),
    .X(_0778_));
 sky130_fd_sc_hd__and2_0 _3885_ (.A(_2497_),
    .B(_2523_),
    .X(_0779_));
 sky130_fd_sc_hd__buf_4 _3886_ (.A(_2522_),
    .X(_2524_));
 sky130_fd_sc_hd__and2_0 _3887_ (.A(_2498_),
    .B(_2524_),
    .X(_0780_));
 sky130_fd_sc_hd__and2_0 _3888_ (.A(_2500_),
    .B(_2524_),
    .X(_0781_));
 sky130_fd_sc_hd__and2_0 _3889_ (.A(_2501_),
    .B(_2524_),
    .X(_0782_));
 sky130_fd_sc_hd__and2_0 _3890_ (.A(_2502_),
    .B(_2524_),
    .X(_0783_));
 sky130_fd_sc_hd__and2_0 _3891_ (.A(_2503_),
    .B(_2524_),
    .X(_0784_));
 sky130_fd_sc_hd__and2_0 _3892_ (.A(_2504_),
    .B(_2524_),
    .X(_0785_));
 sky130_fd_sc_hd__and2_0 _3893_ (.A(_2505_),
    .B(_2524_),
    .X(_0786_));
 sky130_fd_sc_hd__and2_0 _3894_ (.A(_2506_),
    .B(_2524_),
    .X(_0787_));
 sky130_fd_sc_hd__and2_0 _3895_ (.A(_2507_),
    .B(_2524_),
    .X(_0788_));
 sky130_fd_sc_hd__and2_0 _3896_ (.A(_2508_),
    .B(_2524_),
    .X(_0789_));
 sky130_fd_sc_hd__buf_4 _3897_ (.A(_2522_),
    .X(_2525_));
 sky130_fd_sc_hd__and2_0 _3898_ (.A(_2509_),
    .B(_2525_),
    .X(_0790_));
 sky130_fd_sc_hd__and2_0 _3899_ (.A(_2511_),
    .B(_2525_),
    .X(_0791_));
 sky130_fd_sc_hd__and2_0 _3900_ (.A(_2512_),
    .B(_2525_),
    .X(_0792_));
 sky130_fd_sc_hd__and2_0 _3901_ (.A(_2513_),
    .B(_2525_),
    .X(_0793_));
 sky130_fd_sc_hd__and2_0 _3902_ (.A(_2514_),
    .B(_2525_),
    .X(_0794_));
 sky130_fd_sc_hd__and2_0 _3903_ (.A(_2515_),
    .B(_2525_),
    .X(_0795_));
 sky130_fd_sc_hd__and2_0 _3904_ (.A(_2516_),
    .B(_2525_),
    .X(_0796_));
 sky130_fd_sc_hd__and2_0 _3905_ (.A(_2517_),
    .B(_2525_),
    .X(_0797_));
 sky130_fd_sc_hd__and2_0 _3906_ (.A(_2518_),
    .B(_2525_),
    .X(_0798_));
 sky130_fd_sc_hd__and2_0 _3907_ (.A(_2519_),
    .B(_2525_),
    .X(_0799_));
 sky130_fd_sc_hd__and2_0 _3908_ (.A(_2520_),
    .B(_2522_),
    .X(_0800_));
 sky130_fd_sc_hd__and2_0 _3909_ (.A(_2521_),
    .B(_2522_),
    .X(_0801_));
 sky130_fd_sc_hd__nor2_4 _3910_ (.A(_1124_),
    .B(_1133_),
    .Y(_2526_));
 sky130_fd_sc_hd__buf_4 _3911_ (.A(_2526_),
    .X(_2527_));
 sky130_fd_sc_hd__and2_0 _3912_ (.A(_2486_),
    .B(_2527_),
    .X(_0802_));
 sky130_fd_sc_hd__and2_0 _3913_ (.A(_2489_),
    .B(_2527_),
    .X(_0803_));
 sky130_fd_sc_hd__and2_0 _3914_ (.A(_2490_),
    .B(_2527_),
    .X(_0804_));
 sky130_fd_sc_hd__and2_0 _3915_ (.A(_2491_),
    .B(_2527_),
    .X(_0805_));
 sky130_fd_sc_hd__and2_0 _3916_ (.A(_2492_),
    .B(_2527_),
    .X(_0806_));
 sky130_fd_sc_hd__and2_0 _3917_ (.A(_2493_),
    .B(_2527_),
    .X(_0807_));
 sky130_fd_sc_hd__and2_0 _3918_ (.A(_2494_),
    .B(_2527_),
    .X(_0808_));
 sky130_fd_sc_hd__and2_0 _3919_ (.A(_2495_),
    .B(_2527_),
    .X(_0809_));
 sky130_fd_sc_hd__and2_0 _3920_ (.A(_2496_),
    .B(_2527_),
    .X(_0810_));
 sky130_fd_sc_hd__and2_0 _3921_ (.A(_2497_),
    .B(_2527_),
    .X(_0811_));
 sky130_fd_sc_hd__buf_4 _3922_ (.A(_2526_),
    .X(_2528_));
 sky130_fd_sc_hd__and2_0 _3923_ (.A(_2498_),
    .B(_2528_),
    .X(_0812_));
 sky130_fd_sc_hd__and2_0 _3924_ (.A(_2500_),
    .B(_2528_),
    .X(_0813_));
 sky130_fd_sc_hd__and2_0 _3925_ (.A(_2501_),
    .B(_2528_),
    .X(_0814_));
 sky130_fd_sc_hd__and2_0 _3926_ (.A(_2502_),
    .B(_2528_),
    .X(_0815_));
 sky130_fd_sc_hd__and2_0 _3927_ (.A(_2503_),
    .B(_2528_),
    .X(_0816_));
 sky130_fd_sc_hd__and2_0 _3928_ (.A(_2504_),
    .B(_2528_),
    .X(_0817_));
 sky130_fd_sc_hd__and2_0 _3929_ (.A(_2505_),
    .B(_2528_),
    .X(_0818_));
 sky130_fd_sc_hd__and2_0 _3930_ (.A(_2506_),
    .B(_2528_),
    .X(_0819_));
 sky130_fd_sc_hd__and2_0 _3931_ (.A(_2507_),
    .B(_2528_),
    .X(_0820_));
 sky130_fd_sc_hd__and2_0 _3932_ (.A(_2508_),
    .B(_2528_),
    .X(_0821_));
 sky130_fd_sc_hd__buf_4 _3933_ (.A(_2526_),
    .X(_2529_));
 sky130_fd_sc_hd__and2_0 _3934_ (.A(_2509_),
    .B(_2529_),
    .X(_0822_));
 sky130_fd_sc_hd__and2_0 _3935_ (.A(_2511_),
    .B(_2529_),
    .X(_0823_));
 sky130_fd_sc_hd__and2_0 _3936_ (.A(_2512_),
    .B(_2529_),
    .X(_0824_));
 sky130_fd_sc_hd__and2_0 _3937_ (.A(_2513_),
    .B(_2529_),
    .X(_0825_));
 sky130_fd_sc_hd__and2_0 _3938_ (.A(_2514_),
    .B(_2529_),
    .X(_0826_));
 sky130_fd_sc_hd__and2_0 _3939_ (.A(_2515_),
    .B(_2529_),
    .X(_0827_));
 sky130_fd_sc_hd__and2_0 _3940_ (.A(_2516_),
    .B(_2529_),
    .X(_0828_));
 sky130_fd_sc_hd__and2_0 _3941_ (.A(_2517_),
    .B(_2529_),
    .X(_0829_));
 sky130_fd_sc_hd__and2_0 _3942_ (.A(_2518_),
    .B(_2529_),
    .X(_0830_));
 sky130_fd_sc_hd__and2_0 _3943_ (.A(_2519_),
    .B(_2529_),
    .X(_0831_));
 sky130_fd_sc_hd__and2_0 _3944_ (.A(_2520_),
    .B(_2526_),
    .X(_0832_));
 sky130_fd_sc_hd__and2_0 _3945_ (.A(_2521_),
    .B(_2526_),
    .X(_0833_));
 sky130_fd_sc_hd__nor2_2 _3946_ (.A(_1132_),
    .B(_1144_),
    .Y(_2530_));
 sky130_fd_sc_hd__clkbuf_4 _3947_ (.A(_2530_),
    .X(_2531_));
 sky130_fd_sc_hd__and2_0 _3948_ (.A(_2486_),
    .B(_2531_),
    .X(_0834_));
 sky130_fd_sc_hd__and2_0 _3949_ (.A(_2489_),
    .B(_2531_),
    .X(_0835_));
 sky130_fd_sc_hd__and2_0 _3950_ (.A(_2490_),
    .B(_2531_),
    .X(_0836_));
 sky130_fd_sc_hd__and2_0 _3951_ (.A(_2491_),
    .B(_2531_),
    .X(_0837_));
 sky130_fd_sc_hd__and2_0 _3952_ (.A(_2492_),
    .B(_2531_),
    .X(_0838_));
 sky130_fd_sc_hd__and2_0 _3953_ (.A(_2493_),
    .B(_2531_),
    .X(_0839_));
 sky130_fd_sc_hd__and2_0 _3954_ (.A(_2494_),
    .B(_2531_),
    .X(_0840_));
 sky130_fd_sc_hd__and2_0 _3955_ (.A(_2495_),
    .B(_2531_),
    .X(_0841_));
 sky130_fd_sc_hd__and2_0 _3956_ (.A(_2496_),
    .B(_2531_),
    .X(_0842_));
 sky130_fd_sc_hd__and2_0 _3957_ (.A(_2497_),
    .B(_2531_),
    .X(_0843_));
 sky130_fd_sc_hd__buf_4 _3958_ (.A(_2530_),
    .X(_2532_));
 sky130_fd_sc_hd__and2_0 _3959_ (.A(_2498_),
    .B(_2532_),
    .X(_0844_));
 sky130_fd_sc_hd__and2_0 _3960_ (.A(_2500_),
    .B(_2532_),
    .X(_0845_));
 sky130_fd_sc_hd__and2_0 _3961_ (.A(_2501_),
    .B(_2532_),
    .X(_0846_));
 sky130_fd_sc_hd__and2_0 _3962_ (.A(_2502_),
    .B(_2532_),
    .X(_0847_));
 sky130_fd_sc_hd__and2_0 _3963_ (.A(_2503_),
    .B(_2532_),
    .X(_0848_));
 sky130_fd_sc_hd__and2_0 _3964_ (.A(_2504_),
    .B(_2532_),
    .X(_0849_));
 sky130_fd_sc_hd__and2_0 _3965_ (.A(_2505_),
    .B(_2532_),
    .X(_0850_));
 sky130_fd_sc_hd__and2_0 _3966_ (.A(_2506_),
    .B(_2532_),
    .X(_0851_));
 sky130_fd_sc_hd__and2_0 _3967_ (.A(_2507_),
    .B(_2532_),
    .X(_0852_));
 sky130_fd_sc_hd__and2_0 _3968_ (.A(_2508_),
    .B(_2532_),
    .X(_0853_));
 sky130_fd_sc_hd__clkbuf_4 _3969_ (.A(_2530_),
    .X(_2533_));
 sky130_fd_sc_hd__and2_0 _3970_ (.A(_2509_),
    .B(_2533_),
    .X(_0854_));
 sky130_fd_sc_hd__and2_0 _3971_ (.A(_2511_),
    .B(_2533_),
    .X(_0855_));
 sky130_fd_sc_hd__and2_0 _3972_ (.A(_2512_),
    .B(_2533_),
    .X(_0856_));
 sky130_fd_sc_hd__and2_0 _3973_ (.A(_2513_),
    .B(_2533_),
    .X(_0857_));
 sky130_fd_sc_hd__and2_0 _3974_ (.A(_2514_),
    .B(_2533_),
    .X(_0858_));
 sky130_fd_sc_hd__and2_0 _3975_ (.A(_2515_),
    .B(_2533_),
    .X(_0859_));
 sky130_fd_sc_hd__and2_0 _3976_ (.A(_2516_),
    .B(_2533_),
    .X(_0860_));
 sky130_fd_sc_hd__and2_0 _3977_ (.A(_2517_),
    .B(_2533_),
    .X(_0861_));
 sky130_fd_sc_hd__and2_0 _3978_ (.A(_2518_),
    .B(_2533_),
    .X(_0862_));
 sky130_fd_sc_hd__and2_0 _3979_ (.A(_2519_),
    .B(_2533_),
    .X(_0863_));
 sky130_fd_sc_hd__and2_0 _3980_ (.A(_2520_),
    .B(_2530_),
    .X(_0864_));
 sky130_fd_sc_hd__and2_0 _3981_ (.A(_2521_),
    .B(_2530_),
    .X(_0865_));
 sky130_fd_sc_hd__nor2_2 _3982_ (.A(_1134_),
    .B(_1144_),
    .Y(_2534_));
 sky130_fd_sc_hd__buf_4 _3983_ (.A(_2534_),
    .X(_2535_));
 sky130_fd_sc_hd__and2_0 _3984_ (.A(_2486_),
    .B(_2535_),
    .X(_0866_));
 sky130_fd_sc_hd__and2_0 _3985_ (.A(_2489_),
    .B(_2535_),
    .X(_0867_));
 sky130_fd_sc_hd__and2_0 _3986_ (.A(_2490_),
    .B(_2535_),
    .X(_0868_));
 sky130_fd_sc_hd__and2_0 _3987_ (.A(_2491_),
    .B(_2535_),
    .X(_0869_));
 sky130_fd_sc_hd__and2_0 _3988_ (.A(_2492_),
    .B(_2535_),
    .X(_0870_));
 sky130_fd_sc_hd__and2_0 _3989_ (.A(_2493_),
    .B(_2535_),
    .X(_0871_));
 sky130_fd_sc_hd__and2_0 _3990_ (.A(_2494_),
    .B(_2535_),
    .X(_0872_));
 sky130_fd_sc_hd__and2_0 _3991_ (.A(_2495_),
    .B(_2535_),
    .X(_0873_));
 sky130_fd_sc_hd__and2_0 _3992_ (.A(_2496_),
    .B(_2535_),
    .X(_0874_));
 sky130_fd_sc_hd__and2_0 _3993_ (.A(_2497_),
    .B(_2535_),
    .X(_0875_));
 sky130_fd_sc_hd__buf_4 _3994_ (.A(_2534_),
    .X(_2536_));
 sky130_fd_sc_hd__and2_0 _3995_ (.A(_2498_),
    .B(_2536_),
    .X(_0876_));
 sky130_fd_sc_hd__and2_0 _3996_ (.A(_2500_),
    .B(_2536_),
    .X(_0877_));
 sky130_fd_sc_hd__and2_0 _3997_ (.A(_2501_),
    .B(_2536_),
    .X(_0878_));
 sky130_fd_sc_hd__and2_0 _3998_ (.A(_2502_),
    .B(_2536_),
    .X(_0879_));
 sky130_fd_sc_hd__and2_0 _3999_ (.A(_2503_),
    .B(_2536_),
    .X(_0880_));
 sky130_fd_sc_hd__and2_0 _4000_ (.A(_2504_),
    .B(_2536_),
    .X(_0881_));
 sky130_fd_sc_hd__and2_0 _4001_ (.A(_2505_),
    .B(_2536_),
    .X(_0882_));
 sky130_fd_sc_hd__and2_0 _4002_ (.A(_2506_),
    .B(_2536_),
    .X(_0883_));
 sky130_fd_sc_hd__and2_0 _4003_ (.A(_2507_),
    .B(_2536_),
    .X(_0884_));
 sky130_fd_sc_hd__and2_0 _4004_ (.A(_2508_),
    .B(_2536_),
    .X(_0885_));
 sky130_fd_sc_hd__buf_4 _4005_ (.A(_2534_),
    .X(_2537_));
 sky130_fd_sc_hd__and2_0 _4006_ (.A(_2509_),
    .B(_2537_),
    .X(_0886_));
 sky130_fd_sc_hd__and2_0 _4007_ (.A(_2511_),
    .B(_2537_),
    .X(_0887_));
 sky130_fd_sc_hd__and2_0 _4008_ (.A(_2512_),
    .B(_2537_),
    .X(_0888_));
 sky130_fd_sc_hd__and2_0 _4009_ (.A(_2513_),
    .B(_2537_),
    .X(_0889_));
 sky130_fd_sc_hd__and2_0 _4010_ (.A(_2514_),
    .B(_2537_),
    .X(_0890_));
 sky130_fd_sc_hd__and2_0 _4011_ (.A(_2515_),
    .B(_2537_),
    .X(_0891_));
 sky130_fd_sc_hd__and2_0 _4012_ (.A(_2516_),
    .B(_2537_),
    .X(_0892_));
 sky130_fd_sc_hd__and2_0 _4013_ (.A(_2517_),
    .B(_2537_),
    .X(_0893_));
 sky130_fd_sc_hd__and2_0 _4014_ (.A(_2518_),
    .B(_2537_),
    .X(_0894_));
 sky130_fd_sc_hd__and2_0 _4015_ (.A(_2519_),
    .B(_2537_),
    .X(_0895_));
 sky130_fd_sc_hd__and2_0 _4016_ (.A(_2520_),
    .B(_2534_),
    .X(_0896_));
 sky130_fd_sc_hd__and2_0 _4017_ (.A(_2521_),
    .B(_2534_),
    .X(_0897_));
 sky130_fd_sc_hd__nor2_4 _4018_ (.A(_1124_),
    .B(_1135_),
    .Y(_2538_));
 sky130_fd_sc_hd__buf_4 _4019_ (.A(_2538_),
    .X(_2539_));
 sky130_fd_sc_hd__and2_0 _4020_ (.A(_2486_),
    .B(_2539_),
    .X(_0898_));
 sky130_fd_sc_hd__and2_0 _4021_ (.A(_2489_),
    .B(_2539_),
    .X(_0899_));
 sky130_fd_sc_hd__and2_0 _4022_ (.A(_2490_),
    .B(_2539_),
    .X(_0900_));
 sky130_fd_sc_hd__and2_0 _4023_ (.A(_2491_),
    .B(_2539_),
    .X(_0901_));
 sky130_fd_sc_hd__and2_0 _4024_ (.A(_2492_),
    .B(_2539_),
    .X(_0902_));
 sky130_fd_sc_hd__and2_0 _4025_ (.A(_2493_),
    .B(_2539_),
    .X(_0903_));
 sky130_fd_sc_hd__and2_0 _4026_ (.A(_2494_),
    .B(_2539_),
    .X(_0904_));
 sky130_fd_sc_hd__and2_0 _4027_ (.A(_2495_),
    .B(_2539_),
    .X(_0905_));
 sky130_fd_sc_hd__and2_0 _4028_ (.A(_2496_),
    .B(_2539_),
    .X(_0906_));
 sky130_fd_sc_hd__and2_0 _4029_ (.A(_2497_),
    .B(_2539_),
    .X(_0907_));
 sky130_fd_sc_hd__buf_4 _4030_ (.A(_2538_),
    .X(_2540_));
 sky130_fd_sc_hd__and2_0 _4031_ (.A(_2498_),
    .B(_2540_),
    .X(_0908_));
 sky130_fd_sc_hd__and2_0 _4032_ (.A(_2500_),
    .B(_2540_),
    .X(_0909_));
 sky130_fd_sc_hd__and2_0 _4033_ (.A(_2501_),
    .B(_2540_),
    .X(_0910_));
 sky130_fd_sc_hd__and2_0 _4034_ (.A(_2502_),
    .B(_2540_),
    .X(_0911_));
 sky130_fd_sc_hd__and2_0 _4035_ (.A(_2503_),
    .B(_2540_),
    .X(_0912_));
 sky130_fd_sc_hd__and2_0 _4036_ (.A(_2504_),
    .B(_2540_),
    .X(_0913_));
 sky130_fd_sc_hd__and2_0 _4037_ (.A(_2505_),
    .B(_2540_),
    .X(_0914_));
 sky130_fd_sc_hd__and2_0 _4038_ (.A(_2506_),
    .B(_2540_),
    .X(_0915_));
 sky130_fd_sc_hd__and2_0 _4039_ (.A(_2507_),
    .B(_2540_),
    .X(_0916_));
 sky130_fd_sc_hd__and2_0 _4040_ (.A(_2508_),
    .B(_2540_),
    .X(_0917_));
 sky130_fd_sc_hd__buf_4 _4041_ (.A(_2538_),
    .X(_2541_));
 sky130_fd_sc_hd__and2_0 _4042_ (.A(_2509_),
    .B(_2541_),
    .X(_0918_));
 sky130_fd_sc_hd__and2_0 _4043_ (.A(_2511_),
    .B(_2541_),
    .X(_0919_));
 sky130_fd_sc_hd__and2_0 _4044_ (.A(_2512_),
    .B(_2541_),
    .X(_0920_));
 sky130_fd_sc_hd__and2_0 _4045_ (.A(_2513_),
    .B(_2541_),
    .X(_0921_));
 sky130_fd_sc_hd__and2_0 _4046_ (.A(_2514_),
    .B(_2541_),
    .X(_0922_));
 sky130_fd_sc_hd__and2_0 _4047_ (.A(_2515_),
    .B(_2541_),
    .X(_0923_));
 sky130_fd_sc_hd__and2_0 _4048_ (.A(_2516_),
    .B(_2541_),
    .X(_0924_));
 sky130_fd_sc_hd__and2_0 _4049_ (.A(_2517_),
    .B(_2541_),
    .X(_0925_));
 sky130_fd_sc_hd__and2_0 _4050_ (.A(_2518_),
    .B(_2541_),
    .X(_0926_));
 sky130_fd_sc_hd__and2_0 _4051_ (.A(_2519_),
    .B(_2541_),
    .X(_0927_));
 sky130_fd_sc_hd__and2_0 _4052_ (.A(_2520_),
    .B(_2538_),
    .X(_0928_));
 sky130_fd_sc_hd__and2_0 _4053_ (.A(_2521_),
    .B(_2538_),
    .X(_0929_));
 sky130_fd_sc_hd__nor2_2 _4054_ (.A(_1127_),
    .B(_1147_),
    .Y(_2542_));
 sky130_fd_sc_hd__buf_4 _4055_ (.A(_2542_),
    .X(_2543_));
 sky130_fd_sc_hd__and2_0 _4056_ (.A(_2486_),
    .B(_2543_),
    .X(_0930_));
 sky130_fd_sc_hd__and2_0 _4057_ (.A(_2489_),
    .B(_2543_),
    .X(_0931_));
 sky130_fd_sc_hd__and2_0 _4058_ (.A(_2490_),
    .B(_2543_),
    .X(_0932_));
 sky130_fd_sc_hd__and2_0 _4059_ (.A(_2491_),
    .B(_2543_),
    .X(_0933_));
 sky130_fd_sc_hd__and2_0 _4060_ (.A(_2492_),
    .B(_2543_),
    .X(_0934_));
 sky130_fd_sc_hd__and2_0 _4061_ (.A(_2493_),
    .B(_2543_),
    .X(_0935_));
 sky130_fd_sc_hd__and2_0 _4062_ (.A(_2494_),
    .B(_2543_),
    .X(_0936_));
 sky130_fd_sc_hd__and2_0 _4063_ (.A(_2495_),
    .B(_2543_),
    .X(_0937_));
 sky130_fd_sc_hd__and2_0 _4064_ (.A(_2496_),
    .B(_2543_),
    .X(_0938_));
 sky130_fd_sc_hd__and2_0 _4065_ (.A(_2497_),
    .B(_2543_),
    .X(_0939_));
 sky130_fd_sc_hd__buf_4 _4066_ (.A(_2542_),
    .X(_2544_));
 sky130_fd_sc_hd__and2_0 _4067_ (.A(_2498_),
    .B(_2544_),
    .X(_0940_));
 sky130_fd_sc_hd__and2_0 _4068_ (.A(_2500_),
    .B(_2544_),
    .X(_0941_));
 sky130_fd_sc_hd__and2_0 _4069_ (.A(_2501_),
    .B(_2544_),
    .X(_0942_));
 sky130_fd_sc_hd__and2_0 _4070_ (.A(_2502_),
    .B(_2544_),
    .X(_0943_));
 sky130_fd_sc_hd__and2_0 _4071_ (.A(_2503_),
    .B(_2544_),
    .X(_0944_));
 sky130_fd_sc_hd__and2_0 _4072_ (.A(_2504_),
    .B(_2544_),
    .X(_0945_));
 sky130_fd_sc_hd__and2_0 _4073_ (.A(_2505_),
    .B(_2544_),
    .X(_0946_));
 sky130_fd_sc_hd__and2_0 _4074_ (.A(_2506_),
    .B(_2544_),
    .X(_0947_));
 sky130_fd_sc_hd__and2_0 _4075_ (.A(_2507_),
    .B(_2544_),
    .X(_0948_));
 sky130_fd_sc_hd__and2_0 _4076_ (.A(_2508_),
    .B(_2544_),
    .X(_0949_));
 sky130_fd_sc_hd__buf_4 _4077_ (.A(_2542_),
    .X(_2545_));
 sky130_fd_sc_hd__and2_0 _4078_ (.A(_2509_),
    .B(_2545_),
    .X(_0950_));
 sky130_fd_sc_hd__and2_0 _4079_ (.A(_2511_),
    .B(_2545_),
    .X(_0951_));
 sky130_fd_sc_hd__and2_0 _4080_ (.A(_2512_),
    .B(_2545_),
    .X(_0952_));
 sky130_fd_sc_hd__and2_0 _4081_ (.A(_2513_),
    .B(_2545_),
    .X(_0953_));
 sky130_fd_sc_hd__and2_0 _4082_ (.A(_2514_),
    .B(_2545_),
    .X(_0954_));
 sky130_fd_sc_hd__and2_0 _4083_ (.A(_2515_),
    .B(_2545_),
    .X(_0955_));
 sky130_fd_sc_hd__and2_0 _4084_ (.A(_2516_),
    .B(_2545_),
    .X(_0956_));
 sky130_fd_sc_hd__and2_0 _4085_ (.A(_2517_),
    .B(_2545_),
    .X(_0957_));
 sky130_fd_sc_hd__and2_0 _4086_ (.A(_2518_),
    .B(_2545_),
    .X(_0958_));
 sky130_fd_sc_hd__and2_0 _4087_ (.A(_2519_),
    .B(_2545_),
    .X(_0959_));
 sky130_fd_sc_hd__and2_0 _4088_ (.A(_2520_),
    .B(_2542_),
    .X(_0960_));
 sky130_fd_sc_hd__and2_0 _4089_ (.A(_2521_),
    .B(_2542_),
    .X(_0961_));
 sky130_fd_sc_hd__nor2_2 _4090_ (.A(_1137_),
    .B(_1147_),
    .Y(_2546_));
 sky130_fd_sc_hd__buf_4 _4091_ (.A(_2546_),
    .X(_2547_));
 sky130_fd_sc_hd__and2_0 _4092_ (.A(_2486_),
    .B(_2547_),
    .X(_0962_));
 sky130_fd_sc_hd__and2_0 _4093_ (.A(_2489_),
    .B(_2547_),
    .X(_0963_));
 sky130_fd_sc_hd__and2_0 _4094_ (.A(_2490_),
    .B(_2547_),
    .X(_0964_));
 sky130_fd_sc_hd__and2_0 _4095_ (.A(_2491_),
    .B(_2547_),
    .X(_0965_));
 sky130_fd_sc_hd__and2_0 _4096_ (.A(_2492_),
    .B(_2547_),
    .X(_0966_));
 sky130_fd_sc_hd__and2_0 _4097_ (.A(_2493_),
    .B(_2547_),
    .X(_0967_));
 sky130_fd_sc_hd__and2_0 _4098_ (.A(_2494_),
    .B(_2547_),
    .X(_0968_));
 sky130_fd_sc_hd__and2_0 _4099_ (.A(_2495_),
    .B(_2547_),
    .X(_0969_));
 sky130_fd_sc_hd__and2_0 _4100_ (.A(_2496_),
    .B(_2547_),
    .X(_0970_));
 sky130_fd_sc_hd__and2_0 _4101_ (.A(_2497_),
    .B(_2547_),
    .X(_0971_));
 sky130_fd_sc_hd__buf_4 _4102_ (.A(_2546_),
    .X(_2548_));
 sky130_fd_sc_hd__and2_0 _4103_ (.A(_2498_),
    .B(_2548_),
    .X(_0972_));
 sky130_fd_sc_hd__and2_0 _4104_ (.A(_2500_),
    .B(_2548_),
    .X(_0973_));
 sky130_fd_sc_hd__and2_0 _4105_ (.A(_2501_),
    .B(_2548_),
    .X(_0974_));
 sky130_fd_sc_hd__and2_0 _4106_ (.A(_2502_),
    .B(_2548_),
    .X(_0975_));
 sky130_fd_sc_hd__and2_0 _4107_ (.A(_2503_),
    .B(_2548_),
    .X(_0976_));
 sky130_fd_sc_hd__and2_0 _4108_ (.A(_2504_),
    .B(_2548_),
    .X(_0977_));
 sky130_fd_sc_hd__and2_0 _4109_ (.A(_2505_),
    .B(_2548_),
    .X(_0978_));
 sky130_fd_sc_hd__and2_0 _4110_ (.A(_2506_),
    .B(_2548_),
    .X(_0979_));
 sky130_fd_sc_hd__and2_0 _4111_ (.A(_2507_),
    .B(_2548_),
    .X(_0980_));
 sky130_fd_sc_hd__and2_0 _4112_ (.A(_2508_),
    .B(_2548_),
    .X(_0981_));
 sky130_fd_sc_hd__buf_4 _4113_ (.A(_2546_),
    .X(_2549_));
 sky130_fd_sc_hd__and2_0 _4114_ (.A(_2509_),
    .B(_2549_),
    .X(_0982_));
 sky130_fd_sc_hd__and2_0 _4115_ (.A(_2511_),
    .B(_2549_),
    .X(_0983_));
 sky130_fd_sc_hd__and2_0 _4116_ (.A(_2512_),
    .B(_2549_),
    .X(_0984_));
 sky130_fd_sc_hd__and2_0 _4117_ (.A(_2513_),
    .B(_2549_),
    .X(_0985_));
 sky130_fd_sc_hd__and2_0 _4118_ (.A(_2514_),
    .B(_2549_),
    .X(_0986_));
 sky130_fd_sc_hd__and2_0 _4119_ (.A(_2515_),
    .B(_2549_),
    .X(_0987_));
 sky130_fd_sc_hd__and2_0 _4120_ (.A(_2516_),
    .B(_2549_),
    .X(_0988_));
 sky130_fd_sc_hd__and2_0 _4121_ (.A(_2517_),
    .B(_2549_),
    .X(_0989_));
 sky130_fd_sc_hd__and2_0 _4122_ (.A(_2518_),
    .B(_2549_),
    .X(_0990_));
 sky130_fd_sc_hd__and2_0 _4123_ (.A(_2519_),
    .B(_2549_),
    .X(_0991_));
 sky130_fd_sc_hd__and2_0 _4124_ (.A(_2520_),
    .B(_2546_),
    .X(_0992_));
 sky130_fd_sc_hd__and2_0 _4125_ (.A(_2521_),
    .B(_2546_),
    .X(_0993_));
 sky130_fd_sc_hd__nor2_2 _4126_ (.A(_1132_),
    .B(_1147_),
    .Y(_2550_));
 sky130_fd_sc_hd__buf_4 _4127_ (.A(_2550_),
    .X(_2551_));
 sky130_fd_sc_hd__and2_0 _4128_ (.A(_2486_),
    .B(_2551_),
    .X(_0994_));
 sky130_fd_sc_hd__and2_0 _4129_ (.A(_2489_),
    .B(_2551_),
    .X(_0995_));
 sky130_fd_sc_hd__and2_0 _4130_ (.A(_2490_),
    .B(_2551_),
    .X(_0996_));
 sky130_fd_sc_hd__and2_0 _4131_ (.A(_2491_),
    .B(_2551_),
    .X(_0997_));
 sky130_fd_sc_hd__and2_0 _4132_ (.A(_2492_),
    .B(_2551_),
    .X(_0998_));
 sky130_fd_sc_hd__and2_0 _4133_ (.A(_2493_),
    .B(_2551_),
    .X(_0999_));
 sky130_fd_sc_hd__and2_0 _4134_ (.A(_2494_),
    .B(_2551_),
    .X(_1000_));
 sky130_fd_sc_hd__and2_0 _4135_ (.A(_2495_),
    .B(_2551_),
    .X(_1001_));
 sky130_fd_sc_hd__and2_0 _4136_ (.A(_2496_),
    .B(_2551_),
    .X(_1002_));
 sky130_fd_sc_hd__and2_0 _4137_ (.A(_2497_),
    .B(_2551_),
    .X(_1003_));
 sky130_fd_sc_hd__buf_4 _4138_ (.A(_2550_),
    .X(_2552_));
 sky130_fd_sc_hd__and2_0 _4139_ (.A(_2498_),
    .B(_2552_),
    .X(_1004_));
 sky130_fd_sc_hd__and2_0 _4140_ (.A(_2500_),
    .B(_2552_),
    .X(_1005_));
 sky130_fd_sc_hd__and2_0 _4141_ (.A(_2501_),
    .B(_2552_),
    .X(_1006_));
 sky130_fd_sc_hd__and2_0 _4142_ (.A(_2502_),
    .B(_2552_),
    .X(_1007_));
 sky130_fd_sc_hd__and2_0 _4143_ (.A(_2503_),
    .B(_2552_),
    .X(_1008_));
 sky130_fd_sc_hd__and2_0 _4144_ (.A(_2504_),
    .B(_2552_),
    .X(_1009_));
 sky130_fd_sc_hd__and2_0 _4145_ (.A(_2505_),
    .B(_2552_),
    .X(_1010_));
 sky130_fd_sc_hd__and2_0 _4146_ (.A(_2506_),
    .B(_2552_),
    .X(_1011_));
 sky130_fd_sc_hd__and2_0 _4147_ (.A(_2507_),
    .B(_2552_),
    .X(_1012_));
 sky130_fd_sc_hd__and2_0 _4148_ (.A(_2508_),
    .B(_2552_),
    .X(_1013_));
 sky130_fd_sc_hd__buf_4 _4149_ (.A(_2550_),
    .X(_2553_));
 sky130_fd_sc_hd__and2_0 _4150_ (.A(_2509_),
    .B(_2553_),
    .X(_1014_));
 sky130_fd_sc_hd__and2_0 _4151_ (.A(_2511_),
    .B(_2553_),
    .X(_1015_));
 sky130_fd_sc_hd__and2_0 _4152_ (.A(_2512_),
    .B(_2553_),
    .X(_1016_));
 sky130_fd_sc_hd__and2_0 _4153_ (.A(_2513_),
    .B(_2553_),
    .X(_1017_));
 sky130_fd_sc_hd__and2_0 _4154_ (.A(_2514_),
    .B(_2553_),
    .X(_1018_));
 sky130_fd_sc_hd__and2_0 _4155_ (.A(_2515_),
    .B(_2553_),
    .X(_1019_));
 sky130_fd_sc_hd__and2_0 _4156_ (.A(_2516_),
    .B(_2553_),
    .X(_1020_));
 sky130_fd_sc_hd__and2_0 _4157_ (.A(_2517_),
    .B(_2553_),
    .X(_1021_));
 sky130_fd_sc_hd__and2_0 _4158_ (.A(_2518_),
    .B(_2553_),
    .X(_1022_));
 sky130_fd_sc_hd__and2_0 _4159_ (.A(_2519_),
    .B(_2553_),
    .X(_1023_));
 sky130_fd_sc_hd__and2_0 _4160_ (.A(_2520_),
    .B(_2550_),
    .X(_1024_));
 sky130_fd_sc_hd__and2_0 _4161_ (.A(_2521_),
    .B(_2550_),
    .X(_1025_));
 sky130_fd_sc_hd__nor2_2 _4162_ (.A(_1134_),
    .B(_1147_),
    .Y(_2554_));
 sky130_fd_sc_hd__buf_4 _4163_ (.A(_2554_),
    .X(_2555_));
 sky130_fd_sc_hd__and2_0 _4164_ (.A(_2486_),
    .B(_2555_),
    .X(_1026_));
 sky130_fd_sc_hd__and2_0 _4165_ (.A(_2489_),
    .B(_2555_),
    .X(_1027_));
 sky130_fd_sc_hd__and2_0 _4166_ (.A(_2490_),
    .B(_2555_),
    .X(_1028_));
 sky130_fd_sc_hd__and2_0 _4167_ (.A(_2491_),
    .B(_2555_),
    .X(_1029_));
 sky130_fd_sc_hd__and2_0 _4168_ (.A(_2492_),
    .B(_2555_),
    .X(_1030_));
 sky130_fd_sc_hd__and2_0 _4169_ (.A(_2493_),
    .B(_2555_),
    .X(_1031_));
 sky130_fd_sc_hd__and2_0 _4170_ (.A(_2494_),
    .B(_2555_),
    .X(_1032_));
 sky130_fd_sc_hd__and2_0 _4171_ (.A(_2495_),
    .B(_2555_),
    .X(_1033_));
 sky130_fd_sc_hd__and2_0 _4172_ (.A(_2496_),
    .B(_2555_),
    .X(_1034_));
 sky130_fd_sc_hd__and2_0 _4173_ (.A(_2497_),
    .B(_2555_),
    .X(_1035_));
 sky130_fd_sc_hd__buf_4 _4174_ (.A(_2554_),
    .X(_2556_));
 sky130_fd_sc_hd__and2_0 _4175_ (.A(_2498_),
    .B(_2556_),
    .X(_1036_));
 sky130_fd_sc_hd__and2_0 _4176_ (.A(_2500_),
    .B(_2556_),
    .X(_1037_));
 sky130_fd_sc_hd__and2_0 _4177_ (.A(_2501_),
    .B(_2556_),
    .X(_1038_));
 sky130_fd_sc_hd__and2_0 _4178_ (.A(_2502_),
    .B(_2556_),
    .X(_1039_));
 sky130_fd_sc_hd__and2_0 _4179_ (.A(_2503_),
    .B(_2556_),
    .X(_1040_));
 sky130_fd_sc_hd__and2_0 _4180_ (.A(_2504_),
    .B(_2556_),
    .X(_1041_));
 sky130_fd_sc_hd__and2_0 _4181_ (.A(_2505_),
    .B(_2556_),
    .X(_1042_));
 sky130_fd_sc_hd__and2_0 _4182_ (.A(_2506_),
    .B(_2556_),
    .X(_1043_));
 sky130_fd_sc_hd__and2_0 _4183_ (.A(_2507_),
    .B(_2556_),
    .X(_1044_));
 sky130_fd_sc_hd__and2_0 _4184_ (.A(_2508_),
    .B(_2556_),
    .X(_1045_));
 sky130_fd_sc_hd__buf_4 _4185_ (.A(_2554_),
    .X(_2557_));
 sky130_fd_sc_hd__and2_0 _4186_ (.A(_2509_),
    .B(_2557_),
    .X(_1046_));
 sky130_fd_sc_hd__and2_0 _4187_ (.A(_2511_),
    .B(_2557_),
    .X(_1047_));
 sky130_fd_sc_hd__and2_0 _4188_ (.A(_2512_),
    .B(_2557_),
    .X(_1048_));
 sky130_fd_sc_hd__and2_0 _4189_ (.A(_2513_),
    .B(_2557_),
    .X(_1049_));
 sky130_fd_sc_hd__and2_0 _4190_ (.A(_2514_),
    .B(_2557_),
    .X(_1050_));
 sky130_fd_sc_hd__and2_0 _4191_ (.A(_2515_),
    .B(_2557_),
    .X(_1051_));
 sky130_fd_sc_hd__and2_0 _4192_ (.A(_2516_),
    .B(_2557_),
    .X(_1052_));
 sky130_fd_sc_hd__and2_0 _4193_ (.A(_2517_),
    .B(_2557_),
    .X(_1053_));
 sky130_fd_sc_hd__and2_0 _4194_ (.A(_2518_),
    .B(_2557_),
    .X(_1054_));
 sky130_fd_sc_hd__and2_0 _4195_ (.A(_2519_),
    .B(_2557_),
    .X(_1055_));
 sky130_fd_sc_hd__and2_0 _4196_ (.A(_2520_),
    .B(_2554_),
    .X(_1056_));
 sky130_fd_sc_hd__and2_0 _4197_ (.A(_2521_),
    .B(_2554_),
    .X(_1057_));
 sky130_fd_sc_hd__nor2_8 _4198_ (.A(_1127_),
    .B(_1131_),
    .Y(_2558_));
 sky130_fd_sc_hd__buf_4 _4199_ (.A(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__and2_0 _4200_ (.A(net11),
    .B(_2559_),
    .X(_1058_));
 sky130_fd_sc_hd__and2_0 _4201_ (.A(net12),
    .B(_2559_),
    .X(_1059_));
 sky130_fd_sc_hd__and2_0 _4202_ (.A(net13),
    .B(_2559_),
    .X(_1060_));
 sky130_fd_sc_hd__and2_0 _4203_ (.A(net14),
    .B(_2559_),
    .X(_1061_));
 sky130_fd_sc_hd__and2_0 _4204_ (.A(net15),
    .B(_2559_),
    .X(_1062_));
 sky130_fd_sc_hd__and2_0 _4205_ (.A(net16),
    .B(_2559_),
    .X(_1063_));
 sky130_fd_sc_hd__and2_0 _4206_ (.A(net17),
    .B(_2559_),
    .X(_1064_));
 sky130_fd_sc_hd__and2_0 _4207_ (.A(net18),
    .B(_2559_),
    .X(_1065_));
 sky130_fd_sc_hd__and2_0 _4208_ (.A(net19),
    .B(_2559_),
    .X(_1066_));
 sky130_fd_sc_hd__and2_0 _4209_ (.A(net20),
    .B(_2559_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_4 _4210_ (.A(_2558_),
    .X(_2560_));
 sky130_fd_sc_hd__and2_0 _4211_ (.A(net21),
    .B(_2560_),
    .X(_1068_));
 sky130_fd_sc_hd__and2_0 _4212_ (.A(net22),
    .B(_2560_),
    .X(_1069_));
 sky130_fd_sc_hd__and2_0 _4213_ (.A(net23),
    .B(_2560_),
    .X(_1070_));
 sky130_fd_sc_hd__and2_0 _4214_ (.A(net24),
    .B(_2560_),
    .X(_1071_));
 sky130_fd_sc_hd__and2_0 _4215_ (.A(net25),
    .B(_2560_),
    .X(_1072_));
 sky130_fd_sc_hd__and2_0 _4216_ (.A(net26),
    .B(_2560_),
    .X(_1073_));
 sky130_fd_sc_hd__and2_0 _4217_ (.A(net27),
    .B(_2560_),
    .X(_1074_));
 sky130_fd_sc_hd__and2_0 _4218_ (.A(net28),
    .B(_2560_),
    .X(_1075_));
 sky130_fd_sc_hd__and2_0 _4219_ (.A(net29),
    .B(_2560_),
    .X(_1076_));
 sky130_fd_sc_hd__and2_0 _4220_ (.A(net30),
    .B(_2560_),
    .X(_1077_));
 sky130_fd_sc_hd__buf_4 _4221_ (.A(_2558_),
    .X(_2561_));
 sky130_fd_sc_hd__and2_0 _4222_ (.A(net31),
    .B(_2561_),
    .X(_1078_));
 sky130_fd_sc_hd__and2_0 _4223_ (.A(net32),
    .B(_2561_),
    .X(_1079_));
 sky130_fd_sc_hd__and2_0 _4224_ (.A(net33),
    .B(_2561_),
    .X(_1080_));
 sky130_fd_sc_hd__and2_0 _4225_ (.A(net34),
    .B(_2561_),
    .X(_1081_));
 sky130_fd_sc_hd__and2_0 _4226_ (.A(net35),
    .B(_2561_),
    .X(_1082_));
 sky130_fd_sc_hd__and2_0 _4227_ (.A(net36),
    .B(_2561_),
    .X(_1083_));
 sky130_fd_sc_hd__and2_0 _4228_ (.A(net37),
    .B(_2561_),
    .X(_1084_));
 sky130_fd_sc_hd__and2_0 _4229_ (.A(net38),
    .B(_2561_),
    .X(_1085_));
 sky130_fd_sc_hd__and2_0 _4230_ (.A(net39),
    .B(_2561_),
    .X(_1086_));
 sky130_fd_sc_hd__and2_0 _4231_ (.A(net40),
    .B(_2561_),
    .X(_1087_));
 sky130_fd_sc_hd__and2_0 _4232_ (.A(net41),
    .B(_2558_),
    .X(_1088_));
 sky130_fd_sc_hd__and2_0 _4233_ (.A(net42),
    .B(_2558_),
    .X(_1089_));
 sky130_fd_sc_hd__nor2_8 _4234_ (.A(_1131_),
    .B(_1137_),
    .Y(_2562_));
 sky130_fd_sc_hd__buf_4 _4235_ (.A(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__and2_0 _4236_ (.A(net11),
    .B(_2563_),
    .X(_1090_));
 sky130_fd_sc_hd__and2_0 _4237_ (.A(net12),
    .B(_2563_),
    .X(_1091_));
 sky130_fd_sc_hd__and2_0 _4238_ (.A(net13),
    .B(_2563_),
    .X(_1092_));
 sky130_fd_sc_hd__and2_0 _4239_ (.A(net14),
    .B(_2563_),
    .X(_1093_));
 sky130_fd_sc_hd__and2_0 _4240_ (.A(net15),
    .B(_2563_),
    .X(_1094_));
 sky130_fd_sc_hd__and2_0 _4241_ (.A(net16),
    .B(_2563_),
    .X(_1095_));
 sky130_fd_sc_hd__and2_0 _4242_ (.A(net17),
    .B(_2563_),
    .X(_1096_));
 sky130_fd_sc_hd__and2_0 _4243_ (.A(net18),
    .B(_2563_),
    .X(_1097_));
 sky130_fd_sc_hd__and2_0 _4244_ (.A(net19),
    .B(_2563_),
    .X(_1098_));
 sky130_fd_sc_hd__and2_0 _4245_ (.A(net20),
    .B(_2563_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_4 _4246_ (.A(_2562_),
    .X(_2564_));
 sky130_fd_sc_hd__and2_0 _4247_ (.A(net21),
    .B(_2564_),
    .X(_1100_));
 sky130_fd_sc_hd__and2_0 _4248_ (.A(net22),
    .B(_2564_),
    .X(_1101_));
 sky130_fd_sc_hd__and2_0 _4249_ (.A(net23),
    .B(_2564_),
    .X(_1102_));
 sky130_fd_sc_hd__and2_0 _4250_ (.A(net24),
    .B(_2564_),
    .X(_1103_));
 sky130_fd_sc_hd__and2_0 _4251_ (.A(net25),
    .B(_2564_),
    .X(_1104_));
 sky130_fd_sc_hd__and2_0 _4252_ (.A(net26),
    .B(_2564_),
    .X(_1105_));
 sky130_fd_sc_hd__and2_0 _4253_ (.A(net27),
    .B(_2564_),
    .X(_1106_));
 sky130_fd_sc_hd__and2_0 _4254_ (.A(net28),
    .B(_2564_),
    .X(_1107_));
 sky130_fd_sc_hd__and2_0 _4255_ (.A(net29),
    .B(_2564_),
    .X(_1108_));
 sky130_fd_sc_hd__and2_0 _4256_ (.A(net30),
    .B(_2564_),
    .X(_1109_));
 sky130_fd_sc_hd__buf_4 _4257_ (.A(_2562_),
    .X(_2565_));
 sky130_fd_sc_hd__and2_0 _4258_ (.A(net31),
    .B(_2565_),
    .X(_1110_));
 sky130_fd_sc_hd__and2_0 _4259_ (.A(net32),
    .B(_2565_),
    .X(_1111_));
 sky130_fd_sc_hd__and2_0 _4260_ (.A(net33),
    .B(_2565_),
    .X(_1112_));
 sky130_fd_sc_hd__and2_0 _4261_ (.A(net34),
    .B(_2565_),
    .X(_1113_));
 sky130_fd_sc_hd__and2_0 _4262_ (.A(net35),
    .B(_2565_),
    .X(_1114_));
 sky130_fd_sc_hd__and2_0 _4263_ (.A(net36),
    .B(_2565_),
    .X(_1115_));
 sky130_fd_sc_hd__and2_0 _4264_ (.A(net37),
    .B(_2565_),
    .X(_1116_));
 sky130_fd_sc_hd__and2_0 _4265_ (.A(net38),
    .B(_2565_),
    .X(_1117_));
 sky130_fd_sc_hd__and2_0 _4266_ (.A(net39),
    .B(_2565_),
    .X(_1118_));
 sky130_fd_sc_hd__and2_0 _4267_ (.A(net40),
    .B(_2565_),
    .X(_1119_));
 sky130_fd_sc_hd__and2_0 _4268_ (.A(net41),
    .B(_2562_),
    .X(_1120_));
 sky130_fd_sc_hd__and2_0 _4269_ (.A(net42),
    .B(_2562_),
    .X(_1121_));
 sky130_fd_sc_hd__buf_8 _4270_ (.A(net5),
    .X(_1122_));
 sky130_fd_sc_hd__nand2b_4 _4271_ (.A_N(net3),
    .B(_1122_),
    .Y(_0032_));
 sky130_fd_sc_hd__nand2b_4 _4272_ (.A_N(net4),
    .B(_1122_),
    .Y(_0033_));
 sky130_fd_sc_hd__or3_1 _4273_ (.A(net9),
    .B(net10),
    .C(net8),
    .X(_1123_));
 sky130_fd_sc_hd__buf_6 _4274_ (.A(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__nand2_1 _4275_ (.A(net5),
    .B(net43),
    .Y(_1125_));
 sky130_fd_sc_hd__or3_1 _4276_ (.A(net6),
    .B(net7),
    .C(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__buf_8 _4277_ (.A(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__buf_16 _4278_ (.A(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__buf_8 _4279_ (.A(_1122_),
    .X(_1129_));
 sky130_fd_sc_hd__o21ai_4 _4280_ (.A1(_1124_),
    .A2(_1128_),
    .B1(_1129_),
    .Y(_0031_));
 sky130_fd_sc_hd__nor2_2 _4281_ (.A(net10),
    .B(net8),
    .Y(_1130_));
 sky130_fd_sc_hd__nand2_8 _4282_ (.A(net9),
    .B(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__nand4b_4 _4283_ (.A_N(net6),
    .B(net7),
    .C(net43),
    .D(net5),
    .Y(_1132_));
 sky130_fd_sc_hd__buf_8 _4284_ (.A(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__o21ai_4 _4285_ (.A1(_1131_),
    .A2(_1133_),
    .B1(_1129_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand4_4 _4286_ (.A(_1122_),
    .B(net6),
    .C(net7),
    .D(net43),
    .Y(_1134_));
 sky130_fd_sc_hd__buf_8 _4287_ (.A(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__o21ai_4 _4288_ (.A1(_1131_),
    .A2(_1135_),
    .B1(_1129_),
    .Y(_0029_));
 sky130_fd_sc_hd__nand3b_4 _4289_ (.A_N(net10),
    .B(net8),
    .C(net9),
    .Y(_1136_));
 sky130_fd_sc_hd__o21ai_4 _4290_ (.A1(_1128_),
    .A2(_1136_),
    .B1(_1129_),
    .Y(_0028_));
 sky130_fd_sc_hd__nand4b_4 _4291_ (.A_N(net7),
    .B(net43),
    .C(net5),
    .D(net6),
    .Y(_1137_));
 sky130_fd_sc_hd__clkbuf_16 _4292_ (.A(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__o21ai_4 _4293_ (.A1(_1136_),
    .A2(_1138_),
    .B1(_1129_),
    .Y(_0027_));
 sky130_fd_sc_hd__o21ai_4 _4294_ (.A1(_1133_),
    .A2(_1136_),
    .B1(_1129_),
    .Y(_0026_));
 sky130_fd_sc_hd__o21ai_4 _4295_ (.A1(_1135_),
    .A2(_1136_),
    .B1(_1129_),
    .Y(_0025_));
 sky130_fd_sc_hd__nor2_2 _4296_ (.A(net9),
    .B(net8),
    .Y(_1139_));
 sky130_fd_sc_hd__nand2_8 _4297_ (.A(net10),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__o21ai_4 _4298_ (.A1(_1128_),
    .A2(_1140_),
    .B1(_1129_),
    .Y(_0024_));
 sky130_fd_sc_hd__o21ai_4 _4299_ (.A1(_1138_),
    .A2(_1140_),
    .B1(_1129_),
    .Y(_0023_));
 sky130_fd_sc_hd__o21ai_4 _4300_ (.A1(_1133_),
    .A2(_1140_),
    .B1(_1129_),
    .Y(_0022_));
 sky130_fd_sc_hd__buf_8 _4301_ (.A(_1122_),
    .X(_1141_));
 sky130_fd_sc_hd__o21ai_4 _4302_ (.A1(_1135_),
    .A2(_1140_),
    .B1(_1141_),
    .Y(_0021_));
 sky130_fd_sc_hd__o21ai_4 _4303_ (.A1(_1124_),
    .A2(_1138_),
    .B1(_1141_),
    .Y(_0020_));
 sky130_fd_sc_hd__nand3b_4 _4304_ (.A_N(net9),
    .B(net10),
    .C(net8),
    .Y(_1142_));
 sky130_fd_sc_hd__o21ai_4 _4305_ (.A1(_1128_),
    .A2(_1142_),
    .B1(_1141_),
    .Y(_0019_));
 sky130_fd_sc_hd__o21ai_4 _4306_ (.A1(_1138_),
    .A2(_1142_),
    .B1(_1141_),
    .Y(_0018_));
 sky130_fd_sc_hd__o21ai_4 _4307_ (.A1(_1133_),
    .A2(_1142_),
    .B1(_1141_),
    .Y(_0017_));
 sky130_fd_sc_hd__o21ai_4 _4308_ (.A1(_1135_),
    .A2(_1142_),
    .B1(_1141_),
    .Y(_0016_));
 sky130_fd_sc_hd__nand3b_4 _4309_ (.A_N(net8),
    .B(net10),
    .C(net9),
    .Y(_1143_));
 sky130_fd_sc_hd__o21ai_4 _4310_ (.A1(_1128_),
    .A2(_1143_),
    .B1(_1141_),
    .Y(_0015_));
 sky130_fd_sc_hd__o21ai_4 _4311_ (.A1(_1138_),
    .A2(_1143_),
    .B1(_1141_),
    .Y(_0014_));
 sky130_fd_sc_hd__o21ai_4 _4312_ (.A1(_1133_),
    .A2(_1143_),
    .B1(_1141_),
    .Y(_0013_));
 sky130_fd_sc_hd__o21ai_4 _4313_ (.A1(_1135_),
    .A2(_1143_),
    .B1(_1141_),
    .Y(_0012_));
 sky130_fd_sc_hd__nand3_4 _4314_ (.A(net9),
    .B(net10),
    .C(net8),
    .Y(_1144_));
 sky130_fd_sc_hd__buf_8 _4315_ (.A(_1122_),
    .X(_1145_));
 sky130_fd_sc_hd__o21ai_4 _4316_ (.A1(_1128_),
    .A2(_1144_),
    .B1(_1145_),
    .Y(_0011_));
 sky130_fd_sc_hd__o21ai_4 _4317_ (.A1(_1138_),
    .A2(_1144_),
    .B1(_1145_),
    .Y(_0010_));
 sky130_fd_sc_hd__o21ai_4 _4318_ (.A1(_1124_),
    .A2(_1133_),
    .B1(_1145_),
    .Y(_0009_));
 sky130_fd_sc_hd__o21ai_4 _4319_ (.A1(_1133_),
    .A2(_1144_),
    .B1(_1145_),
    .Y(_0008_));
 sky130_fd_sc_hd__o21ai_4 _4320_ (.A1(_1135_),
    .A2(_1144_),
    .B1(_1145_),
    .Y(_0007_));
 sky130_fd_sc_hd__o21ai_4 _4321_ (.A1(_1124_),
    .A2(_1135_),
    .B1(_1145_),
    .Y(_0006_));
 sky130_fd_sc_hd__or3b_1 _4322_ (.A(net9),
    .B(net10),
    .C_N(net8),
    .X(_1146_));
 sky130_fd_sc_hd__buf_4 _4323_ (.A(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__o21ai_4 _4324_ (.A1(_1128_),
    .A2(_1147_),
    .B1(_1145_),
    .Y(_0005_));
 sky130_fd_sc_hd__o21ai_4 _4325_ (.A1(_1138_),
    .A2(_1147_),
    .B1(_1145_),
    .Y(_0004_));
 sky130_fd_sc_hd__o21ai_4 _4326_ (.A1(_1133_),
    .A2(_1147_),
    .B1(_1145_),
    .Y(_0003_));
 sky130_fd_sc_hd__o21ai_4 _4327_ (.A1(_1135_),
    .A2(_1147_),
    .B1(_1145_),
    .Y(_0002_));
 sky130_fd_sc_hd__o21ai_4 _4328_ (.A1(_1128_),
    .A2(_1131_),
    .B1(_1122_),
    .Y(_0001_));
 sky130_fd_sc_hd__o21ai_4 _4329_ (.A1(_1131_),
    .A2(_1138_),
    .B1(_1122_),
    .Y(_0000_));
 sky130_fd_sc_hd__buf_8 _4330_ (.A(net168),
    .X(_1148_));
 sky130_fd_sc_hd__buf_4 _4331_ (.A(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__buf_6 _4332_ (.A(read_addr1[0]),
    .X(_1150_));
 sky130_fd_sc_hd__clkinvlp_4 _4333_ (.A(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__buf_16 _4334_ (.A(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__buf_12 _4335_ (.A(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__buf_16 _4336_ (.A(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__buf_8 _4337_ (.A(read_addr1[1]),
    .X(_1155_));
 sky130_fd_sc_hd__buf_16 _4338_ (.A(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__buf_8 _4339_ (.A(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__buf_2 _4340_ (.A(read_addr1[2]),
    .X(_1158_));
 sky130_fd_sc_hd__buf_6 _4341_ (.A(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__buf_6 _4342_ (.A(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__mux4_1 _4343_ (.A0(\registers[25][0] ),
    .A1(\registers[27][0] ),
    .A2(\registers[29][0] ),
    .A3(\registers[31][0] ),
    .S0(_1157_),
    .S1(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__buf_6 _4344_ (.A(_1159_),
    .X(_1162_));
 sky130_fd_sc_hd__buf_6 _4345_ (.A(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__mux2i_1 _4346_ (.A0(\registers[24][0] ),
    .A1(\registers[28][0] ),
    .S(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__buf_6 _4347_ (.A(_1150_),
    .X(_1165_));
 sky130_fd_sc_hd__buf_8 _4348_ (.A(_1155_),
    .X(_1166_));
 sky130_fd_sc_hd__buf_8 _4349_ (.A(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__nor2_2 _4350_ (.A(_1165_),
    .B(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__buf_6 _4351_ (.A(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__nand2_1 _4352_ (.A(_1164_),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__mux2i_1 _4353_ (.A0(\registers[26][0] ),
    .A1(\registers[30][0] ),
    .S(_1163_),
    .Y(_1171_));
 sky130_fd_sc_hd__nor2b_2 _4354_ (.A(_1165_),
    .B_N(_1167_),
    .Y(_1172_));
 sky130_fd_sc_hd__buf_6 _4355_ (.A(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__nand2_1 _4356_ (.A(_1171_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__buf_8 _4357_ (.A(net1),
    .X(_1175_));
 sky130_fd_sc_hd__buf_16 _4358_ (.A(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__o2111ai_4 _4359_ (.A1(_1154_),
    .A2(_1161_),
    .B1(_1170_),
    .C1(_1174_),
    .D1(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__buf_6 _4360_ (.A(_1156_),
    .X(_1178_));
 sky130_fd_sc_hd__buf_6 _4361_ (.A(_1162_),
    .X(_1179_));
 sky130_fd_sc_hd__mux4_1 _4362_ (.A0(\registers[16][0] ),
    .A1(\registers[18][0] ),
    .A2(\registers[20][0] ),
    .A3(\registers[22][0] ),
    .S0(_1178_),
    .S1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__nor2_8 _4363_ (.A(_1165_),
    .B(_1175_),
    .Y(_1181_));
 sky130_fd_sc_hd__nor2_8 _4364_ (.A(_1153_),
    .B(_1175_),
    .Y(_1182_));
 sky130_fd_sc_hd__buf_8 _4365_ (.A(_1156_),
    .X(_1183_));
 sky130_fd_sc_hd__mux4_1 _4366_ (.A0(\registers[17][0] ),
    .A1(\registers[19][0] ),
    .A2(\registers[21][0] ),
    .A3(\registers[23][0] ),
    .S0(_1183_),
    .S1(_1179_),
    .X(_1184_));
 sky130_fd_sc_hd__a22oi_1 _4367_ (.A1(_1180_),
    .A2(_1181_),
    .B1(_1182_),
    .B2(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__nor2_4 _4368_ (.A(_1175_),
    .B(_1148_),
    .Y(_1186_));
 sky130_fd_sc_hd__buf_4 _4369_ (.A(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__mux4_1 _4370_ (.A0(\registers[0][0] ),
    .A1(\registers[1][0] ),
    .A2(\registers[2][0] ),
    .A3(\registers[3][0] ),
    .S0(_1165_),
    .S1(_1183_),
    .X(_1188_));
 sky130_fd_sc_hd__buf_6 _4371_ (.A(_1150_),
    .X(_1189_));
 sky130_fd_sc_hd__mux4_1 _4372_ (.A0(\registers[4][0] ),
    .A1(\registers[5][0] ),
    .A2(\registers[6][0] ),
    .A3(\registers[7][0] ),
    .S0(_1189_),
    .S1(_1178_),
    .X(_1190_));
 sky130_fd_sc_hd__buf_8 _4373_ (.A(_1158_),
    .X(_1191_));
 sky130_fd_sc_hd__buf_8 _4374_ (.A(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__mux2i_1 _4375_ (.A0(_1188_),
    .A1(_1190_),
    .S(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__nor2b_1 _4376_ (.A(_1148_),
    .B_N(net1),
    .Y(_1194_));
 sky130_fd_sc_hd__clkbuf_4 _4377_ (.A(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__clkbuf_16 _4378_ (.A(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__mux4_1 _4379_ (.A0(\registers[9][0] ),
    .A1(\registers[11][0] ),
    .A2(\registers[13][0] ),
    .A3(\registers[15][0] ),
    .S0(_1155_),
    .S1(_1159_),
    .X(_1197_));
 sky130_fd_sc_hd__mux4_1 _4380_ (.A0(\registers[8][0] ),
    .A1(\registers[10][0] ),
    .A2(\registers[12][0] ),
    .A3(\registers[14][0] ),
    .S0(_1155_),
    .S1(_1159_),
    .X(_1198_));
 sky130_fd_sc_hd__mux2i_1 _4381_ (.A0(_1197_),
    .A1(_1198_),
    .S(_1152_),
    .Y(_1199_));
 sky130_fd_sc_hd__nand2_4 _4382_ (.A(net3),
    .B(_1122_),
    .Y(_1200_));
 sky130_fd_sc_hd__buf_4 _4383_ (.A(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__a221o_2 _4384_ (.A1(_1187_),
    .A2(_1193_),
    .B1(_1196_),
    .B2(_1199_),
    .C1(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__a31oi_2 _4385_ (.A1(_1149_),
    .A2(_1177_),
    .A3(_1185_),
    .B1(_1202_),
    .Y(_0034_));
 sky130_fd_sc_hd__clkbuf_4 _4386_ (.A(_1152_),
    .X(_1203_));
 sky130_fd_sc_hd__buf_4 _4387_ (.A(_1166_),
    .X(_1204_));
 sky130_fd_sc_hd__buf_6 _4388_ (.A(_1162_),
    .X(_1205_));
 sky130_fd_sc_hd__mux4_1 _4389_ (.A0(\registers[17][10] ),
    .A1(\registers[19][10] ),
    .A2(\registers[21][10] ),
    .A3(\registers[23][10] ),
    .S0(_1204_),
    .S1(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__mux2i_1 _4390_ (.A0(\registers[18][10] ),
    .A1(\registers[22][10] ),
    .S(_1160_),
    .Y(_1207_));
 sky130_fd_sc_hd__mux2i_1 _4391_ (.A0(\registers[16][10] ),
    .A1(\registers[20][10] ),
    .S(_1179_),
    .Y(_1208_));
 sky130_fd_sc_hd__a221oi_1 _4392_ (.A1(_1173_),
    .A2(_1207_),
    .B1(_1208_),
    .B2(_1169_),
    .C1(_1176_),
    .Y(_1209_));
 sky130_fd_sc_hd__o21ai_1 _4393_ (.A1(_1203_),
    .A2(_1206_),
    .B1(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__mux4_1 _4394_ (.A0(\registers[24][10] ),
    .A1(\registers[26][10] ),
    .A2(\registers[28][10] ),
    .A3(\registers[30][10] ),
    .S0(_1178_),
    .S1(_1179_),
    .X(_1211_));
 sky130_fd_sc_hd__nor2b_4 _4395_ (.A(_1165_),
    .B_N(_1175_),
    .Y(_1212_));
 sky130_fd_sc_hd__and2_0 _4396_ (.A(_1165_),
    .B(_1175_),
    .X(_1213_));
 sky130_fd_sc_hd__clkbuf_4 _4397_ (.A(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__buf_6 _4398_ (.A(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__mux4_1 _4399_ (.A0(\registers[25][10] ),
    .A1(\registers[27][10] ),
    .A2(\registers[29][10] ),
    .A3(\registers[31][10] ),
    .S0(_1183_),
    .S1(_1179_),
    .X(_1216_));
 sky130_fd_sc_hd__a22oi_2 _4400_ (.A1(_1211_),
    .A2(_1212_),
    .B1(_1215_),
    .B2(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__mux4_1 _4401_ (.A0(\registers[0][10] ),
    .A1(\registers[1][10] ),
    .A2(\registers[2][10] ),
    .A3(\registers[3][10] ),
    .S0(_1165_),
    .S1(_1183_),
    .X(_1218_));
 sky130_fd_sc_hd__buf_6 _4402_ (.A(_1156_),
    .X(_1219_));
 sky130_fd_sc_hd__mux4_1 _4403_ (.A0(\registers[4][10] ),
    .A1(\registers[5][10] ),
    .A2(\registers[6][10] ),
    .A3(\registers[7][10] ),
    .S0(_1189_),
    .S1(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__mux2i_1 _4404_ (.A0(_1218_),
    .A1(_1220_),
    .S(_1192_),
    .Y(_1221_));
 sky130_fd_sc_hd__buf_8 _4405_ (.A(_1159_),
    .X(_1222_));
 sky130_fd_sc_hd__mux4_1 _4406_ (.A0(\registers[9][10] ),
    .A1(\registers[11][10] ),
    .A2(\registers[13][10] ),
    .A3(\registers[15][10] ),
    .S0(_1156_),
    .S1(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__buf_8 _4407_ (.A(_1155_),
    .X(_1224_));
 sky130_fd_sc_hd__buf_6 _4408_ (.A(_1159_),
    .X(_1225_));
 sky130_fd_sc_hd__mux4_1 _4409_ (.A0(\registers[8][10] ),
    .A1(\registers[10][10] ),
    .A2(\registers[12][10] ),
    .A3(\registers[14][10] ),
    .S0(_1224_),
    .S1(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__mux2i_1 _4410_ (.A0(_1223_),
    .A1(_1226_),
    .S(_1153_),
    .Y(_1227_));
 sky130_fd_sc_hd__buf_4 _4411_ (.A(_1195_),
    .X(_1228_));
 sky130_fd_sc_hd__a221o_2 _4412_ (.A1(_1187_),
    .A2(_1221_),
    .B1(_1227_),
    .B2(_1228_),
    .C1(_1201_),
    .X(_1229_));
 sky130_fd_sc_hd__a31oi_4 _4413_ (.A1(_1149_),
    .A2(_1210_),
    .A3(_1217_),
    .B1(_1229_),
    .Y(_0035_));
 sky130_fd_sc_hd__mux4_1 _4414_ (.A0(\registers[17][11] ),
    .A1(\registers[19][11] ),
    .A2(\registers[21][11] ),
    .A3(\registers[23][11] ),
    .S0(_1204_),
    .S1(_1205_),
    .X(_1230_));
 sky130_fd_sc_hd__buf_4 _4415_ (.A(_1172_),
    .X(_1231_));
 sky130_fd_sc_hd__buf_6 _4416_ (.A(_1159_),
    .X(_1232_));
 sky130_fd_sc_hd__mux2i_1 _4417_ (.A0(\registers[18][11] ),
    .A1(\registers[22][11] ),
    .S(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__mux2i_1 _4418_ (.A0(\registers[16][11] ),
    .A1(\registers[20][11] ),
    .S(_1179_),
    .Y(_1234_));
 sky130_fd_sc_hd__buf_4 _4419_ (.A(_1168_),
    .X(_1235_));
 sky130_fd_sc_hd__buf_4 _4420_ (.A(_1175_),
    .X(_1236_));
 sky130_fd_sc_hd__a221oi_2 _4421_ (.A1(_1231_),
    .A2(_1233_),
    .B1(_1234_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__o21ai_0 _4422_ (.A1(_1203_),
    .A2(_1230_),
    .B1(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__buf_6 _4423_ (.A(_1212_),
    .X(_1239_));
 sky130_fd_sc_hd__buf_6 _4424_ (.A(_1222_),
    .X(_1240_));
 sky130_fd_sc_hd__mux4_1 _4425_ (.A0(\registers[24][11] ),
    .A1(\registers[26][11] ),
    .A2(\registers[28][11] ),
    .A3(\registers[30][11] ),
    .S0(_1167_),
    .S1(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__buf_6 _4426_ (.A(_1166_),
    .X(_1242_));
 sky130_fd_sc_hd__buf_8 _4427_ (.A(_1162_),
    .X(_1243_));
 sky130_fd_sc_hd__mux4_1 _4428_ (.A0(\registers[25][11] ),
    .A1(\registers[27][11] ),
    .A2(\registers[29][11] ),
    .A3(\registers[31][11] ),
    .S0(_1242_),
    .S1(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__a22oi_2 _4429_ (.A1(_1239_),
    .A2(_1241_),
    .B1(_1244_),
    .B2(_1215_),
    .Y(_1245_));
 sky130_fd_sc_hd__mux4_1 _4430_ (.A0(\registers[0][11] ),
    .A1(\registers[1][11] ),
    .A2(\registers[2][11] ),
    .A3(\registers[3][11] ),
    .S0(_1165_),
    .S1(_1183_),
    .X(_1246_));
 sky130_fd_sc_hd__mux4_1 _4431_ (.A0(\registers[4][11] ),
    .A1(\registers[5][11] ),
    .A2(\registers[6][11] ),
    .A3(\registers[7][11] ),
    .S0(_1189_),
    .S1(_1219_),
    .X(_1247_));
 sky130_fd_sc_hd__buf_8 _4432_ (.A(_1222_),
    .X(_1248_));
 sky130_fd_sc_hd__mux2i_1 _4433_ (.A0(_1246_),
    .A1(_1247_),
    .S(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__mux4_1 _4434_ (.A0(\registers[9][11] ),
    .A1(\registers[11][11] ),
    .A2(\registers[13][11] ),
    .A3(\registers[15][11] ),
    .S0(_1156_),
    .S1(_1222_),
    .X(_1250_));
 sky130_fd_sc_hd__buf_6 _4435_ (.A(_1155_),
    .X(_1251_));
 sky130_fd_sc_hd__mux4_1 _4436_ (.A0(\registers[8][11] ),
    .A1(\registers[10][11] ),
    .A2(\registers[12][11] ),
    .A3(\registers[14][11] ),
    .S0(_1251_),
    .S1(_1225_),
    .X(_1252_));
 sky130_fd_sc_hd__mux2i_1 _4437_ (.A0(_1250_),
    .A1(_1252_),
    .S(_1153_),
    .Y(_1253_));
 sky130_fd_sc_hd__a221o_1 _4438_ (.A1(_1187_),
    .A2(_1249_),
    .B1(_1253_),
    .B2(_1228_),
    .C1(_1201_),
    .X(_1254_));
 sky130_fd_sc_hd__a31oi_2 _4439_ (.A1(_1149_),
    .A2(_1238_),
    .A3(_1245_),
    .B1(_1254_),
    .Y(_0036_));
 sky130_fd_sc_hd__mux4_1 _4440_ (.A0(\registers[25][12] ),
    .A1(\registers[27][12] ),
    .A2(\registers[29][12] ),
    .A3(\registers[31][12] ),
    .S0(_1157_),
    .S1(_1160_),
    .X(_1255_));
 sky130_fd_sc_hd__mux2i_1 _4441_ (.A0(\registers[24][12] ),
    .A1(\registers[28][12] ),
    .S(_1243_),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_1 _4442_ (.A(_1169_),
    .B(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__mux2i_1 _4443_ (.A0(\registers[26][12] ),
    .A1(\registers[30][12] ),
    .S(_1163_),
    .Y(_1258_));
 sky130_fd_sc_hd__nand2_1 _4444_ (.A(_1173_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__o2111ai_4 _4445_ (.A1(_1154_),
    .A2(_1255_),
    .B1(_1257_),
    .C1(_1259_),
    .D1(_1176_),
    .Y(_1260_));
 sky130_fd_sc_hd__mux4_1 _4446_ (.A0(\registers[16][12] ),
    .A1(\registers[18][12] ),
    .A2(\registers[20][12] ),
    .A3(\registers[22][12] ),
    .S0(_1167_),
    .S1(_1240_),
    .X(_1261_));
 sky130_fd_sc_hd__mux4_1 _4447_ (.A0(\registers[17][12] ),
    .A1(\registers[19][12] ),
    .A2(\registers[21][12] ),
    .A3(\registers[23][12] ),
    .S0(_1242_),
    .S1(_1243_),
    .X(_1262_));
 sky130_fd_sc_hd__a22oi_1 _4448_ (.A1(_1181_),
    .A2(_1261_),
    .B1(_1262_),
    .B2(_1182_),
    .Y(_1263_));
 sky130_fd_sc_hd__mux4_1 _4449_ (.A0(\registers[0][12] ),
    .A1(\registers[1][12] ),
    .A2(\registers[2][12] ),
    .A3(\registers[3][12] ),
    .S0(_1165_),
    .S1(_1183_),
    .X(_1264_));
 sky130_fd_sc_hd__buf_8 _4450_ (.A(_1150_),
    .X(_1265_));
 sky130_fd_sc_hd__mux4_1 _4451_ (.A0(\registers[4][12] ),
    .A1(\registers[5][12] ),
    .A2(\registers[6][12] ),
    .A3(\registers[7][12] ),
    .S0(_1265_),
    .S1(_1219_),
    .X(_1266_));
 sky130_fd_sc_hd__mux2i_1 _4452_ (.A0(_1264_),
    .A1(_1266_),
    .S(_1248_),
    .Y(_1267_));
 sky130_fd_sc_hd__buf_6 _4453_ (.A(_1155_),
    .X(_1268_));
 sky130_fd_sc_hd__mux4_1 _4454_ (.A0(\registers[9][12] ),
    .A1(\registers[11][12] ),
    .A2(\registers[13][12] ),
    .A3(\registers[15][12] ),
    .S0(_1268_),
    .S1(_1222_),
    .X(_1269_));
 sky130_fd_sc_hd__buf_4 _4455_ (.A(_1158_),
    .X(_1270_));
 sky130_fd_sc_hd__mux4_1 _4456_ (.A0(\registers[8][12] ),
    .A1(\registers[10][12] ),
    .A2(\registers[12][12] ),
    .A3(\registers[14][12] ),
    .S0(_1251_),
    .S1(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__mux2i_4 _4457_ (.A0(_1269_),
    .A1(_1271_),
    .S(_1153_),
    .Y(_1272_));
 sky130_fd_sc_hd__a221o_2 _4458_ (.A1(_1187_),
    .A2(_1267_),
    .B1(_1272_),
    .B2(_1228_),
    .C1(_1201_),
    .X(_1273_));
 sky130_fd_sc_hd__a31oi_2 _4459_ (.A1(_1149_),
    .A2(_1260_),
    .A3(_1263_),
    .B1(_1273_),
    .Y(_0037_));
 sky130_fd_sc_hd__buf_4 _4460_ (.A(_1162_),
    .X(_1274_));
 sky130_fd_sc_hd__mux4_1 _4461_ (.A0(\registers[17][13] ),
    .A1(\registers[19][13] ),
    .A2(\registers[21][13] ),
    .A3(\registers[23][13] ),
    .S0(_1204_),
    .S1(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__mux2i_1 _4462_ (.A0(\registers[18][13] ),
    .A1(\registers[22][13] ),
    .S(_1232_),
    .Y(_1276_));
 sky130_fd_sc_hd__mux2i_1 _4463_ (.A0(\registers[16][13] ),
    .A1(\registers[20][13] ),
    .S(_1179_),
    .Y(_1277_));
 sky130_fd_sc_hd__a221oi_1 _4464_ (.A1(_1231_),
    .A2(_1276_),
    .B1(_1277_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1278_));
 sky130_fd_sc_hd__o21ai_0 _4465_ (.A1(_1203_),
    .A2(_1275_),
    .B1(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__buf_6 _4466_ (.A(_1222_),
    .X(_1280_));
 sky130_fd_sc_hd__mux4_1 _4467_ (.A0(\registers[24][13] ),
    .A1(\registers[26][13] ),
    .A2(\registers[28][13] ),
    .A3(\registers[30][13] ),
    .S0(_1167_),
    .S1(_1280_),
    .X(_1281_));
 sky130_fd_sc_hd__buf_6 _4468_ (.A(_1162_),
    .X(_1282_));
 sky130_fd_sc_hd__mux4_1 _4469_ (.A0(\registers[25][13] ),
    .A1(\registers[27][13] ),
    .A2(\registers[29][13] ),
    .A3(\registers[31][13] ),
    .S0(_1242_),
    .S1(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__a22oi_2 _4470_ (.A1(_1239_),
    .A2(_1281_),
    .B1(_1283_),
    .B2(_1215_),
    .Y(_1284_));
 sky130_fd_sc_hd__mux4_1 _4471_ (.A0(\registers[0][13] ),
    .A1(\registers[1][13] ),
    .A2(\registers[2][13] ),
    .A3(\registers[3][13] ),
    .S0(_1165_),
    .S1(_1183_),
    .X(_1285_));
 sky130_fd_sc_hd__mux4_1 _4472_ (.A0(\registers[4][13] ),
    .A1(\registers[5][13] ),
    .A2(\registers[6][13] ),
    .A3(\registers[7][13] ),
    .S0(_1265_),
    .S1(_1219_),
    .X(_1286_));
 sky130_fd_sc_hd__mux2i_1 _4473_ (.A0(_1285_),
    .A1(_1286_),
    .S(_1248_),
    .Y(_1287_));
 sky130_fd_sc_hd__buf_6 _4474_ (.A(_1159_),
    .X(_1288_));
 sky130_fd_sc_hd__mux4_1 _4475_ (.A0(\registers[9][13] ),
    .A1(\registers[11][13] ),
    .A2(\registers[13][13] ),
    .A3(\registers[15][13] ),
    .S0(_1268_),
    .S1(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__mux4_1 _4476_ (.A0(\registers[8][13] ),
    .A1(\registers[10][13] ),
    .A2(\registers[12][13] ),
    .A3(\registers[14][13] ),
    .S0(_1251_),
    .S1(_1270_),
    .X(_1290_));
 sky130_fd_sc_hd__mux2i_4 _4477_ (.A0(_1289_),
    .A1(_1290_),
    .S(_1153_),
    .Y(_1291_));
 sky130_fd_sc_hd__a221o_1 _4478_ (.A1(_1187_),
    .A2(_1287_),
    .B1(_1291_),
    .B2(_1228_),
    .C1(_1201_),
    .X(_1292_));
 sky130_fd_sc_hd__a31oi_1 _4479_ (.A1(_1149_),
    .A2(_1279_),
    .A3(_1284_),
    .B1(_1292_),
    .Y(_0038_));
 sky130_fd_sc_hd__mux4_1 _4480_ (.A0(\registers[17][14] ),
    .A1(\registers[19][14] ),
    .A2(\registers[21][14] ),
    .A3(\registers[23][14] ),
    .S0(_1204_),
    .S1(_1274_),
    .X(_1293_));
 sky130_fd_sc_hd__mux2i_1 _4481_ (.A0(\registers[18][14] ),
    .A1(\registers[22][14] ),
    .S(_1232_),
    .Y(_1294_));
 sky130_fd_sc_hd__mux2i_1 _4482_ (.A0(\registers[16][14] ),
    .A1(\registers[20][14] ),
    .S(_1179_),
    .Y(_1295_));
 sky130_fd_sc_hd__a221oi_2 _4483_ (.A1(_1231_),
    .A2(_1294_),
    .B1(_1295_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1296_));
 sky130_fd_sc_hd__o21ai_0 _4484_ (.A1(_1203_),
    .A2(_1293_),
    .B1(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__mux4_1 _4485_ (.A0(\registers[24][14] ),
    .A1(\registers[26][14] ),
    .A2(\registers[28][14] ),
    .A3(\registers[30][14] ),
    .S0(_1167_),
    .S1(_1280_),
    .X(_1298_));
 sky130_fd_sc_hd__mux4_1 _4486_ (.A0(\registers[25][14] ),
    .A1(\registers[27][14] ),
    .A2(\registers[29][14] ),
    .A3(\registers[31][14] ),
    .S0(_1242_),
    .S1(_1282_),
    .X(_1299_));
 sky130_fd_sc_hd__a22oi_2 _4487_ (.A1(_1239_),
    .A2(_1298_),
    .B1(_1299_),
    .B2(_1215_),
    .Y(_1300_));
 sky130_fd_sc_hd__buf_16 _4488_ (.A(_1150_),
    .X(_1301_));
 sky130_fd_sc_hd__buf_16 _4489_ (.A(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__buf_6 _4490_ (.A(_1166_),
    .X(_1303_));
 sky130_fd_sc_hd__mux4_1 _4491_ (.A0(\registers[8][14] ),
    .A1(\registers[9][14] ),
    .A2(\registers[10][14] ),
    .A3(\registers[11][14] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__mux4_1 _4492_ (.A0(\registers[12][14] ),
    .A1(\registers[13][14] ),
    .A2(\registers[14][14] ),
    .A3(\registers[15][14] ),
    .S0(_1265_),
    .S1(_1219_),
    .X(_1305_));
 sky130_fd_sc_hd__mux2i_1 _4493_ (.A0(_1304_),
    .A1(_1305_),
    .S(_1248_),
    .Y(_1306_));
 sky130_fd_sc_hd__mux4_1 _4494_ (.A0(\registers[1][14] ),
    .A1(\registers[3][14] ),
    .A2(\registers[5][14] ),
    .A3(\registers[7][14] ),
    .S0(_1268_),
    .S1(_1288_),
    .X(_1307_));
 sky130_fd_sc_hd__mux4_1 _4495_ (.A0(\registers[0][14] ),
    .A1(\registers[2][14] ),
    .A2(\registers[4][14] ),
    .A3(\registers[6][14] ),
    .S0(_1251_),
    .S1(_1270_),
    .X(_1308_));
 sky130_fd_sc_hd__mux2i_1 _4496_ (.A0(_1307_),
    .A1(_1308_),
    .S(_1153_),
    .Y(_1309_));
 sky130_fd_sc_hd__buf_8 _4497_ (.A(_1186_),
    .X(_1310_));
 sky130_fd_sc_hd__a221o_2 _4498_ (.A1(_1196_),
    .A2(_1306_),
    .B1(_1309_),
    .B2(_1310_),
    .C1(_1201_),
    .X(_1311_));
 sky130_fd_sc_hd__a31oi_1 _4499_ (.A1(_1149_),
    .A2(_1297_),
    .A3(_1300_),
    .B1(_1311_),
    .Y(_0039_));
 sky130_fd_sc_hd__mux4_1 _4500_ (.A0(\registers[17][15] ),
    .A1(\registers[19][15] ),
    .A2(\registers[21][15] ),
    .A3(\registers[23][15] ),
    .S0(_1204_),
    .S1(_1274_),
    .X(_1312_));
 sky130_fd_sc_hd__mux2i_1 _4501_ (.A0(\registers[18][15] ),
    .A1(\registers[22][15] ),
    .S(_1232_),
    .Y(_1313_));
 sky130_fd_sc_hd__mux2i_1 _4502_ (.A0(\registers[16][15] ),
    .A1(\registers[20][15] ),
    .S(_1179_),
    .Y(_1314_));
 sky130_fd_sc_hd__a221oi_2 _4503_ (.A1(_1231_),
    .A2(_1313_),
    .B1(_1314_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1315_));
 sky130_fd_sc_hd__o21ai_0 _4504_ (.A1(_1203_),
    .A2(_1312_),
    .B1(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__mux4_1 _4505_ (.A0(\registers[24][15] ),
    .A1(\registers[26][15] ),
    .A2(\registers[28][15] ),
    .A3(\registers[30][15] ),
    .S0(_1167_),
    .S1(_1280_),
    .X(_1317_));
 sky130_fd_sc_hd__mux4_1 _4506_ (.A0(\registers[25][15] ),
    .A1(\registers[27][15] ),
    .A2(\registers[29][15] ),
    .A3(\registers[31][15] ),
    .S0(_1242_),
    .S1(_1282_),
    .X(_1318_));
 sky130_fd_sc_hd__a22oi_2 _4507_ (.A1(_1239_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_1215_),
    .Y(_1319_));
 sky130_fd_sc_hd__mux4_1 _4508_ (.A0(\registers[0][15] ),
    .A1(\registers[1][15] ),
    .A2(\registers[2][15] ),
    .A3(\registers[3][15] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1320_));
 sky130_fd_sc_hd__mux4_1 _4509_ (.A0(\registers[4][15] ),
    .A1(\registers[5][15] ),
    .A2(\registers[6][15] ),
    .A3(\registers[7][15] ),
    .S0(_1265_),
    .S1(_1219_),
    .X(_1321_));
 sky130_fd_sc_hd__mux2i_1 _4510_ (.A0(_1320_),
    .A1(_1321_),
    .S(_1248_),
    .Y(_1322_));
 sky130_fd_sc_hd__mux4_1 _4511_ (.A0(\registers[9][15] ),
    .A1(\registers[11][15] ),
    .A2(\registers[13][15] ),
    .A3(\registers[15][15] ),
    .S0(_1268_),
    .S1(_1288_),
    .X(_1323_));
 sky130_fd_sc_hd__mux4_1 _4512_ (.A0(\registers[8][15] ),
    .A1(\registers[10][15] ),
    .A2(\registers[12][15] ),
    .A3(\registers[14][15] ),
    .S0(_1251_),
    .S1(_1270_),
    .X(_1324_));
 sky130_fd_sc_hd__mux2i_2 _4513_ (.A0(_1323_),
    .A1(_1324_),
    .S(_1153_),
    .Y(_1325_));
 sky130_fd_sc_hd__a221o_2 _4514_ (.A1(_1187_),
    .A2(_1322_),
    .B1(_1325_),
    .B2(_1228_),
    .C1(_1201_),
    .X(_1326_));
 sky130_fd_sc_hd__a31oi_1 _4515_ (.A1(_1149_),
    .A2(_1316_),
    .A3(_1319_),
    .B1(_1326_),
    .Y(_0040_));
 sky130_fd_sc_hd__mux4_1 _4516_ (.A0(\registers[17][16] ),
    .A1(\registers[19][16] ),
    .A2(\registers[21][16] ),
    .A3(\registers[23][16] ),
    .S0(_1204_),
    .S1(_1274_),
    .X(_1327_));
 sky130_fd_sc_hd__mux2i_1 _4517_ (.A0(\registers[18][16] ),
    .A1(\registers[22][16] ),
    .S(_1232_),
    .Y(_1328_));
 sky130_fd_sc_hd__buf_6 _4518_ (.A(_1222_),
    .X(_1329_));
 sky130_fd_sc_hd__mux2i_1 _4519_ (.A0(\registers[16][16] ),
    .A1(\registers[20][16] ),
    .S(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__a221oi_1 _4520_ (.A1(_1231_),
    .A2(_1328_),
    .B1(_1330_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1331_));
 sky130_fd_sc_hd__o21ai_0 _4521_ (.A1(_1203_),
    .A2(_1327_),
    .B1(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__mux4_1 _4522_ (.A0(\registers[24][16] ),
    .A1(\registers[26][16] ),
    .A2(\registers[28][16] ),
    .A3(\registers[30][16] ),
    .S0(_1167_),
    .S1(_1280_),
    .X(_1333_));
 sky130_fd_sc_hd__mux4_1 _4523_ (.A0(\registers[25][16] ),
    .A1(\registers[27][16] ),
    .A2(\registers[29][16] ),
    .A3(\registers[31][16] ),
    .S0(_1242_),
    .S1(_1282_),
    .X(_1334_));
 sky130_fd_sc_hd__a22oi_2 _4524_ (.A1(_1239_),
    .A2(_1333_),
    .B1(_1334_),
    .B2(_1215_),
    .Y(_1335_));
 sky130_fd_sc_hd__mux4_1 _4525_ (.A0(\registers[0][16] ),
    .A1(\registers[1][16] ),
    .A2(\registers[2][16] ),
    .A3(\registers[3][16] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1336_));
 sky130_fd_sc_hd__mux4_1 _4526_ (.A0(\registers[4][16] ),
    .A1(\registers[5][16] ),
    .A2(\registers[6][16] ),
    .A3(\registers[7][16] ),
    .S0(_1265_),
    .S1(_1219_),
    .X(_1337_));
 sky130_fd_sc_hd__mux2i_1 _4527_ (.A0(_1336_),
    .A1(_1337_),
    .S(_1248_),
    .Y(_1338_));
 sky130_fd_sc_hd__mux4_1 _4528_ (.A0(\registers[9][16] ),
    .A1(\registers[11][16] ),
    .A2(\registers[13][16] ),
    .A3(\registers[15][16] ),
    .S0(_1268_),
    .S1(_1288_),
    .X(_1339_));
 sky130_fd_sc_hd__mux4_1 _4529_ (.A0(\registers[8][16] ),
    .A1(\registers[10][16] ),
    .A2(\registers[12][16] ),
    .A3(\registers[14][16] ),
    .S0(_1251_),
    .S1(_1270_),
    .X(_1340_));
 sky130_fd_sc_hd__buf_16 _4530_ (.A(_1152_),
    .X(_1341_));
 sky130_fd_sc_hd__mux2i_4 _4531_ (.A0(_1339_),
    .A1(_1340_),
    .S(_1341_),
    .Y(_1342_));
 sky130_fd_sc_hd__a221o_2 _4532_ (.A1(_1187_),
    .A2(_1338_),
    .B1(_1342_),
    .B2(_1228_),
    .C1(_1201_),
    .X(_1343_));
 sky130_fd_sc_hd__a31oi_1 _4533_ (.A1(_1149_),
    .A2(_1332_),
    .A3(_1335_),
    .B1(_1343_),
    .Y(_0041_));
 sky130_fd_sc_hd__mux4_1 _4534_ (.A0(\registers[25][17] ),
    .A1(\registers[27][17] ),
    .A2(\registers[29][17] ),
    .A3(\registers[31][17] ),
    .S0(_1157_),
    .S1(_1160_),
    .X(_1344_));
 sky130_fd_sc_hd__mux2i_1 _4535_ (.A0(\registers[24][17] ),
    .A1(\registers[28][17] ),
    .S(_1243_),
    .Y(_1345_));
 sky130_fd_sc_hd__nand2_1 _4536_ (.A(_1169_),
    .B(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__mux2i_1 _4537_ (.A0(\registers[26][17] ),
    .A1(\registers[30][17] ),
    .S(_1163_),
    .Y(_1347_));
 sky130_fd_sc_hd__nand2_1 _4538_ (.A(_1173_),
    .B(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__o2111ai_4 _4539_ (.A1(_1154_),
    .A2(_1344_),
    .B1(_1346_),
    .C1(_1348_),
    .D1(_1176_),
    .Y(_1349_));
 sky130_fd_sc_hd__mux4_1 _4540_ (.A0(\registers[16][17] ),
    .A1(\registers[18][17] ),
    .A2(\registers[20][17] ),
    .A3(\registers[22][17] ),
    .S0(_1167_),
    .S1(_1280_),
    .X(_1350_));
 sky130_fd_sc_hd__mux4_1 _4541_ (.A0(\registers[17][17] ),
    .A1(\registers[19][17] ),
    .A2(\registers[21][17] ),
    .A3(\registers[23][17] ),
    .S0(_1242_),
    .S1(_1282_),
    .X(_1351_));
 sky130_fd_sc_hd__a22oi_1 _4542_ (.A1(_1181_),
    .A2(_1350_),
    .B1(_1351_),
    .B2(_1182_),
    .Y(_1352_));
 sky130_fd_sc_hd__mux4_1 _4543_ (.A0(\registers[8][17] ),
    .A1(\registers[9][17] ),
    .A2(\registers[10][17] ),
    .A3(\registers[11][17] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1353_));
 sky130_fd_sc_hd__mux4_1 _4544_ (.A0(\registers[12][17] ),
    .A1(\registers[13][17] ),
    .A2(\registers[14][17] ),
    .A3(\registers[15][17] ),
    .S0(_1265_),
    .S1(_1219_),
    .X(_1354_));
 sky130_fd_sc_hd__mux2i_2 _4545_ (.A0(_1353_),
    .A1(_1354_),
    .S(_1248_),
    .Y(_1355_));
 sky130_fd_sc_hd__mux4_1 _4546_ (.A0(\registers[1][17] ),
    .A1(\registers[3][17] ),
    .A2(\registers[5][17] ),
    .A3(\registers[7][17] ),
    .S0(_1268_),
    .S1(_1288_),
    .X(_1356_));
 sky130_fd_sc_hd__mux4_1 _4547_ (.A0(\registers[0][17] ),
    .A1(\registers[2][17] ),
    .A2(\registers[4][17] ),
    .A3(\registers[6][17] ),
    .S0(_1251_),
    .S1(_1270_),
    .X(_1357_));
 sky130_fd_sc_hd__mux2i_1 _4548_ (.A0(_1356_),
    .A1(_1357_),
    .S(_1341_),
    .Y(_1358_));
 sky130_fd_sc_hd__a221o_2 _4549_ (.A1(_1196_),
    .A2(_1355_),
    .B1(_1358_),
    .B2(_1310_),
    .C1(_1201_),
    .X(_1359_));
 sky130_fd_sc_hd__a31oi_2 _4550_ (.A1(_1149_),
    .A2(_1349_),
    .A3(_1352_),
    .B1(_1359_),
    .Y(_0042_));
 sky130_fd_sc_hd__mux4_1 _4551_ (.A0(\registers[17][18] ),
    .A1(\registers[19][18] ),
    .A2(\registers[21][18] ),
    .A3(\registers[23][18] ),
    .S0(_1204_),
    .S1(_1274_),
    .X(_1360_));
 sky130_fd_sc_hd__mux2i_1 _4552_ (.A0(\registers[18][18] ),
    .A1(\registers[22][18] ),
    .S(_1232_),
    .Y(_1361_));
 sky130_fd_sc_hd__mux2i_1 _4553_ (.A0(\registers[16][18] ),
    .A1(\registers[20][18] ),
    .S(_1329_),
    .Y(_1362_));
 sky130_fd_sc_hd__a221oi_1 _4554_ (.A1(_1231_),
    .A2(_1361_),
    .B1(_1362_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1363_));
 sky130_fd_sc_hd__o21ai_0 _4555_ (.A1(_1203_),
    .A2(_1360_),
    .B1(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__buf_8 _4556_ (.A(_1156_),
    .X(_1365_));
 sky130_fd_sc_hd__mux4_1 _4557_ (.A0(\registers[24][18] ),
    .A1(\registers[26][18] ),
    .A2(\registers[28][18] ),
    .A3(\registers[30][18] ),
    .S0(_1365_),
    .S1(_1280_),
    .X(_1366_));
 sky130_fd_sc_hd__mux4_1 _4558_ (.A0(\registers[25][18] ),
    .A1(\registers[27][18] ),
    .A2(\registers[29][18] ),
    .A3(\registers[31][18] ),
    .S0(_1242_),
    .S1(_1282_),
    .X(_1367_));
 sky130_fd_sc_hd__a22oi_2 _4559_ (.A1(_1239_),
    .A2(_1366_),
    .B1(_1367_),
    .B2(_1215_),
    .Y(_1368_));
 sky130_fd_sc_hd__mux4_1 _4560_ (.A0(\registers[0][18] ),
    .A1(\registers[1][18] ),
    .A2(\registers[2][18] ),
    .A3(\registers[3][18] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1369_));
 sky130_fd_sc_hd__mux4_1 _4561_ (.A0(\registers[4][18] ),
    .A1(\registers[5][18] ),
    .A2(\registers[6][18] ),
    .A3(\registers[7][18] ),
    .S0(_1265_),
    .S1(_1219_),
    .X(_1370_));
 sky130_fd_sc_hd__mux2i_1 _4562_ (.A0(_1369_),
    .A1(_1370_),
    .S(_1248_),
    .Y(_1371_));
 sky130_fd_sc_hd__mux4_1 _4563_ (.A0(\registers[9][18] ),
    .A1(\registers[11][18] ),
    .A2(\registers[13][18] ),
    .A3(\registers[15][18] ),
    .S0(_1268_),
    .S1(_1288_),
    .X(_1372_));
 sky130_fd_sc_hd__mux4_1 _4564_ (.A0(\registers[8][18] ),
    .A1(\registers[10][18] ),
    .A2(\registers[12][18] ),
    .A3(\registers[14][18] ),
    .S0(_1251_),
    .S1(_1270_),
    .X(_1373_));
 sky130_fd_sc_hd__mux2i_4 _4565_ (.A0(_1372_),
    .A1(_1373_),
    .S(_1341_),
    .Y(_1374_));
 sky130_fd_sc_hd__a221o_1 _4566_ (.A1(_1187_),
    .A2(_1371_),
    .B1(_1374_),
    .B2(_1228_),
    .C1(_1201_),
    .X(_1375_));
 sky130_fd_sc_hd__a31oi_1 _4567_ (.A1(_1149_),
    .A2(_1364_),
    .A3(_1368_),
    .B1(_1375_),
    .Y(_0043_));
 sky130_fd_sc_hd__buf_6 _4568_ (.A(_1148_),
    .X(_1376_));
 sky130_fd_sc_hd__mux4_1 _4569_ (.A0(\registers[25][19] ),
    .A1(\registers[27][19] ),
    .A2(\registers[29][19] ),
    .A3(\registers[31][19] ),
    .S0(_1157_),
    .S1(_1160_),
    .X(_1377_));
 sky130_fd_sc_hd__mux2i_1 _4570_ (.A0(\registers[24][19] ),
    .A1(\registers[28][19] ),
    .S(_1243_),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _4571_ (.A(_1169_),
    .B(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__mux2i_1 _4572_ (.A0(\registers[26][19] ),
    .A1(\registers[30][19] ),
    .S(_1163_),
    .Y(_1380_));
 sky130_fd_sc_hd__nand2_1 _4573_ (.A(_1173_),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__o2111ai_4 _4574_ (.A1(_1154_),
    .A2(_1377_),
    .B1(_1379_),
    .C1(_1381_),
    .D1(_1176_),
    .Y(_1382_));
 sky130_fd_sc_hd__mux4_1 _4575_ (.A0(\registers[16][19] ),
    .A1(\registers[18][19] ),
    .A2(\registers[20][19] ),
    .A3(\registers[22][19] ),
    .S0(_1365_),
    .S1(_1280_),
    .X(_1383_));
 sky130_fd_sc_hd__mux4_1 _4576_ (.A0(\registers[17][19] ),
    .A1(\registers[19][19] ),
    .A2(\registers[21][19] ),
    .A3(\registers[23][19] ),
    .S0(_1242_),
    .S1(_1282_),
    .X(_1384_));
 sky130_fd_sc_hd__a22oi_1 _4577_ (.A1(_1181_),
    .A2(_1383_),
    .B1(_1384_),
    .B2(_1182_),
    .Y(_1385_));
 sky130_fd_sc_hd__mux4_1 _4578_ (.A0(\registers[0][19] ),
    .A1(\registers[1][19] ),
    .A2(\registers[2][19] ),
    .A3(\registers[3][19] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1386_));
 sky130_fd_sc_hd__mux4_1 _4579_ (.A0(\registers[4][19] ),
    .A1(\registers[5][19] ),
    .A2(\registers[6][19] ),
    .A3(\registers[7][19] ),
    .S0(_1265_),
    .S1(_1219_),
    .X(_1387_));
 sky130_fd_sc_hd__mux2i_1 _4580_ (.A0(_1386_),
    .A1(_1387_),
    .S(_1248_),
    .Y(_1388_));
 sky130_fd_sc_hd__mux4_1 _4581_ (.A0(\registers[9][19] ),
    .A1(\registers[11][19] ),
    .A2(\registers[13][19] ),
    .A3(\registers[15][19] ),
    .S0(_1268_),
    .S1(_1288_),
    .X(_1389_));
 sky130_fd_sc_hd__mux4_1 _4582_ (.A0(\registers[8][19] ),
    .A1(\registers[10][19] ),
    .A2(\registers[12][19] ),
    .A3(\registers[14][19] ),
    .S0(_1251_),
    .S1(_1270_),
    .X(_1390_));
 sky130_fd_sc_hd__mux2i_4 _4583_ (.A0(_1389_),
    .A1(_1390_),
    .S(_1341_),
    .Y(_1391_));
 sky130_fd_sc_hd__buf_6 _4584_ (.A(_1200_),
    .X(_1392_));
 sky130_fd_sc_hd__a221o_2 _4585_ (.A1(_1187_),
    .A2(_1388_),
    .B1(_1391_),
    .B2(_1228_),
    .C1(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__a31oi_2 _4586_ (.A1(_1376_),
    .A2(_1382_),
    .A3(_1385_),
    .B1(_1393_),
    .Y(_0044_));
 sky130_fd_sc_hd__mux4_1 _4587_ (.A0(\registers[25][1] ),
    .A1(\registers[27][1] ),
    .A2(\registers[29][1] ),
    .A3(\registers[31][1] ),
    .S0(_1157_),
    .S1(_1160_),
    .X(_1394_));
 sky130_fd_sc_hd__mux2i_1 _4588_ (.A0(\registers[24][1] ),
    .A1(\registers[28][1] ),
    .S(_1243_),
    .Y(_1395_));
 sky130_fd_sc_hd__nand2_1 _4589_ (.A(_1169_),
    .B(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__mux2i_1 _4590_ (.A0(\registers[26][1] ),
    .A1(\registers[30][1] ),
    .S(_1163_),
    .Y(_1397_));
 sky130_fd_sc_hd__nand2_1 _4591_ (.A(_1173_),
    .B(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__o2111ai_4 _4592_ (.A1(_1154_),
    .A2(_1394_),
    .B1(_1396_),
    .C1(_1398_),
    .D1(_1176_),
    .Y(_1399_));
 sky130_fd_sc_hd__mux4_1 _4593_ (.A0(\registers[16][1] ),
    .A1(\registers[18][1] ),
    .A2(\registers[20][1] ),
    .A3(\registers[22][1] ),
    .S0(_1365_),
    .S1(_1280_),
    .X(_1400_));
 sky130_fd_sc_hd__mux4_1 _4594_ (.A0(\registers[17][1] ),
    .A1(\registers[19][1] ),
    .A2(\registers[21][1] ),
    .A3(\registers[23][1] ),
    .S0(_1242_),
    .S1(_1282_),
    .X(_1401_));
 sky130_fd_sc_hd__a22oi_2 _4595_ (.A1(_1181_),
    .A2(_1400_),
    .B1(_1401_),
    .B2(_1182_),
    .Y(_1402_));
 sky130_fd_sc_hd__mux4_1 _4596_ (.A0(\registers[0][1] ),
    .A1(\registers[1][1] ),
    .A2(\registers[2][1] ),
    .A3(\registers[3][1] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1403_));
 sky130_fd_sc_hd__buf_6 _4597_ (.A(_1156_),
    .X(_1404_));
 sky130_fd_sc_hd__mux4_1 _4598_ (.A0(\registers[4][1] ),
    .A1(\registers[5][1] ),
    .A2(\registers[6][1] ),
    .A3(\registers[7][1] ),
    .S0(_1265_),
    .S1(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2i_1 _4599_ (.A0(_1403_),
    .A1(_1405_),
    .S(_1248_),
    .Y(_1406_));
 sky130_fd_sc_hd__mux4_1 _4600_ (.A0(\registers[9][1] ),
    .A1(\registers[11][1] ),
    .A2(\registers[13][1] ),
    .A3(\registers[15][1] ),
    .S0(_1268_),
    .S1(_1288_),
    .X(_1407_));
 sky130_fd_sc_hd__mux4_1 _4601_ (.A0(\registers[8][1] ),
    .A1(\registers[10][1] ),
    .A2(\registers[12][1] ),
    .A3(\registers[14][1] ),
    .S0(_1251_),
    .S1(_1270_),
    .X(_1408_));
 sky130_fd_sc_hd__mux2i_4 _4602_ (.A0(_1407_),
    .A1(_1408_),
    .S(_1341_),
    .Y(_1409_));
 sky130_fd_sc_hd__a221o_4 _4603_ (.A1(_1187_),
    .A2(_1406_),
    .B1(_1409_),
    .B2(_1228_),
    .C1(_1392_),
    .X(_1410_));
 sky130_fd_sc_hd__a31oi_4 _4604_ (.A1(_1376_),
    .A2(_1399_),
    .A3(_1402_),
    .B1(_1410_),
    .Y(_0045_));
 sky130_fd_sc_hd__mux4_1 _4605_ (.A0(\registers[17][20] ),
    .A1(\registers[19][20] ),
    .A2(\registers[21][20] ),
    .A3(\registers[23][20] ),
    .S0(_1204_),
    .S1(_1274_),
    .X(_1411_));
 sky130_fd_sc_hd__mux2i_1 _4606_ (.A0(\registers[18][20] ),
    .A1(\registers[22][20] ),
    .S(_1232_),
    .Y(_1412_));
 sky130_fd_sc_hd__mux2i_1 _4607_ (.A0(\registers[16][20] ),
    .A1(\registers[20][20] ),
    .S(_1329_),
    .Y(_1413_));
 sky130_fd_sc_hd__a221oi_2 _4608_ (.A1(_1231_),
    .A2(_1412_),
    .B1(_1413_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1414_));
 sky130_fd_sc_hd__o21ai_1 _4609_ (.A1(_1203_),
    .A2(_1411_),
    .B1(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__mux4_1 _4610_ (.A0(\registers[24][20] ),
    .A1(\registers[26][20] ),
    .A2(\registers[28][20] ),
    .A3(\registers[30][20] ),
    .S0(_1365_),
    .S1(_1280_),
    .X(_1416_));
 sky130_fd_sc_hd__buf_8 _4611_ (.A(_1166_),
    .X(_1417_));
 sky130_fd_sc_hd__mux4_1 _4612_ (.A0(\registers[25][20] ),
    .A1(\registers[27][20] ),
    .A2(\registers[29][20] ),
    .A3(\registers[31][20] ),
    .S0(_1417_),
    .S1(_1282_),
    .X(_1418_));
 sky130_fd_sc_hd__a22oi_2 _4613_ (.A1(_1239_),
    .A2(_1416_),
    .B1(_1418_),
    .B2(_1215_),
    .Y(_1419_));
 sky130_fd_sc_hd__buf_6 _4614_ (.A(_1186_),
    .X(_1420_));
 sky130_fd_sc_hd__mux4_1 _4615_ (.A0(\registers[0][20] ),
    .A1(\registers[1][20] ),
    .A2(\registers[2][20] ),
    .A3(\registers[3][20] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1421_));
 sky130_fd_sc_hd__mux4_1 _4616_ (.A0(\registers[4][20] ),
    .A1(\registers[5][20] ),
    .A2(\registers[6][20] ),
    .A3(\registers[7][20] ),
    .S0(_1265_),
    .S1(_1404_),
    .X(_1422_));
 sky130_fd_sc_hd__buf_8 _4617_ (.A(_1222_),
    .X(_1423_));
 sky130_fd_sc_hd__mux2i_1 _4618_ (.A0(_1421_),
    .A1(_1422_),
    .S(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__mux4_1 _4619_ (.A0(\registers[9][20] ),
    .A1(\registers[11][20] ),
    .A2(\registers[13][20] ),
    .A3(\registers[15][20] ),
    .S0(_1268_),
    .S1(_1288_),
    .X(_1425_));
 sky130_fd_sc_hd__buf_8 _4620_ (.A(_1155_),
    .X(_1426_));
 sky130_fd_sc_hd__mux4_1 _4621_ (.A0(\registers[8][20] ),
    .A1(\registers[10][20] ),
    .A2(\registers[12][20] ),
    .A3(\registers[14][20] ),
    .S0(_1426_),
    .S1(_1270_),
    .X(_1427_));
 sky130_fd_sc_hd__mux2i_4 _4622_ (.A0(_1425_),
    .A1(_1427_),
    .S(_1341_),
    .Y(_1428_));
 sky130_fd_sc_hd__buf_6 _4623_ (.A(_1195_),
    .X(_1429_));
 sky130_fd_sc_hd__a221o_2 _4624_ (.A1(_1420_),
    .A2(_1424_),
    .B1(_1428_),
    .B2(_1429_),
    .C1(_1392_),
    .X(_1430_));
 sky130_fd_sc_hd__a31oi_2 _4625_ (.A1(_1376_),
    .A2(_1415_),
    .A3(_1419_),
    .B1(_1430_),
    .Y(_0046_));
 sky130_fd_sc_hd__mux4_1 _4626_ (.A0(\registers[17][21] ),
    .A1(\registers[19][21] ),
    .A2(\registers[21][21] ),
    .A3(\registers[23][21] ),
    .S0(_1204_),
    .S1(_1274_),
    .X(_1431_));
 sky130_fd_sc_hd__mux2i_1 _4627_ (.A0(\registers[18][21] ),
    .A1(\registers[22][21] ),
    .S(_1232_),
    .Y(_1432_));
 sky130_fd_sc_hd__mux2i_1 _4628_ (.A0(\registers[16][21] ),
    .A1(\registers[20][21] ),
    .S(_1329_),
    .Y(_1433_));
 sky130_fd_sc_hd__a221oi_2 _4629_ (.A1(_1231_),
    .A2(_1432_),
    .B1(_1433_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1434_));
 sky130_fd_sc_hd__o21ai_1 _4630_ (.A1(_1203_),
    .A2(_1431_),
    .B1(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__mux4_1 _4631_ (.A0(\registers[24][21] ),
    .A1(\registers[26][21] ),
    .A2(\registers[28][21] ),
    .A3(\registers[30][21] ),
    .S0(_1365_),
    .S1(_1280_),
    .X(_1436_));
 sky130_fd_sc_hd__mux4_1 _4632_ (.A0(\registers[25][21] ),
    .A1(\registers[27][21] ),
    .A2(\registers[29][21] ),
    .A3(\registers[31][21] ),
    .S0(_1417_),
    .S1(_1282_),
    .X(_1437_));
 sky130_fd_sc_hd__a22oi_2 _4633_ (.A1(_1239_),
    .A2(_1436_),
    .B1(_1437_),
    .B2(_1215_),
    .Y(_1438_));
 sky130_fd_sc_hd__mux4_1 _4634_ (.A0(\registers[8][21] ),
    .A1(\registers[9][21] ),
    .A2(\registers[10][21] ),
    .A3(\registers[11][21] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1439_));
 sky130_fd_sc_hd__buf_6 _4635_ (.A(_1150_),
    .X(_1440_));
 sky130_fd_sc_hd__mux4_1 _4636_ (.A0(\registers[12][21] ),
    .A1(\registers[13][21] ),
    .A2(\registers[14][21] ),
    .A3(\registers[15][21] ),
    .S0(_1440_),
    .S1(_1404_),
    .X(_1441_));
 sky130_fd_sc_hd__mux2i_2 _4637_ (.A0(_1439_),
    .A1(_1441_),
    .S(_1423_),
    .Y(_1442_));
 sky130_fd_sc_hd__buf_6 _4638_ (.A(_1155_),
    .X(_1443_));
 sky130_fd_sc_hd__mux4_1 _4639_ (.A0(\registers[1][21] ),
    .A1(\registers[3][21] ),
    .A2(\registers[5][21] ),
    .A3(\registers[7][21] ),
    .S0(_1443_),
    .S1(_1288_),
    .X(_1444_));
 sky130_fd_sc_hd__buf_6 _4640_ (.A(_1158_),
    .X(_1445_));
 sky130_fd_sc_hd__mux4_1 _4641_ (.A0(\registers[0][21] ),
    .A1(\registers[2][21] ),
    .A2(\registers[4][21] ),
    .A3(\registers[6][21] ),
    .S0(_1426_),
    .S1(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__mux2i_1 _4642_ (.A0(_1444_),
    .A1(_1446_),
    .S(_1341_),
    .Y(_1447_));
 sky130_fd_sc_hd__a221o_4 _4643_ (.A1(_1196_),
    .A2(_1442_),
    .B1(_1447_),
    .B2(_1310_),
    .C1(_1392_),
    .X(_1448_));
 sky130_fd_sc_hd__a31oi_4 _4644_ (.A1(_1376_),
    .A2(_1435_),
    .A3(_1438_),
    .B1(_1448_),
    .Y(_0047_));
 sky130_fd_sc_hd__mux4_1 _4645_ (.A0(\registers[17][22] ),
    .A1(\registers[19][22] ),
    .A2(\registers[21][22] ),
    .A3(\registers[23][22] ),
    .S0(_1204_),
    .S1(_1274_),
    .X(_1449_));
 sky130_fd_sc_hd__mux2i_1 _4646_ (.A0(\registers[18][22] ),
    .A1(\registers[22][22] ),
    .S(_1232_),
    .Y(_1450_));
 sky130_fd_sc_hd__mux2i_1 _4647_ (.A0(\registers[16][22] ),
    .A1(\registers[20][22] ),
    .S(_1329_),
    .Y(_1451_));
 sky130_fd_sc_hd__a221oi_2 _4648_ (.A1(_1231_),
    .A2(_1450_),
    .B1(_1451_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1452_));
 sky130_fd_sc_hd__o21ai_0 _4649_ (.A1(_1203_),
    .A2(_1449_),
    .B1(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__buf_6 _4650_ (.A(_1222_),
    .X(_1454_));
 sky130_fd_sc_hd__mux4_1 _4651_ (.A0(\registers[24][22] ),
    .A1(\registers[26][22] ),
    .A2(\registers[28][22] ),
    .A3(\registers[30][22] ),
    .S0(_1365_),
    .S1(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__buf_6 _4652_ (.A(_1162_),
    .X(_1456_));
 sky130_fd_sc_hd__mux4_1 _4653_ (.A0(\registers[25][22] ),
    .A1(\registers[27][22] ),
    .A2(\registers[29][22] ),
    .A3(\registers[31][22] ),
    .S0(_1417_),
    .S1(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__a22oi_2 _4654_ (.A1(_1239_),
    .A2(_1455_),
    .B1(_1457_),
    .B2(_1215_),
    .Y(_1458_));
 sky130_fd_sc_hd__mux4_1 _4655_ (.A0(\registers[0][22] ),
    .A1(\registers[1][22] ),
    .A2(\registers[2][22] ),
    .A3(\registers[3][22] ),
    .S0(_1302_),
    .S1(_1303_),
    .X(_1459_));
 sky130_fd_sc_hd__mux4_1 _4656_ (.A0(\registers[4][22] ),
    .A1(\registers[5][22] ),
    .A2(\registers[6][22] ),
    .A3(\registers[7][22] ),
    .S0(_1440_),
    .S1(_1404_),
    .X(_1460_));
 sky130_fd_sc_hd__mux2i_1 _4657_ (.A0(_1459_),
    .A1(_1460_),
    .S(_1423_),
    .Y(_1461_));
 sky130_fd_sc_hd__buf_6 _4658_ (.A(_1159_),
    .X(_1462_));
 sky130_fd_sc_hd__mux4_1 _4659_ (.A0(\registers[9][22] ),
    .A1(\registers[11][22] ),
    .A2(\registers[13][22] ),
    .A3(\registers[15][22] ),
    .S0(_1443_),
    .S1(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__mux4_1 _4660_ (.A0(\registers[8][22] ),
    .A1(\registers[10][22] ),
    .A2(\registers[12][22] ),
    .A3(\registers[14][22] ),
    .S0(_1426_),
    .S1(_1445_),
    .X(_1464_));
 sky130_fd_sc_hd__mux2i_2 _4661_ (.A0(_1463_),
    .A1(_1464_),
    .S(_1341_),
    .Y(_1465_));
 sky130_fd_sc_hd__a221o_2 _4662_ (.A1(_1420_),
    .A2(_1461_),
    .B1(_1465_),
    .B2(_1429_),
    .C1(_1392_),
    .X(_1466_));
 sky130_fd_sc_hd__a31oi_2 _4663_ (.A1(_1376_),
    .A2(_1453_),
    .A3(_1458_),
    .B1(_1466_),
    .Y(_0048_));
 sky130_fd_sc_hd__clkbuf_4 _4664_ (.A(_1151_),
    .X(_1467_));
 sky130_fd_sc_hd__buf_4 _4665_ (.A(_1166_),
    .X(_1468_));
 sky130_fd_sc_hd__mux4_1 _4666_ (.A0(\registers[17][23] ),
    .A1(\registers[19][23] ),
    .A2(\registers[21][23] ),
    .A3(\registers[23][23] ),
    .S0(_1468_),
    .S1(_1274_),
    .X(_1469_));
 sky130_fd_sc_hd__mux2i_1 _4667_ (.A0(\registers[18][23] ),
    .A1(\registers[22][23] ),
    .S(_1232_),
    .Y(_1470_));
 sky130_fd_sc_hd__mux2i_1 _4668_ (.A0(\registers[16][23] ),
    .A1(\registers[20][23] ),
    .S(_1329_),
    .Y(_1471_));
 sky130_fd_sc_hd__a221oi_2 _4669_ (.A1(_1231_),
    .A2(_1470_),
    .B1(_1471_),
    .B2(_1235_),
    .C1(_1236_),
    .Y(_1472_));
 sky130_fd_sc_hd__o21ai_1 _4670_ (.A1(_1467_),
    .A2(_1469_),
    .B1(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__mux4_1 _4671_ (.A0(\registers[24][23] ),
    .A1(\registers[26][23] ),
    .A2(\registers[28][23] ),
    .A3(\registers[30][23] ),
    .S0(_1365_),
    .S1(_1454_),
    .X(_1474_));
 sky130_fd_sc_hd__mux4_1 _4672_ (.A0(\registers[25][23] ),
    .A1(\registers[27][23] ),
    .A2(\registers[29][23] ),
    .A3(\registers[31][23] ),
    .S0(_1417_),
    .S1(_1456_),
    .X(_1475_));
 sky130_fd_sc_hd__buf_8 _4673_ (.A(_1214_),
    .X(_1476_));
 sky130_fd_sc_hd__a22oi_4 _4674_ (.A1(_1239_),
    .A2(_1474_),
    .B1(_1475_),
    .B2(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__buf_6 _4675_ (.A(_1150_),
    .X(_1478_));
 sky130_fd_sc_hd__buf_6 _4676_ (.A(_1166_),
    .X(_1479_));
 sky130_fd_sc_hd__mux4_1 _4677_ (.A0(\registers[8][23] ),
    .A1(\registers[9][23] ),
    .A2(\registers[10][23] ),
    .A3(\registers[11][23] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__mux4_1 _4678_ (.A0(\registers[12][23] ),
    .A1(\registers[13][23] ),
    .A2(\registers[14][23] ),
    .A3(\registers[15][23] ),
    .S0(_1440_),
    .S1(_1404_),
    .X(_1481_));
 sky130_fd_sc_hd__mux2i_2 _4679_ (.A0(_1480_),
    .A1(_1481_),
    .S(_1423_),
    .Y(_1482_));
 sky130_fd_sc_hd__mux4_1 _4680_ (.A0(\registers[1][23] ),
    .A1(\registers[3][23] ),
    .A2(\registers[5][23] ),
    .A3(\registers[7][23] ),
    .S0(_1443_),
    .S1(_1462_),
    .X(_1483_));
 sky130_fd_sc_hd__mux4_1 _4681_ (.A0(\registers[0][23] ),
    .A1(\registers[2][23] ),
    .A2(\registers[4][23] ),
    .A3(\registers[6][23] ),
    .S0(_1426_),
    .S1(_1445_),
    .X(_1484_));
 sky130_fd_sc_hd__mux2i_1 _4682_ (.A0(_1483_),
    .A1(_1484_),
    .S(_1341_),
    .Y(_1485_));
 sky130_fd_sc_hd__a221o_4 _4683_ (.A1(_1196_),
    .A2(_1482_),
    .B1(_1485_),
    .B2(_1310_),
    .C1(_1392_),
    .X(_1486_));
 sky130_fd_sc_hd__a31oi_4 _4684_ (.A1(_1376_),
    .A2(_1473_),
    .A3(_1477_),
    .B1(_1486_),
    .Y(_0049_));
 sky130_fd_sc_hd__mux4_1 _4685_ (.A0(\registers[17][24] ),
    .A1(\registers[19][24] ),
    .A2(\registers[21][24] ),
    .A3(\registers[23][24] ),
    .S0(_1468_),
    .S1(_1274_),
    .X(_1487_));
 sky130_fd_sc_hd__buf_4 _4686_ (.A(_1172_),
    .X(_1488_));
 sky130_fd_sc_hd__buf_6 _4687_ (.A(_1159_),
    .X(_1489_));
 sky130_fd_sc_hd__mux2i_1 _4688_ (.A0(\registers[18][24] ),
    .A1(\registers[22][24] ),
    .S(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__mux2i_1 _4689_ (.A0(\registers[16][24] ),
    .A1(\registers[20][24] ),
    .S(_1329_),
    .Y(_1491_));
 sky130_fd_sc_hd__buf_4 _4690_ (.A(_1168_),
    .X(_1492_));
 sky130_fd_sc_hd__buf_4 _4691_ (.A(_1175_),
    .X(_1493_));
 sky130_fd_sc_hd__a221oi_2 _4692_ (.A1(_1488_),
    .A2(_1490_),
    .B1(_1491_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__o21ai_1 _4693_ (.A1(_1467_),
    .A2(_1487_),
    .B1(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__buf_8 _4694_ (.A(_1212_),
    .X(_1496_));
 sky130_fd_sc_hd__mux4_1 _4695_ (.A0(\registers[24][24] ),
    .A1(\registers[26][24] ),
    .A2(\registers[28][24] ),
    .A3(\registers[30][24] ),
    .S0(_1365_),
    .S1(_1454_),
    .X(_1497_));
 sky130_fd_sc_hd__mux4_1 _4696_ (.A0(\registers[25][24] ),
    .A1(\registers[27][24] ),
    .A2(\registers[29][24] ),
    .A3(\registers[31][24] ),
    .S0(_1417_),
    .S1(_1456_),
    .X(_1498_));
 sky130_fd_sc_hd__a22oi_4 _4697_ (.A1(_1496_),
    .A2(_1497_),
    .B1(_1498_),
    .B2(_1476_),
    .Y(_1499_));
 sky130_fd_sc_hd__mux4_1 _4698_ (.A0(\registers[8][24] ),
    .A1(\registers[9][24] ),
    .A2(\registers[10][24] ),
    .A3(\registers[11][24] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1500_));
 sky130_fd_sc_hd__mux4_1 _4699_ (.A0(\registers[12][24] ),
    .A1(\registers[13][24] ),
    .A2(\registers[14][24] ),
    .A3(\registers[15][24] ),
    .S0(_1440_),
    .S1(_1404_),
    .X(_1501_));
 sky130_fd_sc_hd__mux2i_4 _4700_ (.A0(_1500_),
    .A1(_1501_),
    .S(_1423_),
    .Y(_1502_));
 sky130_fd_sc_hd__mux4_1 _4701_ (.A0(\registers[1][24] ),
    .A1(\registers[3][24] ),
    .A2(\registers[5][24] ),
    .A3(\registers[7][24] ),
    .S0(_1443_),
    .S1(_1462_),
    .X(_1503_));
 sky130_fd_sc_hd__mux4_1 _4702_ (.A0(\registers[0][24] ),
    .A1(\registers[2][24] ),
    .A2(\registers[4][24] ),
    .A3(\registers[6][24] ),
    .S0(_1426_),
    .S1(_1445_),
    .X(_1504_));
 sky130_fd_sc_hd__mux2i_1 _4703_ (.A0(_1503_),
    .A1(_1504_),
    .S(_1341_),
    .Y(_1505_));
 sky130_fd_sc_hd__a221o_4 _4704_ (.A1(_1196_),
    .A2(_1502_),
    .B1(_1505_),
    .B2(_1310_),
    .C1(_1392_),
    .X(_1506_));
 sky130_fd_sc_hd__a31oi_4 _4705_ (.A1(_1376_),
    .A2(_1495_),
    .A3(_1499_),
    .B1(_1506_),
    .Y(_0050_));
 sky130_fd_sc_hd__mux4_1 _4706_ (.A0(\registers[25][25] ),
    .A1(\registers[27][25] ),
    .A2(\registers[29][25] ),
    .A3(\registers[31][25] ),
    .S0(_1157_),
    .S1(_1160_),
    .X(_1507_));
 sky130_fd_sc_hd__mux2i_1 _4707_ (.A0(\registers[24][25] ),
    .A1(\registers[28][25] ),
    .S(_1243_),
    .Y(_1508_));
 sky130_fd_sc_hd__nand2_1 _4708_ (.A(_1169_),
    .B(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__mux2i_1 _4709_ (.A0(\registers[26][25] ),
    .A1(\registers[30][25] ),
    .S(_1163_),
    .Y(_1510_));
 sky130_fd_sc_hd__nand2_1 _4710_ (.A(_1173_),
    .B(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__o2111ai_4 _4711_ (.A1(_1154_),
    .A2(_1507_),
    .B1(_1509_),
    .C1(_1511_),
    .D1(_1176_),
    .Y(_1512_));
 sky130_fd_sc_hd__mux4_1 _4712_ (.A0(\registers[16][25] ),
    .A1(\registers[18][25] ),
    .A2(\registers[20][25] ),
    .A3(\registers[22][25] ),
    .S0(_1365_),
    .S1(_1454_),
    .X(_1513_));
 sky130_fd_sc_hd__mux4_1 _4713_ (.A0(\registers[17][25] ),
    .A1(\registers[19][25] ),
    .A2(\registers[21][25] ),
    .A3(\registers[23][25] ),
    .S0(_1417_),
    .S1(_1456_),
    .X(_1514_));
 sky130_fd_sc_hd__a22oi_1 _4714_ (.A1(_1181_),
    .A2(_1513_),
    .B1(_1514_),
    .B2(_1182_),
    .Y(_1515_));
 sky130_fd_sc_hd__mux4_1 _4715_ (.A0(\registers[0][25] ),
    .A1(\registers[1][25] ),
    .A2(\registers[2][25] ),
    .A3(\registers[3][25] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1516_));
 sky130_fd_sc_hd__mux4_1 _4716_ (.A0(\registers[4][25] ),
    .A1(\registers[5][25] ),
    .A2(\registers[6][25] ),
    .A3(\registers[7][25] ),
    .S0(_1440_),
    .S1(_1404_),
    .X(_1517_));
 sky130_fd_sc_hd__mux2i_1 _4717_ (.A0(_1516_),
    .A1(_1517_),
    .S(_1423_),
    .Y(_1518_));
 sky130_fd_sc_hd__mux4_1 _4718_ (.A0(\registers[9][25] ),
    .A1(\registers[11][25] ),
    .A2(\registers[13][25] ),
    .A3(\registers[15][25] ),
    .S0(_1443_),
    .S1(_1462_),
    .X(_1519_));
 sky130_fd_sc_hd__mux4_1 _4719_ (.A0(\registers[8][25] ),
    .A1(\registers[10][25] ),
    .A2(\registers[12][25] ),
    .A3(\registers[14][25] ),
    .S0(_1426_),
    .S1(_1445_),
    .X(_1520_));
 sky130_fd_sc_hd__buf_8 _4720_ (.A(_1152_),
    .X(_1521_));
 sky130_fd_sc_hd__mux2i_2 _4721_ (.A0(_1519_),
    .A1(_1520_),
    .S(_1521_),
    .Y(_1522_));
 sky130_fd_sc_hd__a221o_4 _4722_ (.A1(_1420_),
    .A2(_1518_),
    .B1(_1522_),
    .B2(_1429_),
    .C1(_1392_),
    .X(_1523_));
 sky130_fd_sc_hd__a31oi_2 _4723_ (.A1(_1376_),
    .A2(_1512_),
    .A3(_1515_),
    .B1(_1523_),
    .Y(_0051_));
 sky130_fd_sc_hd__buf_4 _4724_ (.A(_1162_),
    .X(_1524_));
 sky130_fd_sc_hd__mux4_1 _4725_ (.A0(\registers[17][26] ),
    .A1(\registers[19][26] ),
    .A2(\registers[21][26] ),
    .A3(\registers[23][26] ),
    .S0(_1468_),
    .S1(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__mux2i_1 _4726_ (.A0(\registers[18][26] ),
    .A1(\registers[22][26] ),
    .S(_1489_),
    .Y(_1526_));
 sky130_fd_sc_hd__mux2i_1 _4727_ (.A0(\registers[16][26] ),
    .A1(\registers[20][26] ),
    .S(_1329_),
    .Y(_1527_));
 sky130_fd_sc_hd__a221oi_2 _4728_ (.A1(_1488_),
    .A2(_1526_),
    .B1(_1527_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1528_));
 sky130_fd_sc_hd__o21ai_1 _4729_ (.A1(_1467_),
    .A2(_1525_),
    .B1(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__mux4_1 _4730_ (.A0(\registers[24][26] ),
    .A1(\registers[26][26] ),
    .A2(\registers[28][26] ),
    .A3(\registers[30][26] ),
    .S0(_1365_),
    .S1(_1454_),
    .X(_1530_));
 sky130_fd_sc_hd__mux4_1 _4731_ (.A0(\registers[25][26] ),
    .A1(\registers[27][26] ),
    .A2(\registers[29][26] ),
    .A3(\registers[31][26] ),
    .S0(_1417_),
    .S1(_1456_),
    .X(_1531_));
 sky130_fd_sc_hd__a22oi_4 _4732_ (.A1(_1496_),
    .A2(_1530_),
    .B1(_1531_),
    .B2(_1476_),
    .Y(_1532_));
 sky130_fd_sc_hd__mux4_1 _4733_ (.A0(\registers[0][26] ),
    .A1(\registers[1][26] ),
    .A2(\registers[2][26] ),
    .A3(\registers[3][26] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1533_));
 sky130_fd_sc_hd__mux4_1 _4734_ (.A0(\registers[4][26] ),
    .A1(\registers[5][26] ),
    .A2(\registers[6][26] ),
    .A3(\registers[7][26] ),
    .S0(_1440_),
    .S1(_1404_),
    .X(_1534_));
 sky130_fd_sc_hd__mux2i_1 _4735_ (.A0(_1533_),
    .A1(_1534_),
    .S(_1423_),
    .Y(_1535_));
 sky130_fd_sc_hd__mux4_1 _4736_ (.A0(\registers[9][26] ),
    .A1(\registers[11][26] ),
    .A2(\registers[13][26] ),
    .A3(\registers[15][26] ),
    .S0(_1443_),
    .S1(_1462_),
    .X(_1536_));
 sky130_fd_sc_hd__mux4_1 _4737_ (.A0(\registers[8][26] ),
    .A1(\registers[10][26] ),
    .A2(\registers[12][26] ),
    .A3(\registers[14][26] ),
    .S0(_1426_),
    .S1(_1445_),
    .X(_1537_));
 sky130_fd_sc_hd__mux2i_4 _4738_ (.A0(_1536_),
    .A1(_1537_),
    .S(_1521_),
    .Y(_1538_));
 sky130_fd_sc_hd__a221o_4 _4739_ (.A1(_1420_),
    .A2(_1535_),
    .B1(_1538_),
    .B2(_1429_),
    .C1(_1392_),
    .X(_1539_));
 sky130_fd_sc_hd__a31oi_4 _4740_ (.A1(_1376_),
    .A2(_1529_),
    .A3(_1532_),
    .B1(_1539_),
    .Y(_0052_));
 sky130_fd_sc_hd__mux4_1 _4741_ (.A0(\registers[25][27] ),
    .A1(\registers[27][27] ),
    .A2(\registers[29][27] ),
    .A3(\registers[31][27] ),
    .S0(_1157_),
    .S1(_1160_),
    .X(_1540_));
 sky130_fd_sc_hd__mux2i_1 _4742_ (.A0(\registers[24][27] ),
    .A1(\registers[28][27] ),
    .S(_1243_),
    .Y(_1541_));
 sky130_fd_sc_hd__nand2_1 _4743_ (.A(_1169_),
    .B(_1541_),
    .Y(_1542_));
 sky130_fd_sc_hd__mux2i_1 _4744_ (.A0(\registers[26][27] ),
    .A1(\registers[30][27] ),
    .S(_1163_),
    .Y(_1543_));
 sky130_fd_sc_hd__nand2_1 _4745_ (.A(_1173_),
    .B(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__o2111ai_4 _4746_ (.A1(_1154_),
    .A2(_1540_),
    .B1(_1542_),
    .C1(_1544_),
    .D1(_1176_),
    .Y(_1545_));
 sky130_fd_sc_hd__buf_6 _4747_ (.A(_1156_),
    .X(_1546_));
 sky130_fd_sc_hd__mux4_1 _4748_ (.A0(\registers[16][27] ),
    .A1(\registers[18][27] ),
    .A2(\registers[20][27] ),
    .A3(\registers[22][27] ),
    .S0(_1546_),
    .S1(_1454_),
    .X(_1547_));
 sky130_fd_sc_hd__mux4_1 _4749_ (.A0(\registers[17][27] ),
    .A1(\registers[19][27] ),
    .A2(\registers[21][27] ),
    .A3(\registers[23][27] ),
    .S0(_1417_),
    .S1(_1456_),
    .X(_1548_));
 sky130_fd_sc_hd__a22oi_2 _4750_ (.A1(_1181_),
    .A2(_1547_),
    .B1(_1548_),
    .B2(_1182_),
    .Y(_1549_));
 sky130_fd_sc_hd__mux4_1 _4751_ (.A0(\registers[0][27] ),
    .A1(\registers[1][27] ),
    .A2(\registers[2][27] ),
    .A3(\registers[3][27] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1550_));
 sky130_fd_sc_hd__mux4_1 _4752_ (.A0(\registers[4][27] ),
    .A1(\registers[5][27] ),
    .A2(\registers[6][27] ),
    .A3(\registers[7][27] ),
    .S0(_1440_),
    .S1(_1404_),
    .X(_1551_));
 sky130_fd_sc_hd__mux2i_1 _4753_ (.A0(_1550_),
    .A1(_1551_),
    .S(_1423_),
    .Y(_1552_));
 sky130_fd_sc_hd__mux4_1 _4754_ (.A0(\registers[9][27] ),
    .A1(\registers[11][27] ),
    .A2(\registers[13][27] ),
    .A3(\registers[15][27] ),
    .S0(_1443_),
    .S1(_1462_),
    .X(_1553_));
 sky130_fd_sc_hd__mux4_1 _4755_ (.A0(\registers[8][27] ),
    .A1(\registers[10][27] ),
    .A2(\registers[12][27] ),
    .A3(\registers[14][27] ),
    .S0(_1426_),
    .S1(_1445_),
    .X(_1554_));
 sky130_fd_sc_hd__mux2i_2 _4756_ (.A0(_1553_),
    .A1(_1554_),
    .S(_1521_),
    .Y(_1555_));
 sky130_fd_sc_hd__a221o_4 _4757_ (.A1(_1420_),
    .A2(_1552_),
    .B1(_1555_),
    .B2(_1429_),
    .C1(_1392_),
    .X(_1556_));
 sky130_fd_sc_hd__a31oi_4 _4758_ (.A1(_1376_),
    .A2(_1545_),
    .A3(_1549_),
    .B1(_1556_),
    .Y(_0053_));
 sky130_fd_sc_hd__buf_4 _4759_ (.A(_1148_),
    .X(_1557_));
 sky130_fd_sc_hd__mux4_1 _4760_ (.A0(\registers[17][28] ),
    .A1(\registers[19][28] ),
    .A2(\registers[21][28] ),
    .A3(\registers[23][28] ),
    .S0(_1468_),
    .S1(_1524_),
    .X(_1558_));
 sky130_fd_sc_hd__mux2i_1 _4761_ (.A0(\registers[18][28] ),
    .A1(\registers[22][28] ),
    .S(_1489_),
    .Y(_1559_));
 sky130_fd_sc_hd__mux2i_1 _4762_ (.A0(\registers[16][28] ),
    .A1(\registers[20][28] ),
    .S(_1329_),
    .Y(_1560_));
 sky130_fd_sc_hd__a221oi_1 _4763_ (.A1(_1488_),
    .A2(_1559_),
    .B1(_1560_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1561_));
 sky130_fd_sc_hd__o21ai_0 _4764_ (.A1(_1467_),
    .A2(_1558_),
    .B1(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__mux4_1 _4765_ (.A0(\registers[24][28] ),
    .A1(\registers[26][28] ),
    .A2(\registers[28][28] ),
    .A3(\registers[30][28] ),
    .S0(_1546_),
    .S1(_1454_),
    .X(_1563_));
 sky130_fd_sc_hd__mux4_1 _4766_ (.A0(\registers[25][28] ),
    .A1(\registers[27][28] ),
    .A2(\registers[29][28] ),
    .A3(\registers[31][28] ),
    .S0(_1417_),
    .S1(_1456_),
    .X(_1564_));
 sky130_fd_sc_hd__a22oi_4 _4767_ (.A1(_1496_),
    .A2(_1563_),
    .B1(_1564_),
    .B2(_1476_),
    .Y(_1565_));
 sky130_fd_sc_hd__mux4_1 _4768_ (.A0(\registers[0][28] ),
    .A1(\registers[1][28] ),
    .A2(\registers[2][28] ),
    .A3(\registers[3][28] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1566_));
 sky130_fd_sc_hd__mux4_1 _4769_ (.A0(\registers[4][28] ),
    .A1(\registers[5][28] ),
    .A2(\registers[6][28] ),
    .A3(\registers[7][28] ),
    .S0(_1440_),
    .S1(_1404_),
    .X(_1567_));
 sky130_fd_sc_hd__mux2i_1 _4770_ (.A0(_1566_),
    .A1(_1567_),
    .S(_1423_),
    .Y(_1568_));
 sky130_fd_sc_hd__mux4_1 _4771_ (.A0(\registers[9][28] ),
    .A1(\registers[11][28] ),
    .A2(\registers[13][28] ),
    .A3(\registers[15][28] ),
    .S0(_1443_),
    .S1(_1462_),
    .X(_1569_));
 sky130_fd_sc_hd__mux4_1 _4772_ (.A0(\registers[8][28] ),
    .A1(\registers[10][28] ),
    .A2(\registers[12][28] ),
    .A3(\registers[14][28] ),
    .S0(_1426_),
    .S1(_1445_),
    .X(_1570_));
 sky130_fd_sc_hd__mux2i_2 _4773_ (.A0(_1569_),
    .A1(_1570_),
    .S(_1521_),
    .Y(_1571_));
 sky130_fd_sc_hd__buf_4 _4774_ (.A(_1200_),
    .X(_1572_));
 sky130_fd_sc_hd__a221o_2 _4775_ (.A1(_1420_),
    .A2(_1568_),
    .B1(_1571_),
    .B2(_1429_),
    .C1(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__a31oi_1 _4776_ (.A1(_1557_),
    .A2(_1562_),
    .A3(_1565_),
    .B1(_1573_),
    .Y(_0054_));
 sky130_fd_sc_hd__mux4_1 _4777_ (.A0(\registers[17][29] ),
    .A1(\registers[19][29] ),
    .A2(\registers[21][29] ),
    .A3(\registers[23][29] ),
    .S0(_1468_),
    .S1(_1524_),
    .X(_1574_));
 sky130_fd_sc_hd__mux2i_1 _4778_ (.A0(\registers[18][29] ),
    .A1(\registers[22][29] ),
    .S(_1489_),
    .Y(_1575_));
 sky130_fd_sc_hd__mux2i_1 _4779_ (.A0(\registers[16][29] ),
    .A1(\registers[20][29] ),
    .S(_1329_),
    .Y(_1576_));
 sky130_fd_sc_hd__a221oi_2 _4780_ (.A1(_1488_),
    .A2(_1575_),
    .B1(_1576_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1577_));
 sky130_fd_sc_hd__o21ai_0 _4781_ (.A1(_1467_),
    .A2(_1574_),
    .B1(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__mux4_1 _4782_ (.A0(\registers[24][29] ),
    .A1(\registers[26][29] ),
    .A2(\registers[28][29] ),
    .A3(\registers[30][29] ),
    .S0(_1546_),
    .S1(_1454_),
    .X(_1579_));
 sky130_fd_sc_hd__mux4_1 _4783_ (.A0(\registers[25][29] ),
    .A1(\registers[27][29] ),
    .A2(\registers[29][29] ),
    .A3(\registers[31][29] ),
    .S0(_1417_),
    .S1(_1456_),
    .X(_1580_));
 sky130_fd_sc_hd__a22oi_4 _4784_ (.A1(_1496_),
    .A2(_1579_),
    .B1(_1580_),
    .B2(_1476_),
    .Y(_1581_));
 sky130_fd_sc_hd__mux4_1 _4785_ (.A0(\registers[8][29] ),
    .A1(\registers[9][29] ),
    .A2(\registers[10][29] ),
    .A3(\registers[11][29] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1582_));
 sky130_fd_sc_hd__buf_6 _4786_ (.A(_1156_),
    .X(_1583_));
 sky130_fd_sc_hd__mux4_1 _4787_ (.A0(\registers[12][29] ),
    .A1(\registers[13][29] ),
    .A2(\registers[14][29] ),
    .A3(\registers[15][29] ),
    .S0(_1440_),
    .S1(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__mux2i_2 _4788_ (.A0(_1582_),
    .A1(_1584_),
    .S(_1423_),
    .Y(_1585_));
 sky130_fd_sc_hd__mux4_1 _4789_ (.A0(\registers[1][29] ),
    .A1(\registers[3][29] ),
    .A2(\registers[5][29] ),
    .A3(\registers[7][29] ),
    .S0(_1443_),
    .S1(_1462_),
    .X(_1586_));
 sky130_fd_sc_hd__mux4_1 _4790_ (.A0(\registers[0][29] ),
    .A1(\registers[2][29] ),
    .A2(\registers[4][29] ),
    .A3(\registers[6][29] ),
    .S0(_1426_),
    .S1(_1445_),
    .X(_1587_));
 sky130_fd_sc_hd__mux2i_1 _4791_ (.A0(_1586_),
    .A1(_1587_),
    .S(_1521_),
    .Y(_1588_));
 sky130_fd_sc_hd__a221o_2 _4792_ (.A1(_1196_),
    .A2(_1585_),
    .B1(_1588_),
    .B2(_1310_),
    .C1(_1572_),
    .X(_1589_));
 sky130_fd_sc_hd__a31oi_2 _4793_ (.A1(_1557_),
    .A2(_1578_),
    .A3(_1581_),
    .B1(_1589_),
    .Y(_0055_));
 sky130_fd_sc_hd__mux4_1 _4794_ (.A0(\registers[17][2] ),
    .A1(\registers[19][2] ),
    .A2(\registers[21][2] ),
    .A3(\registers[23][2] ),
    .S0(_1468_),
    .S1(_1524_),
    .X(_1590_));
 sky130_fd_sc_hd__mux2i_1 _4795_ (.A0(\registers[18][2] ),
    .A1(\registers[22][2] ),
    .S(_1489_),
    .Y(_1591_));
 sky130_fd_sc_hd__mux2i_1 _4796_ (.A0(\registers[16][2] ),
    .A1(\registers[20][2] ),
    .S(_1240_),
    .Y(_1592_));
 sky130_fd_sc_hd__a221oi_1 _4797_ (.A1(_1488_),
    .A2(_1591_),
    .B1(_1592_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1593_));
 sky130_fd_sc_hd__o21ai_0 _4798_ (.A1(_1467_),
    .A2(_1590_),
    .B1(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__mux4_1 _4799_ (.A0(\registers[24][2] ),
    .A1(\registers[26][2] ),
    .A2(\registers[28][2] ),
    .A3(\registers[30][2] ),
    .S0(_1546_),
    .S1(_1454_),
    .X(_1595_));
 sky130_fd_sc_hd__buf_6 _4800_ (.A(_1166_),
    .X(_1596_));
 sky130_fd_sc_hd__mux4_1 _4801_ (.A0(\registers[25][2] ),
    .A1(\registers[27][2] ),
    .A2(\registers[29][2] ),
    .A3(\registers[31][2] ),
    .S0(_1596_),
    .S1(_1456_),
    .X(_1597_));
 sky130_fd_sc_hd__a22oi_4 _4802_ (.A1(_1496_),
    .A2(_1595_),
    .B1(_1597_),
    .B2(_1476_),
    .Y(_1598_));
 sky130_fd_sc_hd__mux4_1 _4803_ (.A0(\registers[0][2] ),
    .A1(\registers[1][2] ),
    .A2(\registers[2][2] ),
    .A3(\registers[3][2] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1599_));
 sky130_fd_sc_hd__mux4_1 _4804_ (.A0(\registers[4][2] ),
    .A1(\registers[5][2] ),
    .A2(\registers[6][2] ),
    .A3(\registers[7][2] ),
    .S0(_1440_),
    .S1(_1583_),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_16 _4805_ (.A(_1222_),
    .X(_1601_));
 sky130_fd_sc_hd__mux2i_1 _4806_ (.A0(_1599_),
    .A1(_1600_),
    .S(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__mux4_1 _4807_ (.A0(\registers[9][2] ),
    .A1(\registers[11][2] ),
    .A2(\registers[13][2] ),
    .A3(\registers[15][2] ),
    .S0(_1443_),
    .S1(_1462_),
    .X(_1603_));
 sky130_fd_sc_hd__buf_8 _4808_ (.A(_1155_),
    .X(_1604_));
 sky130_fd_sc_hd__mux4_1 _4809_ (.A0(\registers[8][2] ),
    .A1(\registers[10][2] ),
    .A2(\registers[12][2] ),
    .A3(\registers[14][2] ),
    .S0(_1604_),
    .S1(_1445_),
    .X(_1605_));
 sky130_fd_sc_hd__mux2i_2 _4810_ (.A0(_1603_),
    .A1(_1605_),
    .S(_1521_),
    .Y(_1606_));
 sky130_fd_sc_hd__a221o_2 _4811_ (.A1(_1420_),
    .A2(_1602_),
    .B1(_1606_),
    .B2(_1429_),
    .C1(_1572_),
    .X(_1607_));
 sky130_fd_sc_hd__a31oi_1 _4812_ (.A1(_1557_),
    .A2(_1594_),
    .A3(_1598_),
    .B1(_1607_),
    .Y(_0056_));
 sky130_fd_sc_hd__mux4_1 _4813_ (.A0(\registers[17][30] ),
    .A1(\registers[19][30] ),
    .A2(\registers[21][30] ),
    .A3(\registers[23][30] ),
    .S0(_1468_),
    .S1(_1524_),
    .X(_1608_));
 sky130_fd_sc_hd__mux2i_2 _4814_ (.A0(\registers[18][30] ),
    .A1(\registers[22][30] ),
    .S(_1489_),
    .Y(_1609_));
 sky130_fd_sc_hd__mux2i_1 _4815_ (.A0(\registers[16][30] ),
    .A1(\registers[20][30] ),
    .S(_1240_),
    .Y(_1610_));
 sky130_fd_sc_hd__a221oi_2 _4816_ (.A1(_1488_),
    .A2(_1609_),
    .B1(_1610_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1611_));
 sky130_fd_sc_hd__o21ai_0 _4817_ (.A1(_1467_),
    .A2(_1608_),
    .B1(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__mux4_1 _4818_ (.A0(\registers[24][30] ),
    .A1(\registers[26][30] ),
    .A2(\registers[28][30] ),
    .A3(\registers[30][30] ),
    .S0(_1546_),
    .S1(_1454_),
    .X(_1613_));
 sky130_fd_sc_hd__mux4_1 _4819_ (.A0(\registers[25][30] ),
    .A1(\registers[27][30] ),
    .A2(\registers[29][30] ),
    .A3(\registers[31][30] ),
    .S0(_1596_),
    .S1(_1456_),
    .X(_1614_));
 sky130_fd_sc_hd__a22oi_2 _4820_ (.A1(_1496_),
    .A2(_1613_),
    .B1(_1614_),
    .B2(_1476_),
    .Y(_1615_));
 sky130_fd_sc_hd__mux4_1 _4821_ (.A0(\registers[8][30] ),
    .A1(\registers[9][30] ),
    .A2(\registers[10][30] ),
    .A3(\registers[11][30] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1616_));
 sky130_fd_sc_hd__mux4_1 _4822_ (.A0(\registers[12][30] ),
    .A1(\registers[13][30] ),
    .A2(\registers[14][30] ),
    .A3(\registers[15][30] ),
    .S0(_1301_),
    .S1(_1583_),
    .X(_1617_));
 sky130_fd_sc_hd__mux2i_2 _4823_ (.A0(_1616_),
    .A1(_1617_),
    .S(_1601_),
    .Y(_1618_));
 sky130_fd_sc_hd__mux4_1 _4824_ (.A0(\registers[1][30] ),
    .A1(\registers[3][30] ),
    .A2(\registers[5][30] ),
    .A3(\registers[7][30] ),
    .S0(_1224_),
    .S1(_1462_),
    .X(_1619_));
 sky130_fd_sc_hd__mux4_1 _4825_ (.A0(\registers[0][30] ),
    .A1(\registers[2][30] ),
    .A2(\registers[4][30] ),
    .A3(\registers[6][30] ),
    .S0(_1604_),
    .S1(_1191_),
    .X(_1620_));
 sky130_fd_sc_hd__mux2i_1 _4826_ (.A0(_1619_),
    .A1(_1620_),
    .S(_1521_),
    .Y(_1621_));
 sky130_fd_sc_hd__a221o_2 _4827_ (.A1(_1196_),
    .A2(_1618_),
    .B1(_1621_),
    .B2(_1310_),
    .C1(_1572_),
    .X(_1622_));
 sky130_fd_sc_hd__a31oi_1 _4828_ (.A1(_1557_),
    .A2(_1612_),
    .A3(_1615_),
    .B1(_1622_),
    .Y(_0057_));
 sky130_fd_sc_hd__mux4_1 _4829_ (.A0(\registers[17][31] ),
    .A1(\registers[19][31] ),
    .A2(\registers[21][31] ),
    .A3(\registers[23][31] ),
    .S0(_1468_),
    .S1(_1524_),
    .X(_1623_));
 sky130_fd_sc_hd__mux2i_2 _4830_ (.A0(\registers[18][31] ),
    .A1(\registers[22][31] ),
    .S(_1489_),
    .Y(_1624_));
 sky130_fd_sc_hd__mux2i_1 _4831_ (.A0(\registers[16][31] ),
    .A1(\registers[20][31] ),
    .S(_1240_),
    .Y(_1625_));
 sky130_fd_sc_hd__a221oi_2 _4832_ (.A1(_1488_),
    .A2(_1624_),
    .B1(_1625_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1626_));
 sky130_fd_sc_hd__o21ai_0 _4833_ (.A1(_1467_),
    .A2(_1623_),
    .B1(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__mux4_1 _4834_ (.A0(\registers[24][31] ),
    .A1(\registers[26][31] ),
    .A2(\registers[28][31] ),
    .A3(\registers[30][31] ),
    .S0(_1546_),
    .S1(_1192_),
    .X(_1628_));
 sky130_fd_sc_hd__mux4_1 _4835_ (.A0(\registers[25][31] ),
    .A1(\registers[27][31] ),
    .A2(\registers[29][31] ),
    .A3(\registers[31][31] ),
    .S0(_1596_),
    .S1(_1205_),
    .X(_1629_));
 sky130_fd_sc_hd__a22oi_2 _4836_ (.A1(_1496_),
    .A2(_1628_),
    .B1(_1629_),
    .B2(_1476_),
    .Y(_1630_));
 sky130_fd_sc_hd__mux4_1 _4837_ (.A0(\registers[8][31] ),
    .A1(\registers[9][31] ),
    .A2(\registers[10][31] ),
    .A3(\registers[11][31] ),
    .S0(_1478_),
    .S1(_1479_),
    .X(_1631_));
 sky130_fd_sc_hd__mux4_1 _4838_ (.A0(\registers[12][31] ),
    .A1(\registers[13][31] ),
    .A2(\registers[14][31] ),
    .A3(\registers[15][31] ),
    .S0(_1301_),
    .S1(_1583_),
    .X(_1632_));
 sky130_fd_sc_hd__mux2i_2 _4839_ (.A0(_1631_),
    .A1(_1632_),
    .S(_1601_),
    .Y(_1633_));
 sky130_fd_sc_hd__mux4_1 _4840_ (.A0(\registers[1][31] ),
    .A1(\registers[3][31] ),
    .A2(\registers[5][31] ),
    .A3(\registers[7][31] ),
    .S0(_1224_),
    .S1(_1225_),
    .X(_1634_));
 sky130_fd_sc_hd__mux4_1 _4841_ (.A0(\registers[0][31] ),
    .A1(\registers[2][31] ),
    .A2(\registers[4][31] ),
    .A3(\registers[6][31] ),
    .S0(_1604_),
    .S1(_1191_),
    .X(_1635_));
 sky130_fd_sc_hd__mux2i_1 _4842_ (.A0(_1634_),
    .A1(_1635_),
    .S(_1521_),
    .Y(_1636_));
 sky130_fd_sc_hd__a221o_2 _4843_ (.A1(_1196_),
    .A2(_1633_),
    .B1(_1636_),
    .B2(_1310_),
    .C1(_1572_),
    .X(_1637_));
 sky130_fd_sc_hd__a31oi_1 _4844_ (.A1(_1557_),
    .A2(_1627_),
    .A3(_1630_),
    .B1(_1637_),
    .Y(_0058_));
 sky130_fd_sc_hd__mux4_1 _4845_ (.A0(\registers[25][3] ),
    .A1(\registers[27][3] ),
    .A2(\registers[29][3] ),
    .A3(\registers[31][3] ),
    .S0(_1166_),
    .S1(_1160_),
    .X(_1638_));
 sky130_fd_sc_hd__mux2i_1 _4846_ (.A0(\registers[24][3] ),
    .A1(\registers[28][3] ),
    .S(_1243_),
    .Y(_1639_));
 sky130_fd_sc_hd__nand2_1 _4847_ (.A(_1169_),
    .B(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__mux2i_1 _4848_ (.A0(\registers[26][3] ),
    .A1(\registers[30][3] ),
    .S(_1163_),
    .Y(_1641_));
 sky130_fd_sc_hd__nand2_1 _4849_ (.A(_1173_),
    .B(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__o2111ai_4 _4850_ (.A1(_1153_),
    .A2(_1638_),
    .B1(_1640_),
    .C1(_1642_),
    .D1(_1176_),
    .Y(_1643_));
 sky130_fd_sc_hd__mux4_1 _4851_ (.A0(\registers[16][3] ),
    .A1(\registers[18][3] ),
    .A2(\registers[20][3] ),
    .A3(\registers[22][3] ),
    .S0(_1546_),
    .S1(_1192_),
    .X(_1644_));
 sky130_fd_sc_hd__mux4_1 _4852_ (.A0(\registers[17][3] ),
    .A1(\registers[19][3] ),
    .A2(\registers[21][3] ),
    .A3(\registers[23][3] ),
    .S0(_1596_),
    .S1(_1205_),
    .X(_1645_));
 sky130_fd_sc_hd__a22oi_1 _4853_ (.A1(_1181_),
    .A2(_1644_),
    .B1(_1645_),
    .B2(_1182_),
    .Y(_1646_));
 sky130_fd_sc_hd__mux4_1 _4854_ (.A0(\registers[0][3] ),
    .A1(\registers[1][3] ),
    .A2(\registers[2][3] ),
    .A3(\registers[3][3] ),
    .S0(_1189_),
    .S1(_1178_),
    .X(_1647_));
 sky130_fd_sc_hd__mux4_1 _4855_ (.A0(\registers[4][3] ),
    .A1(\registers[5][3] ),
    .A2(\registers[6][3] ),
    .A3(\registers[7][3] ),
    .S0(_1301_),
    .S1(_1583_),
    .X(_1648_));
 sky130_fd_sc_hd__mux2i_1 _4856_ (.A0(_1647_),
    .A1(_1648_),
    .S(_1601_),
    .Y(_1649_));
 sky130_fd_sc_hd__mux4_1 _4857_ (.A0(\registers[9][3] ),
    .A1(\registers[11][3] ),
    .A2(\registers[13][3] ),
    .A3(\registers[15][3] ),
    .S0(_1224_),
    .S1(_1225_),
    .X(_1650_));
 sky130_fd_sc_hd__mux4_1 _4858_ (.A0(\registers[8][3] ),
    .A1(\registers[10][3] ),
    .A2(\registers[12][3] ),
    .A3(\registers[14][3] ),
    .S0(_1604_),
    .S1(_1191_),
    .X(_1651_));
 sky130_fd_sc_hd__mux2i_4 _4859_ (.A0(_1650_),
    .A1(_1651_),
    .S(_1521_),
    .Y(_1652_));
 sky130_fd_sc_hd__a221o_2 _4860_ (.A1(_1420_),
    .A2(_1649_),
    .B1(_1652_),
    .B2(_1429_),
    .C1(_1572_),
    .X(_1653_));
 sky130_fd_sc_hd__a31oi_2 _4861_ (.A1(_1557_),
    .A2(_1643_),
    .A3(_1646_),
    .B1(_1653_),
    .Y(_0059_));
 sky130_fd_sc_hd__mux4_1 _4862_ (.A0(\registers[17][4] ),
    .A1(\registers[19][4] ),
    .A2(\registers[21][4] ),
    .A3(\registers[23][4] ),
    .S0(_1468_),
    .S1(_1524_),
    .X(_1654_));
 sky130_fd_sc_hd__mux2i_1 _4863_ (.A0(\registers[18][4] ),
    .A1(\registers[22][4] ),
    .S(_1489_),
    .Y(_1655_));
 sky130_fd_sc_hd__mux2i_1 _4864_ (.A0(\registers[16][4] ),
    .A1(\registers[20][4] ),
    .S(_1240_),
    .Y(_1656_));
 sky130_fd_sc_hd__a221oi_1 _4865_ (.A1(_1488_),
    .A2(_1655_),
    .B1(_1656_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1657_));
 sky130_fd_sc_hd__o21ai_0 _4866_ (.A1(_1467_),
    .A2(_1654_),
    .B1(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hd__mux4_1 _4867_ (.A0(\registers[24][4] ),
    .A1(\registers[26][4] ),
    .A2(\registers[28][4] ),
    .A3(\registers[30][4] ),
    .S0(_1546_),
    .S1(_1192_),
    .X(_1659_));
 sky130_fd_sc_hd__mux4_1 _4868_ (.A0(\registers[25][4] ),
    .A1(\registers[27][4] ),
    .A2(\registers[29][4] ),
    .A3(\registers[31][4] ),
    .S0(_1596_),
    .S1(_1205_),
    .X(_1660_));
 sky130_fd_sc_hd__a22oi_2 _4869_ (.A1(_1496_),
    .A2(_1659_),
    .B1(_1660_),
    .B2(_1476_),
    .Y(_1661_));
 sky130_fd_sc_hd__mux4_1 _4870_ (.A0(\registers[0][4] ),
    .A1(\registers[1][4] ),
    .A2(\registers[2][4] ),
    .A3(\registers[3][4] ),
    .S0(_1189_),
    .S1(_1178_),
    .X(_1662_));
 sky130_fd_sc_hd__mux4_1 _4871_ (.A0(\registers[4][4] ),
    .A1(\registers[5][4] ),
    .A2(\registers[6][4] ),
    .A3(\registers[7][4] ),
    .S0(_1301_),
    .S1(_1583_),
    .X(_1663_));
 sky130_fd_sc_hd__mux2i_1 _4872_ (.A0(_1662_),
    .A1(_1663_),
    .S(_1601_),
    .Y(_1664_));
 sky130_fd_sc_hd__mux4_1 _4873_ (.A0(\registers[9][4] ),
    .A1(\registers[11][4] ),
    .A2(\registers[13][4] ),
    .A3(\registers[15][4] ),
    .S0(_1224_),
    .S1(_1225_),
    .X(_1665_));
 sky130_fd_sc_hd__mux4_1 _4874_ (.A0(\registers[8][4] ),
    .A1(\registers[10][4] ),
    .A2(\registers[12][4] ),
    .A3(\registers[14][4] ),
    .S0(_1604_),
    .S1(_1191_),
    .X(_1666_));
 sky130_fd_sc_hd__mux2i_2 _4875_ (.A0(_1665_),
    .A1(_1666_),
    .S(_1521_),
    .Y(_1667_));
 sky130_fd_sc_hd__a221o_1 _4876_ (.A1(_1420_),
    .A2(_1664_),
    .B1(_1667_),
    .B2(_1429_),
    .C1(_1572_),
    .X(_1668_));
 sky130_fd_sc_hd__a31oi_1 _4877_ (.A1(_1557_),
    .A2(_1658_),
    .A3(_1661_),
    .B1(_1668_),
    .Y(_0060_));
 sky130_fd_sc_hd__mux4_1 _4878_ (.A0(\registers[25][5] ),
    .A1(\registers[27][5] ),
    .A2(\registers[29][5] ),
    .A3(\registers[31][5] ),
    .S0(_1166_),
    .S1(_1160_),
    .X(_1669_));
 sky130_fd_sc_hd__mux2i_1 _4879_ (.A0(\registers[24][5] ),
    .A1(\registers[28][5] ),
    .S(_1243_),
    .Y(_1670_));
 sky130_fd_sc_hd__nand2_1 _4880_ (.A(_1169_),
    .B(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__mux2i_1 _4881_ (.A0(\registers[26][5] ),
    .A1(\registers[30][5] ),
    .S(_1163_),
    .Y(_1672_));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(_1173_),
    .B(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__o2111ai_4 _4883_ (.A1(_1153_),
    .A2(_1669_),
    .B1(_1671_),
    .C1(_1673_),
    .D1(_1176_),
    .Y(_1674_));
 sky130_fd_sc_hd__mux4_1 _4884_ (.A0(\registers[16][5] ),
    .A1(\registers[18][5] ),
    .A2(\registers[20][5] ),
    .A3(\registers[22][5] ),
    .S0(_1546_),
    .S1(_1192_),
    .X(_1675_));
 sky130_fd_sc_hd__mux4_1 _4885_ (.A0(\registers[17][5] ),
    .A1(\registers[19][5] ),
    .A2(\registers[21][5] ),
    .A3(\registers[23][5] ),
    .S0(_1596_),
    .S1(_1205_),
    .X(_1676_));
 sky130_fd_sc_hd__a22oi_1 _4886_ (.A1(_1181_),
    .A2(_1675_),
    .B1(_1676_),
    .B2(_1182_),
    .Y(_1677_));
 sky130_fd_sc_hd__mux4_1 _4887_ (.A0(\registers[0][5] ),
    .A1(\registers[1][5] ),
    .A2(\registers[2][5] ),
    .A3(\registers[3][5] ),
    .S0(_1189_),
    .S1(_1178_),
    .X(_1678_));
 sky130_fd_sc_hd__mux4_1 _4888_ (.A0(\registers[4][5] ),
    .A1(\registers[5][5] ),
    .A2(\registers[6][5] ),
    .A3(\registers[7][5] ),
    .S0(_1301_),
    .S1(_1583_),
    .X(_1679_));
 sky130_fd_sc_hd__mux2i_1 _4889_ (.A0(_1678_),
    .A1(_1679_),
    .S(_1601_),
    .Y(_1680_));
 sky130_fd_sc_hd__mux4_1 _4890_ (.A0(\registers[9][5] ),
    .A1(\registers[11][5] ),
    .A2(\registers[13][5] ),
    .A3(\registers[15][5] ),
    .S0(_1224_),
    .S1(_1225_),
    .X(_1681_));
 sky130_fd_sc_hd__mux4_1 _4891_ (.A0(\registers[8][5] ),
    .A1(\registers[10][5] ),
    .A2(\registers[12][5] ),
    .A3(\registers[14][5] ),
    .S0(_1604_),
    .S1(_1191_),
    .X(_1682_));
 sky130_fd_sc_hd__mux2i_2 _4892_ (.A0(_1681_),
    .A1(_1682_),
    .S(_1152_),
    .Y(_1683_));
 sky130_fd_sc_hd__a221o_2 _4893_ (.A1(_1420_),
    .A2(_1680_),
    .B1(_1683_),
    .B2(_1429_),
    .C1(_1572_),
    .X(_1684_));
 sky130_fd_sc_hd__a31oi_2 _4894_ (.A1(_1557_),
    .A2(_1674_),
    .A3(_1677_),
    .B1(_1684_),
    .Y(_0061_));
 sky130_fd_sc_hd__mux4_1 _4895_ (.A0(\registers[17][6] ),
    .A1(\registers[19][6] ),
    .A2(\registers[21][6] ),
    .A3(\registers[23][6] ),
    .S0(_1468_),
    .S1(_1524_),
    .X(_1685_));
 sky130_fd_sc_hd__mux2i_1 _4896_ (.A0(\registers[18][6] ),
    .A1(\registers[22][6] ),
    .S(_1489_),
    .Y(_1686_));
 sky130_fd_sc_hd__mux2i_1 _4897_ (.A0(\registers[16][6] ),
    .A1(\registers[20][6] ),
    .S(_1240_),
    .Y(_1687_));
 sky130_fd_sc_hd__a221oi_1 _4898_ (.A1(_1488_),
    .A2(_1686_),
    .B1(_1687_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1688_));
 sky130_fd_sc_hd__o21ai_0 _4899_ (.A1(_1467_),
    .A2(_1685_),
    .B1(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hd__mux4_1 _4900_ (.A0(\registers[24][6] ),
    .A1(\registers[26][6] ),
    .A2(\registers[28][6] ),
    .A3(\registers[30][6] ),
    .S0(_1546_),
    .S1(_1192_),
    .X(_1690_));
 sky130_fd_sc_hd__mux4_1 _4901_ (.A0(\registers[25][6] ),
    .A1(\registers[27][6] ),
    .A2(\registers[29][6] ),
    .A3(\registers[31][6] ),
    .S0(_1596_),
    .S1(_1205_),
    .X(_1691_));
 sky130_fd_sc_hd__a22oi_2 _4902_ (.A1(_1496_),
    .A2(_1690_),
    .B1(_1691_),
    .B2(_1476_),
    .Y(_1692_));
 sky130_fd_sc_hd__mux4_1 _4903_ (.A0(\registers[0][6] ),
    .A1(\registers[1][6] ),
    .A2(\registers[2][6] ),
    .A3(\registers[3][6] ),
    .S0(_1189_),
    .S1(_1178_),
    .X(_1693_));
 sky130_fd_sc_hd__mux4_1 _4904_ (.A0(\registers[4][6] ),
    .A1(\registers[5][6] ),
    .A2(\registers[6][6] ),
    .A3(\registers[7][6] ),
    .S0(_1301_),
    .S1(_1583_),
    .X(_1694_));
 sky130_fd_sc_hd__mux2i_1 _4905_ (.A0(_1693_),
    .A1(_1694_),
    .S(_1601_),
    .Y(_1695_));
 sky130_fd_sc_hd__mux4_1 _4906_ (.A0(\registers[9][6] ),
    .A1(\registers[11][6] ),
    .A2(\registers[13][6] ),
    .A3(\registers[15][6] ),
    .S0(_1224_),
    .S1(_1225_),
    .X(_1696_));
 sky130_fd_sc_hd__mux4_1 _4907_ (.A0(\registers[8][6] ),
    .A1(\registers[10][6] ),
    .A2(\registers[12][6] ),
    .A3(\registers[14][6] ),
    .S0(_1604_),
    .S1(_1191_),
    .X(_1697_));
 sky130_fd_sc_hd__mux2i_1 _4908_ (.A0(_1696_),
    .A1(_1697_),
    .S(_1152_),
    .Y(_1698_));
 sky130_fd_sc_hd__a221o_1 _4909_ (.A1(_1310_),
    .A2(_1695_),
    .B1(_1698_),
    .B2(_1195_),
    .C1(_1572_),
    .X(_1699_));
 sky130_fd_sc_hd__a31oi_1 _4910_ (.A1(_1557_),
    .A2(_1689_),
    .A3(_1692_),
    .B1(_1699_),
    .Y(_0062_));
 sky130_fd_sc_hd__mux4_1 _4911_ (.A0(\registers[17][7] ),
    .A1(\registers[19][7] ),
    .A2(\registers[21][7] ),
    .A3(\registers[23][7] ),
    .S0(_1183_),
    .S1(_1524_),
    .X(_1700_));
 sky130_fd_sc_hd__mux2i_1 _4912_ (.A0(\registers[18][7] ),
    .A1(\registers[22][7] ),
    .S(_1489_),
    .Y(_1701_));
 sky130_fd_sc_hd__mux2i_1 _4913_ (.A0(\registers[16][7] ),
    .A1(\registers[20][7] ),
    .S(_1240_),
    .Y(_1702_));
 sky130_fd_sc_hd__a221oi_2 _4914_ (.A1(_1488_),
    .A2(_1701_),
    .B1(_1702_),
    .B2(_1492_),
    .C1(_1493_),
    .Y(_1703_));
 sky130_fd_sc_hd__o21ai_1 _4915_ (.A1(_1154_),
    .A2(_1700_),
    .B1(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__mux4_1 _4916_ (.A0(\registers[24][7] ),
    .A1(\registers[26][7] ),
    .A2(\registers[28][7] ),
    .A3(\registers[30][7] ),
    .S0(_1157_),
    .S1(_1192_),
    .X(_1705_));
 sky130_fd_sc_hd__mux4_1 _4917_ (.A0(\registers[25][7] ),
    .A1(\registers[27][7] ),
    .A2(\registers[29][7] ),
    .A3(\registers[31][7] ),
    .S0(_1596_),
    .S1(_1205_),
    .X(_1706_));
 sky130_fd_sc_hd__a22oi_4 _4918_ (.A1(_1496_),
    .A2(_1705_),
    .B1(_1706_),
    .B2(_1214_),
    .Y(_1707_));
 sky130_fd_sc_hd__mux4_1 _4919_ (.A0(\registers[8][7] ),
    .A1(\registers[9][7] ),
    .A2(\registers[10][7] ),
    .A3(\registers[11][7] ),
    .S0(_1189_),
    .S1(_1178_),
    .X(_1708_));
 sky130_fd_sc_hd__mux4_1 _4920_ (.A0(\registers[12][7] ),
    .A1(\registers[13][7] ),
    .A2(\registers[14][7] ),
    .A3(\registers[15][7] ),
    .S0(_1301_),
    .S1(_1583_),
    .X(_1709_));
 sky130_fd_sc_hd__mux2i_1 _4921_ (.A0(_1708_),
    .A1(_1709_),
    .S(_1601_),
    .Y(_1710_));
 sky130_fd_sc_hd__mux4_1 _4922_ (.A0(\registers[1][7] ),
    .A1(\registers[3][7] ),
    .A2(\registers[5][7] ),
    .A3(\registers[7][7] ),
    .S0(_1224_),
    .S1(_1225_),
    .X(_1711_));
 sky130_fd_sc_hd__mux4_1 _4923_ (.A0(\registers[0][7] ),
    .A1(\registers[2][7] ),
    .A2(\registers[4][7] ),
    .A3(\registers[6][7] ),
    .S0(_1604_),
    .S1(_1191_),
    .X(_1712_));
 sky130_fd_sc_hd__mux2i_1 _4924_ (.A0(_1711_),
    .A1(_1712_),
    .S(_1152_),
    .Y(_1713_));
 sky130_fd_sc_hd__a221o_2 _4925_ (.A1(_1196_),
    .A2(_1710_),
    .B1(_1713_),
    .B2(_1186_),
    .C1(_1572_),
    .X(_1714_));
 sky130_fd_sc_hd__a31oi_4 _4926_ (.A1(_1557_),
    .A2(_1704_),
    .A3(_1707_),
    .B1(_1714_),
    .Y(_0063_));
 sky130_fd_sc_hd__mux4_1 _4927_ (.A0(\registers[17][8] ),
    .A1(\registers[19][8] ),
    .A2(\registers[21][8] ),
    .A3(\registers[23][8] ),
    .S0(_1183_),
    .S1(_1524_),
    .X(_1715_));
 sky130_fd_sc_hd__mux2i_1 _4928_ (.A0(\registers[18][8] ),
    .A1(\registers[22][8] ),
    .S(_1162_),
    .Y(_1716_));
 sky130_fd_sc_hd__mux2i_1 _4929_ (.A0(\registers[16][8] ),
    .A1(\registers[20][8] ),
    .S(_1240_),
    .Y(_1717_));
 sky130_fd_sc_hd__a221oi_1 _4930_ (.A1(_1172_),
    .A2(_1716_),
    .B1(_1717_),
    .B2(_1168_),
    .C1(_1175_),
    .Y(_1718_));
 sky130_fd_sc_hd__o21ai_1 _4931_ (.A1(_1154_),
    .A2(_1715_),
    .B1(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__mux4_1 _4932_ (.A0(\registers[24][8] ),
    .A1(\registers[26][8] ),
    .A2(\registers[28][8] ),
    .A3(\registers[30][8] ),
    .S0(_1157_),
    .S1(_1192_),
    .X(_1720_));
 sky130_fd_sc_hd__mux4_1 _4933_ (.A0(\registers[25][8] ),
    .A1(\registers[27][8] ),
    .A2(\registers[29][8] ),
    .A3(\registers[31][8] ),
    .S0(_1596_),
    .S1(_1205_),
    .X(_1721_));
 sky130_fd_sc_hd__a22oi_4 _4934_ (.A1(_1212_),
    .A2(_1720_),
    .B1(_1721_),
    .B2(_1214_),
    .Y(_1722_));
 sky130_fd_sc_hd__mux4_1 _4935_ (.A0(\registers[0][8] ),
    .A1(\registers[1][8] ),
    .A2(\registers[2][8] ),
    .A3(\registers[3][8] ),
    .S0(_1189_),
    .S1(_1178_),
    .X(_1723_));
 sky130_fd_sc_hd__mux4_1 _4936_ (.A0(\registers[4][8] ),
    .A1(\registers[5][8] ),
    .A2(\registers[6][8] ),
    .A3(\registers[7][8] ),
    .S0(_1301_),
    .S1(_1583_),
    .X(_1724_));
 sky130_fd_sc_hd__mux2i_1 _4937_ (.A0(_1723_),
    .A1(_1724_),
    .S(_1601_),
    .Y(_1725_));
 sky130_fd_sc_hd__mux4_1 _4938_ (.A0(\registers[9][8] ),
    .A1(\registers[11][8] ),
    .A2(\registers[13][8] ),
    .A3(\registers[15][8] ),
    .S0(_1224_),
    .S1(_1225_),
    .X(_1726_));
 sky130_fd_sc_hd__mux4_1 _4939_ (.A0(\registers[8][8] ),
    .A1(\registers[10][8] ),
    .A2(\registers[12][8] ),
    .A3(\registers[14][8] ),
    .S0(_1604_),
    .S1(_1191_),
    .X(_1727_));
 sky130_fd_sc_hd__mux2i_1 _4940_ (.A0(_1726_),
    .A1(_1727_),
    .S(_1152_),
    .Y(_1728_));
 sky130_fd_sc_hd__a221o_2 _4941_ (.A1(_1310_),
    .A2(_1725_),
    .B1(_1728_),
    .B2(_1195_),
    .C1(_1200_),
    .X(_1729_));
 sky130_fd_sc_hd__a31oi_4 _4942_ (.A1(_1148_),
    .A2(_1719_),
    .A3(_1722_),
    .B1(_1729_),
    .Y(_0064_));
 sky130_fd_sc_hd__mux4_1 _4943_ (.A0(\registers[17][9] ),
    .A1(\registers[19][9] ),
    .A2(\registers[21][9] ),
    .A3(\registers[23][9] ),
    .S0(_1183_),
    .S1(_1179_),
    .X(_1730_));
 sky130_fd_sc_hd__mux2i_1 _4944_ (.A0(\registers[18][9] ),
    .A1(\registers[22][9] ),
    .S(_1162_),
    .Y(_1731_));
 sky130_fd_sc_hd__mux2i_1 _4945_ (.A0(\registers[16][9] ),
    .A1(\registers[20][9] ),
    .S(_1240_),
    .Y(_1732_));
 sky130_fd_sc_hd__a221oi_1 _4946_ (.A1(_1172_),
    .A2(_1731_),
    .B1(_1732_),
    .B2(_1168_),
    .C1(_1175_),
    .Y(_1733_));
 sky130_fd_sc_hd__o21ai_1 _4947_ (.A1(_1154_),
    .A2(_1730_),
    .B1(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__mux4_1 _4948_ (.A0(\registers[24][9] ),
    .A1(\registers[26][9] ),
    .A2(\registers[28][9] ),
    .A3(\registers[30][9] ),
    .S0(_1157_),
    .S1(_1192_),
    .X(_1735_));
 sky130_fd_sc_hd__mux4_1 _4949_ (.A0(\registers[25][9] ),
    .A1(\registers[27][9] ),
    .A2(\registers[29][9] ),
    .A3(\registers[31][9] ),
    .S0(_1596_),
    .S1(_1205_),
    .X(_1736_));
 sky130_fd_sc_hd__a22oi_2 _4950_ (.A1(_1212_),
    .A2(_1735_),
    .B1(_1736_),
    .B2(_1214_),
    .Y(_1737_));
 sky130_fd_sc_hd__mux4_1 _4951_ (.A0(\registers[8][9] ),
    .A1(\registers[9][9] ),
    .A2(\registers[10][9] ),
    .A3(\registers[11][9] ),
    .S0(_1189_),
    .S1(_1178_),
    .X(_1738_));
 sky130_fd_sc_hd__mux4_1 _4952_ (.A0(\registers[12][9] ),
    .A1(\registers[13][9] ),
    .A2(\registers[14][9] ),
    .A3(\registers[15][9] ),
    .S0(_1301_),
    .S1(_1167_),
    .X(_1739_));
 sky130_fd_sc_hd__mux2i_1 _4953_ (.A0(_1738_),
    .A1(_1739_),
    .S(_1601_),
    .Y(_1740_));
 sky130_fd_sc_hd__mux4_1 _4954_ (.A0(\registers[1][9] ),
    .A1(\registers[3][9] ),
    .A2(\registers[5][9] ),
    .A3(\registers[7][9] ),
    .S0(_1224_),
    .S1(_1225_),
    .X(_1741_));
 sky130_fd_sc_hd__mux4_1 _4955_ (.A0(\registers[0][9] ),
    .A1(\registers[2][9] ),
    .A2(\registers[4][9] ),
    .A3(\registers[6][9] ),
    .S0(_1604_),
    .S1(_1191_),
    .X(_1742_));
 sky130_fd_sc_hd__mux2i_1 _4956_ (.A0(_1741_),
    .A1(_1742_),
    .S(_1152_),
    .Y(_1743_));
 sky130_fd_sc_hd__a221o_2 _4957_ (.A1(_1228_),
    .A2(_1740_),
    .B1(_1743_),
    .B2(_1186_),
    .C1(_1200_),
    .X(_1744_));
 sky130_fd_sc_hd__a31oi_4 _4958_ (.A1(_1148_),
    .A2(_1734_),
    .A3(_1737_),
    .B1(_1744_),
    .Y(_0065_));
 sky130_fd_sc_hd__buf_8 _4959_ (.A(net167),
    .X(_1745_));
 sky130_fd_sc_hd__buf_4 _4960_ (.A(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__buf_6 _4961_ (.A(read_addr2[0]),
    .X(_1747_));
 sky130_fd_sc_hd__clkinvlp_4 _4962_ (.A(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__buf_16 _4963_ (.A(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__buf_12 _4964_ (.A(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__buf_16 _4965_ (.A(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__buf_8 _4966_ (.A(read_addr2[1]),
    .X(_1752_));
 sky130_fd_sc_hd__buf_16 _4967_ (.A(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__buf_8 _4968_ (.A(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__clkbuf_2 _4969_ (.A(read_addr2[2]),
    .X(_1755_));
 sky130_fd_sc_hd__buf_6 _4970_ (.A(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__buf_8 _4971_ (.A(_1756_),
    .X(_1757_));
 sky130_fd_sc_hd__mux4_1 _4972_ (.A0(\registers[25][0] ),
    .A1(\registers[27][0] ),
    .A2(\registers[29][0] ),
    .A3(\registers[31][0] ),
    .S0(_1754_),
    .S1(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__buf_6 _4973_ (.A(_1756_),
    .X(_1759_));
 sky130_fd_sc_hd__buf_6 _4974_ (.A(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__mux2i_1 _4975_ (.A0(\registers[24][0] ),
    .A1(\registers[28][0] ),
    .S(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__buf_6 _4976_ (.A(_1747_),
    .X(_1762_));
 sky130_fd_sc_hd__buf_8 _4977_ (.A(_1752_),
    .X(_1763_));
 sky130_fd_sc_hd__buf_6 _4978_ (.A(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__nor2_2 _4979_ (.A(_1762_),
    .B(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__buf_6 _4980_ (.A(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__nand2_1 _4981_ (.A(_1761_),
    .B(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__mux2i_1 _4982_ (.A0(\registers[26][0] ),
    .A1(\registers[30][0] ),
    .S(_1760_),
    .Y(_1768_));
 sky130_fd_sc_hd__nor2b_2 _4983_ (.A(_1762_),
    .B_N(_1764_),
    .Y(_1769_));
 sky130_fd_sc_hd__buf_6 _4984_ (.A(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__nand2_1 _4985_ (.A(_1768_),
    .B(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__buf_8 _4986_ (.A(net2),
    .X(_1772_));
 sky130_fd_sc_hd__buf_16 _4987_ (.A(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__o2111ai_4 _4988_ (.A1(_1751_),
    .A2(_1758_),
    .B1(_1767_),
    .C1(_1771_),
    .D1(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__buf_6 _4989_ (.A(_1753_),
    .X(_1775_));
 sky130_fd_sc_hd__buf_6 _4990_ (.A(_1759_),
    .X(_1776_));
 sky130_fd_sc_hd__mux4_1 _4991_ (.A0(\registers[16][0] ),
    .A1(\registers[18][0] ),
    .A2(\registers[20][0] ),
    .A3(\registers[22][0] ),
    .S0(_1775_),
    .S1(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__nor2_8 _4992_ (.A(_1762_),
    .B(_1772_),
    .Y(_1778_));
 sky130_fd_sc_hd__nor2_8 _4993_ (.A(_1750_),
    .B(_1772_),
    .Y(_1779_));
 sky130_fd_sc_hd__buf_8 _4994_ (.A(_1753_),
    .X(_1780_));
 sky130_fd_sc_hd__mux4_1 _4995_ (.A0(\registers[17][0] ),
    .A1(\registers[19][0] ),
    .A2(\registers[21][0] ),
    .A3(\registers[23][0] ),
    .S0(_1780_),
    .S1(_1776_),
    .X(_1781_));
 sky130_fd_sc_hd__a22oi_1 _4996_ (.A1(_1777_),
    .A2(_1778_),
    .B1(_1779_),
    .B2(_1781_),
    .Y(_1782_));
 sky130_fd_sc_hd__nor2b_1 _4997_ (.A(_1745_),
    .B_N(net2),
    .Y(_1783_));
 sky130_fd_sc_hd__buf_2 _4998_ (.A(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__buf_8 _4999_ (.A(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__mux4_1 _5000_ (.A0(\registers[8][0] ),
    .A1(\registers[9][0] ),
    .A2(\registers[10][0] ),
    .A3(\registers[11][0] ),
    .S0(_1762_),
    .S1(_1780_),
    .X(_1786_));
 sky130_fd_sc_hd__buf_6 _5001_ (.A(_1747_),
    .X(_1787_));
 sky130_fd_sc_hd__mux4_1 _5002_ (.A0(\registers[12][0] ),
    .A1(\registers[13][0] ),
    .A2(\registers[14][0] ),
    .A3(\registers[15][0] ),
    .S0(_1787_),
    .S1(_1775_),
    .X(_1788_));
 sky130_fd_sc_hd__buf_8 _5003_ (.A(_1755_),
    .X(_1789_));
 sky130_fd_sc_hd__buf_8 _5004_ (.A(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__mux2i_1 _5005_ (.A0(_1786_),
    .A1(_1788_),
    .S(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__nor2_4 _5006_ (.A(_1772_),
    .B(_1745_),
    .Y(_1792_));
 sky130_fd_sc_hd__buf_4 _5007_ (.A(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__mux4_1 _5008_ (.A0(\registers[1][0] ),
    .A1(\registers[3][0] ),
    .A2(\registers[5][0] ),
    .A3(\registers[7][0] ),
    .S0(_1752_),
    .S1(_1756_),
    .X(_1794_));
 sky130_fd_sc_hd__mux4_1 _5009_ (.A0(\registers[0][0] ),
    .A1(\registers[2][0] ),
    .A2(\registers[4][0] ),
    .A3(\registers[6][0] ),
    .S0(_1752_),
    .S1(_1756_),
    .X(_1795_));
 sky130_fd_sc_hd__mux2i_1 _5010_ (.A0(_1794_),
    .A1(_1795_),
    .S(_1749_),
    .Y(_1796_));
 sky130_fd_sc_hd__nand2_4 _5011_ (.A(_1122_),
    .B(net4),
    .Y(_1797_));
 sky130_fd_sc_hd__buf_4 _5012_ (.A(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__a221o_2 _5013_ (.A1(_1785_),
    .A2(_1791_),
    .B1(_1793_),
    .B2(_1796_),
    .C1(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__a31oi_2 _5014_ (.A1(_1746_),
    .A2(_1774_),
    .A3(_1782_),
    .B1(_1799_),
    .Y(_0066_));
 sky130_fd_sc_hd__clkbuf_4 _5015_ (.A(_1749_),
    .X(_1800_));
 sky130_fd_sc_hd__buf_4 _5016_ (.A(_1763_),
    .X(_1801_));
 sky130_fd_sc_hd__buf_6 _5017_ (.A(_1759_),
    .X(_1802_));
 sky130_fd_sc_hd__mux4_1 _5018_ (.A0(\registers[17][10] ),
    .A1(\registers[19][10] ),
    .A2(\registers[21][10] ),
    .A3(\registers[23][10] ),
    .S0(_1801_),
    .S1(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__mux2i_1 _5019_ (.A0(\registers[18][10] ),
    .A1(\registers[22][10] ),
    .S(_1757_),
    .Y(_1804_));
 sky130_fd_sc_hd__mux2i_1 _5020_ (.A0(\registers[16][10] ),
    .A1(\registers[20][10] ),
    .S(_1776_),
    .Y(_1805_));
 sky130_fd_sc_hd__a221oi_1 _5021_ (.A1(_1770_),
    .A2(_1804_),
    .B1(_1805_),
    .B2(_1766_),
    .C1(_1773_),
    .Y(_1806_));
 sky130_fd_sc_hd__o21ai_1 _5022_ (.A1(_1800_),
    .A2(_1803_),
    .B1(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__mux4_1 _5023_ (.A0(\registers[24][10] ),
    .A1(\registers[26][10] ),
    .A2(\registers[28][10] ),
    .A3(\registers[30][10] ),
    .S0(_1775_),
    .S1(_1776_),
    .X(_1808_));
 sky130_fd_sc_hd__nor2b_4 _5024_ (.A(_1762_),
    .B_N(_1772_),
    .Y(_1809_));
 sky130_fd_sc_hd__and2_0 _5025_ (.A(_1762_),
    .B(_1772_),
    .X(_1810_));
 sky130_fd_sc_hd__buf_4 _5026_ (.A(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__buf_8 _5027_ (.A(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__mux4_1 _5028_ (.A0(\registers[25][10] ),
    .A1(\registers[27][10] ),
    .A2(\registers[29][10] ),
    .A3(\registers[31][10] ),
    .S0(_1780_),
    .S1(_1776_),
    .X(_1813_));
 sky130_fd_sc_hd__a22oi_2 _5029_ (.A1(_1808_),
    .A2(_1809_),
    .B1(_1812_),
    .B2(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__mux4_1 _5030_ (.A0(\registers[0][10] ),
    .A1(\registers[1][10] ),
    .A2(\registers[2][10] ),
    .A3(\registers[3][10] ),
    .S0(_1762_),
    .S1(_1780_),
    .X(_1815_));
 sky130_fd_sc_hd__buf_6 _5031_ (.A(_1753_),
    .X(_1816_));
 sky130_fd_sc_hd__mux4_1 _5032_ (.A0(\registers[4][10] ),
    .A1(\registers[5][10] ),
    .A2(\registers[6][10] ),
    .A3(\registers[7][10] ),
    .S0(_1787_),
    .S1(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__mux2i_1 _5033_ (.A0(_1815_),
    .A1(_1817_),
    .S(_1790_),
    .Y(_1818_));
 sky130_fd_sc_hd__buf_8 _5034_ (.A(_1756_),
    .X(_1819_));
 sky130_fd_sc_hd__mux4_1 _5035_ (.A0(\registers[9][10] ),
    .A1(\registers[11][10] ),
    .A2(\registers[13][10] ),
    .A3(\registers[15][10] ),
    .S0(_1753_),
    .S1(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__buf_8 _5036_ (.A(_1752_),
    .X(_1821_));
 sky130_fd_sc_hd__buf_8 _5037_ (.A(_1756_),
    .X(_1822_));
 sky130_fd_sc_hd__mux4_1 _5038_ (.A0(\registers[8][10] ),
    .A1(\registers[10][10] ),
    .A2(\registers[12][10] ),
    .A3(\registers[14][10] ),
    .S0(_1821_),
    .S1(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__mux2i_1 _5039_ (.A0(_1820_),
    .A1(_1823_),
    .S(_1750_),
    .Y(_1824_));
 sky130_fd_sc_hd__clkbuf_8 _5040_ (.A(_1784_),
    .X(_1825_));
 sky130_fd_sc_hd__a221o_2 _5041_ (.A1(_1793_),
    .A2(_1818_),
    .B1(_1824_),
    .B2(_1825_),
    .C1(_1798_),
    .X(_1826_));
 sky130_fd_sc_hd__a31oi_4 _5042_ (.A1(_1746_),
    .A2(_1807_),
    .A3(_1814_),
    .B1(_1826_),
    .Y(_0067_));
 sky130_fd_sc_hd__mux4_1 _5043_ (.A0(\registers[17][11] ),
    .A1(\registers[19][11] ),
    .A2(\registers[21][11] ),
    .A3(\registers[23][11] ),
    .S0(_1801_),
    .S1(_1802_),
    .X(_1827_));
 sky130_fd_sc_hd__buf_4 _5044_ (.A(_1769_),
    .X(_1828_));
 sky130_fd_sc_hd__buf_6 _5045_ (.A(_1756_),
    .X(_1829_));
 sky130_fd_sc_hd__mux2i_1 _5046_ (.A0(\registers[18][11] ),
    .A1(\registers[22][11] ),
    .S(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__mux2i_1 _5047_ (.A0(\registers[16][11] ),
    .A1(\registers[20][11] ),
    .S(_1776_),
    .Y(_1831_));
 sky130_fd_sc_hd__buf_6 _5048_ (.A(_1765_),
    .X(_1832_));
 sky130_fd_sc_hd__buf_4 _5049_ (.A(_1772_),
    .X(_1833_));
 sky130_fd_sc_hd__a221oi_2 _5050_ (.A1(_1828_),
    .A2(_1830_),
    .B1(_1831_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__o21ai_0 _5051_ (.A1(_1800_),
    .A2(_1827_),
    .B1(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__buf_8 _5052_ (.A(_1809_),
    .X(_1836_));
 sky130_fd_sc_hd__buf_6 _5053_ (.A(_1819_),
    .X(_1837_));
 sky130_fd_sc_hd__mux4_1 _5054_ (.A0(\registers[24][11] ),
    .A1(\registers[26][11] ),
    .A2(\registers[28][11] ),
    .A3(\registers[30][11] ),
    .S0(_1764_),
    .S1(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__buf_6 _5055_ (.A(_1763_),
    .X(_1839_));
 sky130_fd_sc_hd__buf_8 _5056_ (.A(_1759_),
    .X(_1840_));
 sky130_fd_sc_hd__mux4_1 _5057_ (.A0(\registers[25][11] ),
    .A1(\registers[27][11] ),
    .A2(\registers[29][11] ),
    .A3(\registers[31][11] ),
    .S0(_1839_),
    .S1(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__a22oi_2 _5058_ (.A1(_1836_),
    .A2(_1838_),
    .B1(_1841_),
    .B2(_1812_),
    .Y(_1842_));
 sky130_fd_sc_hd__mux4_1 _5059_ (.A0(\registers[0][11] ),
    .A1(\registers[1][11] ),
    .A2(\registers[2][11] ),
    .A3(\registers[3][11] ),
    .S0(_1762_),
    .S1(_1780_),
    .X(_1843_));
 sky130_fd_sc_hd__mux4_1 _5060_ (.A0(\registers[4][11] ),
    .A1(\registers[5][11] ),
    .A2(\registers[6][11] ),
    .A3(\registers[7][11] ),
    .S0(_1787_),
    .S1(_1816_),
    .X(_1844_));
 sky130_fd_sc_hd__buf_8 _5061_ (.A(_1819_),
    .X(_1845_));
 sky130_fd_sc_hd__mux2i_1 _5062_ (.A0(_1843_),
    .A1(_1844_),
    .S(_1845_),
    .Y(_1846_));
 sky130_fd_sc_hd__mux4_1 _5063_ (.A0(\registers[9][11] ),
    .A1(\registers[11][11] ),
    .A2(\registers[13][11] ),
    .A3(\registers[15][11] ),
    .S0(_1753_),
    .S1(_1819_),
    .X(_1847_));
 sky130_fd_sc_hd__buf_6 _5064_ (.A(_1752_),
    .X(_1848_));
 sky130_fd_sc_hd__mux4_1 _5065_ (.A0(\registers[8][11] ),
    .A1(\registers[10][11] ),
    .A2(\registers[12][11] ),
    .A3(\registers[14][11] ),
    .S0(_1848_),
    .S1(_1822_),
    .X(_1849_));
 sky130_fd_sc_hd__mux2i_1 _5066_ (.A0(_1847_),
    .A1(_1849_),
    .S(_1750_),
    .Y(_1850_));
 sky130_fd_sc_hd__a221o_1 _5067_ (.A1(_1793_),
    .A2(_1846_),
    .B1(_1850_),
    .B2(_1825_),
    .C1(_1798_),
    .X(_1851_));
 sky130_fd_sc_hd__a31oi_2 _5068_ (.A1(_1746_),
    .A2(_1835_),
    .A3(_1842_),
    .B1(_1851_),
    .Y(_0068_));
 sky130_fd_sc_hd__mux4_1 _5069_ (.A0(\registers[25][12] ),
    .A1(\registers[27][12] ),
    .A2(\registers[29][12] ),
    .A3(\registers[31][12] ),
    .S0(_1754_),
    .S1(_1757_),
    .X(_1852_));
 sky130_fd_sc_hd__mux2i_1 _5070_ (.A0(\registers[24][12] ),
    .A1(\registers[28][12] ),
    .S(_1840_),
    .Y(_1853_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(_1766_),
    .B(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__mux2i_1 _5072_ (.A0(\registers[26][12] ),
    .A1(\registers[30][12] ),
    .S(_1760_),
    .Y(_1855_));
 sky130_fd_sc_hd__nand2_1 _5073_ (.A(_1770_),
    .B(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__o2111ai_4 _5074_ (.A1(_1751_),
    .A2(_1852_),
    .B1(_1854_),
    .C1(_1856_),
    .D1(_1773_),
    .Y(_1857_));
 sky130_fd_sc_hd__mux4_1 _5075_ (.A0(\registers[16][12] ),
    .A1(\registers[18][12] ),
    .A2(\registers[20][12] ),
    .A3(\registers[22][12] ),
    .S0(_1764_),
    .S1(_1837_),
    .X(_1858_));
 sky130_fd_sc_hd__mux4_1 _5076_ (.A0(\registers[17][12] ),
    .A1(\registers[19][12] ),
    .A2(\registers[21][12] ),
    .A3(\registers[23][12] ),
    .S0(_1839_),
    .S1(_1840_),
    .X(_1859_));
 sky130_fd_sc_hd__a22oi_1 _5077_ (.A1(_1778_),
    .A2(_1858_),
    .B1(_1859_),
    .B2(_1779_),
    .Y(_1860_));
 sky130_fd_sc_hd__mux4_1 _5078_ (.A0(\registers[0][12] ),
    .A1(\registers[1][12] ),
    .A2(\registers[2][12] ),
    .A3(\registers[3][12] ),
    .S0(_1762_),
    .S1(_1780_),
    .X(_1861_));
 sky130_fd_sc_hd__buf_6 _5079_ (.A(_1747_),
    .X(_1862_));
 sky130_fd_sc_hd__mux4_1 _5080_ (.A0(\registers[4][12] ),
    .A1(\registers[5][12] ),
    .A2(\registers[6][12] ),
    .A3(\registers[7][12] ),
    .S0(_1862_),
    .S1(_1816_),
    .X(_1863_));
 sky130_fd_sc_hd__mux2i_1 _5081_ (.A0(_1861_),
    .A1(_1863_),
    .S(_1845_),
    .Y(_1864_));
 sky130_fd_sc_hd__buf_6 _5082_ (.A(_1752_),
    .X(_1865_));
 sky130_fd_sc_hd__mux4_1 _5083_ (.A0(\registers[9][12] ),
    .A1(\registers[11][12] ),
    .A2(\registers[13][12] ),
    .A3(\registers[15][12] ),
    .S0(_1865_),
    .S1(_1819_),
    .X(_1866_));
 sky130_fd_sc_hd__buf_6 _5084_ (.A(_1755_),
    .X(_1867_));
 sky130_fd_sc_hd__mux4_1 _5085_ (.A0(\registers[8][12] ),
    .A1(\registers[10][12] ),
    .A2(\registers[12][12] ),
    .A3(\registers[14][12] ),
    .S0(_1848_),
    .S1(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__mux2i_4 _5086_ (.A0(_1866_),
    .A1(_1868_),
    .S(_1750_),
    .Y(_1869_));
 sky130_fd_sc_hd__a221o_2 _5087_ (.A1(_1793_),
    .A2(_1864_),
    .B1(_1869_),
    .B2(_1825_),
    .C1(_1798_),
    .X(_1870_));
 sky130_fd_sc_hd__a31oi_2 _5088_ (.A1(_1746_),
    .A2(_1857_),
    .A3(_1860_),
    .B1(_1870_),
    .Y(_0069_));
 sky130_fd_sc_hd__buf_4 _5089_ (.A(_1759_),
    .X(_1871_));
 sky130_fd_sc_hd__mux4_1 _5090_ (.A0(\registers[17][13] ),
    .A1(\registers[19][13] ),
    .A2(\registers[21][13] ),
    .A3(\registers[23][13] ),
    .S0(_1801_),
    .S1(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__mux2i_1 _5091_ (.A0(\registers[18][13] ),
    .A1(\registers[22][13] ),
    .S(_1829_),
    .Y(_1873_));
 sky130_fd_sc_hd__mux2i_1 _5092_ (.A0(\registers[16][13] ),
    .A1(\registers[20][13] ),
    .S(_1776_),
    .Y(_1874_));
 sky130_fd_sc_hd__a221oi_1 _5093_ (.A1(_1828_),
    .A2(_1873_),
    .B1(_1874_),
    .B2(_1832_),
    .C1(_1833_),
    .Y(_1875_));
 sky130_fd_sc_hd__o21ai_0 _5094_ (.A1(_1800_),
    .A2(_1872_),
    .B1(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__buf_6 _5095_ (.A(_1819_),
    .X(_1877_));
 sky130_fd_sc_hd__mux4_1 _5096_ (.A0(\registers[24][13] ),
    .A1(\registers[26][13] ),
    .A2(\registers[28][13] ),
    .A3(\registers[30][13] ),
    .S0(_1764_),
    .S1(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__buf_6 _5097_ (.A(_1759_),
    .X(_1879_));
 sky130_fd_sc_hd__mux4_1 _5098_ (.A0(\registers[25][13] ),
    .A1(\registers[27][13] ),
    .A2(\registers[29][13] ),
    .A3(\registers[31][13] ),
    .S0(_1839_),
    .S1(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__a22oi_2 _5099_ (.A1(_1836_),
    .A2(_1878_),
    .B1(_1880_),
    .B2(_1812_),
    .Y(_1881_));
 sky130_fd_sc_hd__mux4_1 _5100_ (.A0(\registers[0][13] ),
    .A1(\registers[1][13] ),
    .A2(\registers[2][13] ),
    .A3(\registers[3][13] ),
    .S0(_1762_),
    .S1(_1780_),
    .X(_1882_));
 sky130_fd_sc_hd__mux4_1 _5101_ (.A0(\registers[4][13] ),
    .A1(\registers[5][13] ),
    .A2(\registers[6][13] ),
    .A3(\registers[7][13] ),
    .S0(_1862_),
    .S1(_1816_),
    .X(_1883_));
 sky130_fd_sc_hd__mux2i_1 _5102_ (.A0(_1882_),
    .A1(_1883_),
    .S(_1845_),
    .Y(_1884_));
 sky130_fd_sc_hd__buf_4 _5103_ (.A(_1756_),
    .X(_1885_));
 sky130_fd_sc_hd__mux4_1 _5104_ (.A0(\registers[9][13] ),
    .A1(\registers[11][13] ),
    .A2(\registers[13][13] ),
    .A3(\registers[15][13] ),
    .S0(_1865_),
    .S1(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__mux4_1 _5105_ (.A0(\registers[8][13] ),
    .A1(\registers[10][13] ),
    .A2(\registers[12][13] ),
    .A3(\registers[14][13] ),
    .S0(_1848_),
    .S1(_1867_),
    .X(_1887_));
 sky130_fd_sc_hd__mux2i_4 _5106_ (.A0(_1886_),
    .A1(_1887_),
    .S(_1750_),
    .Y(_1888_));
 sky130_fd_sc_hd__a221o_1 _5107_ (.A1(_1793_),
    .A2(_1884_),
    .B1(_1888_),
    .B2(_1825_),
    .C1(_1798_),
    .X(_1889_));
 sky130_fd_sc_hd__a31oi_1 _5108_ (.A1(_1746_),
    .A2(_1876_),
    .A3(_1881_),
    .B1(_1889_),
    .Y(_0070_));
 sky130_fd_sc_hd__mux4_1 _5109_ (.A0(\registers[25][14] ),
    .A1(\registers[27][14] ),
    .A2(\registers[29][14] ),
    .A3(\registers[31][14] ),
    .S0(_1754_),
    .S1(_1757_),
    .X(_1890_));
 sky130_fd_sc_hd__mux2i_1 _5110_ (.A0(\registers[24][14] ),
    .A1(\registers[28][14] ),
    .S(_1840_),
    .Y(_1891_));
 sky130_fd_sc_hd__nand2_1 _5111_ (.A(_1766_),
    .B(_1891_),
    .Y(_1892_));
 sky130_fd_sc_hd__mux2i_1 _5112_ (.A0(\registers[26][14] ),
    .A1(\registers[30][14] ),
    .S(_1760_),
    .Y(_1893_));
 sky130_fd_sc_hd__nand2_1 _5113_ (.A(_1770_),
    .B(_1893_),
    .Y(_1894_));
 sky130_fd_sc_hd__o2111ai_4 _5114_ (.A1(_1751_),
    .A2(_1890_),
    .B1(_1892_),
    .C1(_1894_),
    .D1(_1773_),
    .Y(_1895_));
 sky130_fd_sc_hd__mux4_1 _5115_ (.A0(\registers[16][14] ),
    .A1(\registers[18][14] ),
    .A2(\registers[20][14] ),
    .A3(\registers[22][14] ),
    .S0(_1764_),
    .S1(_1877_),
    .X(_1896_));
 sky130_fd_sc_hd__mux4_1 _5116_ (.A0(\registers[17][14] ),
    .A1(\registers[19][14] ),
    .A2(\registers[21][14] ),
    .A3(\registers[23][14] ),
    .S0(_1839_),
    .S1(_1879_),
    .X(_1897_));
 sky130_fd_sc_hd__a22oi_1 _5117_ (.A1(_1778_),
    .A2(_1896_),
    .B1(_1897_),
    .B2(_1779_),
    .Y(_1898_));
 sky130_fd_sc_hd__buf_16 _5118_ (.A(_1747_),
    .X(_1899_));
 sky130_fd_sc_hd__buf_16 _5119_ (.A(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__buf_6 _5120_ (.A(_1763_),
    .X(_1901_));
 sky130_fd_sc_hd__mux4_1 _5121_ (.A0(\registers[0][14] ),
    .A1(\registers[1][14] ),
    .A2(\registers[2][14] ),
    .A3(\registers[3][14] ),
    .S0(_1900_),
    .S1(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__mux4_1 _5122_ (.A0(\registers[4][14] ),
    .A1(\registers[5][14] ),
    .A2(\registers[6][14] ),
    .A3(\registers[7][14] ),
    .S0(_1862_),
    .S1(_1816_),
    .X(_1903_));
 sky130_fd_sc_hd__mux2i_1 _5123_ (.A0(_1902_),
    .A1(_1903_),
    .S(_1845_),
    .Y(_1904_));
 sky130_fd_sc_hd__mux4_1 _5124_ (.A0(\registers[9][14] ),
    .A1(\registers[11][14] ),
    .A2(\registers[13][14] ),
    .A3(\registers[15][14] ),
    .S0(_1865_),
    .S1(_1885_),
    .X(_1905_));
 sky130_fd_sc_hd__mux4_1 _5125_ (.A0(\registers[8][14] ),
    .A1(\registers[10][14] ),
    .A2(\registers[12][14] ),
    .A3(\registers[14][14] ),
    .S0(_1848_),
    .S1(_1867_),
    .X(_1906_));
 sky130_fd_sc_hd__mux2i_1 _5126_ (.A0(_1905_),
    .A1(_1906_),
    .S(_1750_),
    .Y(_1907_));
 sky130_fd_sc_hd__a221o_2 _5127_ (.A1(_1793_),
    .A2(_1904_),
    .B1(_1907_),
    .B2(_1825_),
    .C1(_1798_),
    .X(_1908_));
 sky130_fd_sc_hd__a31oi_2 _5128_ (.A1(_1746_),
    .A2(_1895_),
    .A3(_1898_),
    .B1(_1908_),
    .Y(_0071_));
 sky130_fd_sc_hd__mux4_1 _5129_ (.A0(\registers[17][15] ),
    .A1(\registers[19][15] ),
    .A2(\registers[21][15] ),
    .A3(\registers[23][15] ),
    .S0(_1801_),
    .S1(_1871_),
    .X(_1909_));
 sky130_fd_sc_hd__mux2i_1 _5130_ (.A0(\registers[18][15] ),
    .A1(\registers[22][15] ),
    .S(_1829_),
    .Y(_1910_));
 sky130_fd_sc_hd__mux2i_1 _5131_ (.A0(\registers[16][15] ),
    .A1(\registers[20][15] ),
    .S(_1776_),
    .Y(_1911_));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[0]$_SDFFCE_PN0P_  (.D(_0034_),
    .DE(_0032_),
    .Q(net44),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[10]$_SDFFCE_PN0P_  (.D(_0035_),
    .DE(_0032_),
    .Q(net45),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[11]$_SDFFCE_PN0P_  (.D(_0036_),
    .DE(_0032_),
    .Q(net46),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[12]$_SDFFCE_PN0P_  (.D(_0037_),
    .DE(_0032_),
    .Q(net47),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[13]$_SDFFCE_PN0P_  (.D(_0038_),
    .DE(_0032_),
    .Q(net48),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[14]$_SDFFCE_PN0P_  (.D(_0039_),
    .DE(_0032_),
    .Q(net49),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[15]$_SDFFCE_PN0P_  (.D(_0040_),
    .DE(_0032_),
    .Q(net50),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[16]$_SDFFCE_PN0P_  (.D(_0041_),
    .DE(_0032_),
    .Q(net51),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[17]$_SDFFCE_PN0P_  (.D(_0042_),
    .DE(_0032_),
    .Q(net52),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[18]$_SDFFCE_PN0P_  (.D(_0043_),
    .DE(_0032_),
    .Q(net53),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[19]$_SDFFCE_PN0P_  (.D(_0044_),
    .DE(_0032_),
    .Q(net54),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[1]$_SDFFCE_PN0P_  (.D(_0045_),
    .DE(_0032_),
    .Q(net55),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[20]$_SDFFCE_PN0P_  (.D(_0046_),
    .DE(_0032_),
    .Q(net56),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[21]$_SDFFCE_PN0P_  (.D(_0047_),
    .DE(_0032_),
    .Q(net57),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[22]$_SDFFCE_PN0P_  (.D(_0048_),
    .DE(_0032_),
    .Q(net58),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[23]$_SDFFCE_PN0P_  (.D(_0049_),
    .DE(_0032_),
    .Q(net59),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[24]$_SDFFCE_PN0P_  (.D(_0050_),
    .DE(_0032_),
    .Q(net60),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[25]$_SDFFCE_PN0P_  (.D(_0051_),
    .DE(_0032_),
    .Q(net61),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[26]$_SDFFCE_PN0P_  (.D(_0052_),
    .DE(_0032_),
    .Q(net62),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[27]$_SDFFCE_PN0P_  (.D(_0053_),
    .DE(_0032_),
    .Q(net63),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[28]$_SDFFCE_PN0P_  (.D(_0054_),
    .DE(_0032_),
    .Q(net64),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[29]$_SDFFCE_PN0P_  (.D(_0055_),
    .DE(_0032_),
    .Q(net65),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[2]$_SDFFCE_PN0P_  (.D(_0056_),
    .DE(_0032_),
    .Q(net66),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[30]$_SDFFCE_PN0P_  (.D(_0057_),
    .DE(_0032_),
    .Q(net67),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[31]$_SDFFCE_PN0P_  (.D(_0058_),
    .DE(_0032_),
    .Q(net68),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[3]$_SDFFCE_PN0P_  (.D(_0059_),
    .DE(_0032_),
    .Q(net69),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[4]$_SDFFCE_PN0P_  (.D(_0060_),
    .DE(_0032_),
    .Q(net70),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[5]$_SDFFCE_PN0P_  (.D(_0061_),
    .DE(_0032_),
    .Q(net71),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[6]$_SDFFCE_PN0P_  (.D(_0062_),
    .DE(_0032_),
    .Q(net72),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[7]$_SDFFCE_PN0P_  (.D(_0063_),
    .DE(_0032_),
    .Q(net73),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[8]$_SDFFCE_PN0P_  (.D(_0064_),
    .DE(_0032_),
    .Q(net74),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data1[9]$_SDFFCE_PN0P_  (.D(_0065_),
    .DE(_0032_),
    .Q(net75),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[0]$_SDFFCE_PN0P_  (.D(_0066_),
    .DE(_0033_),
    .Q(net76),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[10]$_SDFFCE_PN0P_  (.D(_0067_),
    .DE(_0033_),
    .Q(net77),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[11]$_SDFFCE_PN0P_  (.D(_0068_),
    .DE(_0033_),
    .Q(net78),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[12]$_SDFFCE_PN0P_  (.D(_0069_),
    .DE(_0033_),
    .Q(net79),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[13]$_SDFFCE_PN0P_  (.D(_0070_),
    .DE(_0033_),
    .Q(net80),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[14]$_SDFFCE_PN0P_  (.D(_0071_),
    .DE(_0033_),
    .Q(net81),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[15]$_SDFFCE_PN0P_  (.D(_0072_),
    .DE(_0033_),
    .Q(net82),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[16]$_SDFFCE_PN0P_  (.D(_0073_),
    .DE(_0033_),
    .Q(net83),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[17]$_SDFFCE_PN0P_  (.D(_0074_),
    .DE(_0033_),
    .Q(net84),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[18]$_SDFFCE_PN0P_  (.D(_0075_),
    .DE(_0033_),
    .Q(net85),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[19]$_SDFFCE_PN0P_  (.D(_0076_),
    .DE(_0033_),
    .Q(net86),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[1]$_SDFFCE_PN0P_  (.D(_0077_),
    .DE(_0033_),
    .Q(net87),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[20]$_SDFFCE_PN0P_  (.D(_0078_),
    .DE(_0033_),
    .Q(net88),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[21]$_SDFFCE_PN0P_  (.D(_0079_),
    .DE(_0033_),
    .Q(net89),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[22]$_SDFFCE_PN0P_  (.D(_0080_),
    .DE(_0033_),
    .Q(net90),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[23]$_SDFFCE_PN0P_  (.D(_0081_),
    .DE(_0033_),
    .Q(net91),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[24]$_SDFFCE_PN0P_  (.D(_0082_),
    .DE(_0033_),
    .Q(net92),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[25]$_SDFFCE_PN0P_  (.D(_0083_),
    .DE(_0033_),
    .Q(net93),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[26]$_SDFFCE_PN0P_  (.D(_0084_),
    .DE(_0033_),
    .Q(net94),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[27]$_SDFFCE_PN0P_  (.D(_0085_),
    .DE(_0033_),
    .Q(net95),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[28]$_SDFFCE_PN0P_  (.D(_0086_),
    .DE(_0033_),
    .Q(net96),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[29]$_SDFFCE_PN0P_  (.D(_0087_),
    .DE(_0033_),
    .Q(net97),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[2]$_SDFFCE_PN0P_  (.D(_0088_),
    .DE(_0033_),
    .Q(net98),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[30]$_SDFFCE_PN0P_  (.D(_0089_),
    .DE(_0033_),
    .Q(net99),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[31]$_SDFFCE_PN0P_  (.D(_0090_),
    .DE(_0033_),
    .Q(net100),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[3]$_SDFFCE_PN0P_  (.D(_0091_),
    .DE(_0033_),
    .Q(net101),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[4]$_SDFFCE_PN0P_  (.D(_0092_),
    .DE(_0033_),
    .Q(net102),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[5]$_SDFFCE_PN0P_  (.D(_0093_),
    .DE(_0033_),
    .Q(net103),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[6]$_SDFFCE_PN0P_  (.D(_0094_),
    .DE(_0033_),
    .Q(net104),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[7]$_SDFFCE_PN0P_  (.D(_0095_),
    .DE(_0033_),
    .Q(net105),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[8]$_SDFFCE_PN0P_  (.D(_0096_),
    .DE(_0033_),
    .Q(net106),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \read_data2[9]$_SDFFCE_PN0P_  (.D(_0097_),
    .DE(_0033_),
    .Q(net107),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][0]$_SDFFCE_PN0P_  (.D(_0098_),
    .DE(_0031_),
    .Q(\registers[0][0] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][10]$_SDFFCE_PN0P_  (.D(_0099_),
    .DE(_0031_),
    .Q(\registers[0][10] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][11]$_SDFFCE_PN0P_  (.D(_0100_),
    .DE(_0031_),
    .Q(\registers[0][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][12]$_SDFFCE_PN0P_  (.D(_0101_),
    .DE(_0031_),
    .Q(\registers[0][12] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][13]$_SDFFCE_PN0P_  (.D(_0102_),
    .DE(_0031_),
    .Q(\registers[0][13] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][14]$_SDFFCE_PN0P_  (.D(_0103_),
    .DE(_0031_),
    .Q(\registers[0][14] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][15]$_SDFFCE_PN0P_  (.D(_0104_),
    .DE(_0031_),
    .Q(\registers[0][15] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][16]$_SDFFCE_PN0P_  (.D(_0105_),
    .DE(_0031_),
    .Q(\registers[0][16] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][17]$_SDFFCE_PN0P_  (.D(_0106_),
    .DE(_0031_),
    .Q(\registers[0][17] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][18]$_SDFFCE_PN0P_  (.D(_0107_),
    .DE(_0031_),
    .Q(\registers[0][18] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][19]$_SDFFCE_PN0P_  (.D(_0108_),
    .DE(net113),
    .Q(\registers[0][19] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][1]$_SDFFCE_PN0P_  (.D(_0109_),
    .DE(net113),
    .Q(\registers[0][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][20]$_SDFFCE_PN0P_  (.D(_0110_),
    .DE(net113),
    .Q(\registers[0][20] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][21]$_SDFFCE_PN0P_  (.D(_0111_),
    .DE(net113),
    .Q(\registers[0][21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][22]$_SDFFCE_PN0P_  (.D(_0112_),
    .DE(net113),
    .Q(\registers[0][22] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][23]$_SDFFCE_PN0P_  (.D(_0113_),
    .DE(net113),
    .Q(\registers[0][23] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][24]$_SDFFCE_PN0P_  (.D(_0114_),
    .DE(net113),
    .Q(\registers[0][24] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][25]$_SDFFCE_PN0P_  (.D(_0115_),
    .DE(net113),
    .Q(\registers[0][25] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][26]$_SDFFCE_PN0P_  (.D(_0116_),
    .DE(net113),
    .Q(\registers[0][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][27]$_SDFFCE_PN0P_  (.D(_0117_),
    .DE(net113),
    .Q(\registers[0][27] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][28]$_SDFFCE_PN0P_  (.D(_0118_),
    .DE(_0031_),
    .Q(\registers[0][28] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][29]$_SDFFCE_PN0P_  (.D(_0119_),
    .DE(net113),
    .Q(\registers[0][29] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][2]$_SDFFCE_PN0P_  (.D(_0120_),
    .DE(net113),
    .Q(\registers[0][2] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][30]$_SDFFCE_PN0P_  (.D(_0121_),
    .DE(net113),
    .Q(\registers[0][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][31]$_SDFFCE_PN0P_  (.D(_0122_),
    .DE(net113),
    .Q(\registers[0][31] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][3]$_SDFFCE_PN0P_  (.D(_0123_),
    .DE(_0031_),
    .Q(\registers[0][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][4]$_SDFFCE_PN0P_  (.D(_0124_),
    .DE(_0031_),
    .Q(\registers[0][4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][5]$_SDFFCE_PN0P_  (.D(_0125_),
    .DE(_0031_),
    .Q(\registers[0][5] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][6]$_SDFFCE_PN0P_  (.D(_0126_),
    .DE(_0031_),
    .Q(\registers[0][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][7]$_SDFFCE_PN0P_  (.D(_0127_),
    .DE(_0031_),
    .Q(\registers[0][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][8]$_SDFFCE_PN0P_  (.D(_0128_),
    .DE(_0031_),
    .Q(\registers[0][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[0][9]$_SDFFCE_PN0P_  (.D(_0129_),
    .DE(_0031_),
    .Q(\registers[0][9] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][0]$_SDFFCE_PN0P_  (.D(_0130_),
    .DE(net134),
    .Q(\registers[10][0] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][10]$_SDFFCE_PN0P_  (.D(_0131_),
    .DE(net134),
    .Q(\registers[10][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][11]$_SDFFCE_PN0P_  (.D(_0132_),
    .DE(net134),
    .Q(\registers[10][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][12]$_SDFFCE_PN0P_  (.D(_0133_),
    .DE(net134),
    .Q(\registers[10][12] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][13]$_SDFFCE_PN0P_  (.D(_0134_),
    .DE(net134),
    .Q(\registers[10][13] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][14]$_SDFFCE_PN0P_  (.D(_0135_),
    .DE(net134),
    .Q(\registers[10][14] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][15]$_SDFFCE_PN0P_  (.D(_0136_),
    .DE(net134),
    .Q(\registers[10][15] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][16]$_SDFFCE_PN0P_  (.D(_0137_),
    .DE(net134),
    .Q(\registers[10][16] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][17]$_SDFFCE_PN0P_  (.D(_0138_),
    .DE(net134),
    .Q(\registers[10][17] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][18]$_SDFFCE_PN0P_  (.D(_0139_),
    .DE(net134),
    .Q(\registers[10][18] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][19]$_SDFFCE_PN0P_  (.D(_0140_),
    .DE(net134),
    .Q(\registers[10][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][1]$_SDFFCE_PN0P_  (.D(_0141_),
    .DE(net134),
    .Q(\registers[10][1] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][20]$_SDFFCE_PN0P_  (.D(_0142_),
    .DE(net134),
    .Q(\registers[10][20] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][21]$_SDFFCE_PN0P_  (.D(_0143_),
    .DE(net134),
    .Q(\registers[10][21] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][22]$_SDFFCE_PN0P_  (.D(_0144_),
    .DE(net134),
    .Q(\registers[10][22] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][23]$_SDFFCE_PN0P_  (.D(_0145_),
    .DE(net134),
    .Q(\registers[10][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][24]$_SDFFCE_PN0P_  (.D(_0146_),
    .DE(net134),
    .Q(\registers[10][24] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][25]$_SDFFCE_PN0P_  (.D(_0147_),
    .DE(net134),
    .Q(\registers[10][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][26]$_SDFFCE_PN0P_  (.D(_0148_),
    .DE(_0030_),
    .Q(\registers[10][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][27]$_SDFFCE_PN0P_  (.D(_0149_),
    .DE(net134),
    .Q(\registers[10][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][28]$_SDFFCE_PN0P_  (.D(_0150_),
    .DE(_0030_),
    .Q(\registers[10][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][29]$_SDFFCE_PN0P_  (.D(_0151_),
    .DE(_0030_),
    .Q(\registers[10][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][2]$_SDFFCE_PN0P_  (.D(_0152_),
    .DE(_0030_),
    .Q(\registers[10][2] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][30]$_SDFFCE_PN0P_  (.D(_0153_),
    .DE(_0030_),
    .Q(\registers[10][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][31]$_SDFFCE_PN0P_  (.D(_0154_),
    .DE(_0030_),
    .Q(\registers[10][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][3]$_SDFFCE_PN0P_  (.D(_0155_),
    .DE(_0030_),
    .Q(\registers[10][3] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][4]$_SDFFCE_PN0P_  (.D(_0156_),
    .DE(_0030_),
    .Q(\registers[10][4] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][5]$_SDFFCE_PN0P_  (.D(_0157_),
    .DE(_0030_),
    .Q(\registers[10][5] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][6]$_SDFFCE_PN0P_  (.D(_0158_),
    .DE(_0030_),
    .Q(\registers[10][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][7]$_SDFFCE_PN0P_  (.D(_0159_),
    .DE(_0030_),
    .Q(\registers[10][7] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][8]$_SDFFCE_PN0P_  (.D(_0160_),
    .DE(_0030_),
    .Q(\registers[10][8] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[10][9]$_SDFFCE_PN0P_  (.D(_0161_),
    .DE(_0030_),
    .Q(\registers[10][9] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][0]$_SDFFCE_PN0P_  (.D(_0162_),
    .DE(net121),
    .Q(\registers[11][0] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][10]$_SDFFCE_PN0P_  (.D(_0163_),
    .DE(net121),
    .Q(\registers[11][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][11]$_SDFFCE_PN0P_  (.D(_0164_),
    .DE(net121),
    .Q(\registers[11][11] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][12]$_SDFFCE_PN0P_  (.D(_0165_),
    .DE(net121),
    .Q(\registers[11][12] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][13]$_SDFFCE_PN0P_  (.D(_0166_),
    .DE(net121),
    .Q(\registers[11][13] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][14]$_SDFFCE_PN0P_  (.D(_0167_),
    .DE(net121),
    .Q(\registers[11][14] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][15]$_SDFFCE_PN0P_  (.D(_0168_),
    .DE(net121),
    .Q(\registers[11][15] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][16]$_SDFFCE_PN0P_  (.D(_0169_),
    .DE(net121),
    .Q(\registers[11][16] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][17]$_SDFFCE_PN0P_  (.D(_0170_),
    .DE(net121),
    .Q(\registers[11][17] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][18]$_SDFFCE_PN0P_  (.D(_0171_),
    .DE(net121),
    .Q(\registers[11][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][19]$_SDFFCE_PN0P_  (.D(_0172_),
    .DE(net121),
    .Q(\registers[11][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][1]$_SDFFCE_PN0P_  (.D(_0173_),
    .DE(net121),
    .Q(\registers[11][1] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][20]$_SDFFCE_PN0P_  (.D(_0174_),
    .DE(net121),
    .Q(\registers[11][20] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][21]$_SDFFCE_PN0P_  (.D(_0175_),
    .DE(net121),
    .Q(\registers[11][21] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][22]$_SDFFCE_PN0P_  (.D(_0176_),
    .DE(net121),
    .Q(\registers[11][22] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][23]$_SDFFCE_PN0P_  (.D(_0177_),
    .DE(net121),
    .Q(\registers[11][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][24]$_SDFFCE_PN0P_  (.D(_0178_),
    .DE(net121),
    .Q(\registers[11][24] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][25]$_SDFFCE_PN0P_  (.D(_0179_),
    .DE(net121),
    .Q(\registers[11][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][26]$_SDFFCE_PN0P_  (.D(_0180_),
    .DE(net121),
    .Q(\registers[11][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][27]$_SDFFCE_PN0P_  (.D(_0181_),
    .DE(net121),
    .Q(\registers[11][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][28]$_SDFFCE_PN0P_  (.D(_0182_),
    .DE(_0029_),
    .Q(\registers[11][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][29]$_SDFFCE_PN0P_  (.D(_0183_),
    .DE(net121),
    .Q(\registers[11][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][2]$_SDFFCE_PN0P_  (.D(_0184_),
    .DE(_0029_),
    .Q(\registers[11][2] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][30]$_SDFFCE_PN0P_  (.D(_0185_),
    .DE(_0029_),
    .Q(\registers[11][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][31]$_SDFFCE_PN0P_  (.D(_0186_),
    .DE(_0029_),
    .Q(\registers[11][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][3]$_SDFFCE_PN0P_  (.D(_0187_),
    .DE(_0029_),
    .Q(\registers[11][3] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][4]$_SDFFCE_PN0P_  (.D(_0188_),
    .DE(_0029_),
    .Q(\registers[11][4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][5]$_SDFFCE_PN0P_  (.D(_0189_),
    .DE(_0029_),
    .Q(\registers[11][5] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][6]$_SDFFCE_PN0P_  (.D(_0190_),
    .DE(_0029_),
    .Q(\registers[11][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][7]$_SDFFCE_PN0P_  (.D(_0191_),
    .DE(_0029_),
    .Q(\registers[11][7] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][8]$_SDFFCE_PN0P_  (.D(_0192_),
    .DE(_0029_),
    .Q(\registers[11][8] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[11][9]$_SDFFCE_PN0P_  (.D(_0193_),
    .DE(_0029_),
    .Q(\registers[11][9] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][0]$_SDFFCE_PN0P_  (.D(_0194_),
    .DE(net112),
    .Q(\registers[12][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][10]$_SDFFCE_PN0P_  (.D(_0195_),
    .DE(net112),
    .Q(\registers[12][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][11]$_SDFFCE_PN0P_  (.D(_0196_),
    .DE(net112),
    .Q(\registers[12][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][12]$_SDFFCE_PN0P_  (.D(_0197_),
    .DE(net112),
    .Q(\registers[12][12] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][13]$_SDFFCE_PN0P_  (.D(_0198_),
    .DE(net112),
    .Q(\registers[12][13] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][14]$_SDFFCE_PN0P_  (.D(_0199_),
    .DE(net112),
    .Q(\registers[12][14] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][15]$_SDFFCE_PN0P_  (.D(_0200_),
    .DE(net112),
    .Q(\registers[12][15] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][16]$_SDFFCE_PN0P_  (.D(_0201_),
    .DE(net112),
    .Q(\registers[12][16] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][17]$_SDFFCE_PN0P_  (.D(_0202_),
    .DE(net112),
    .Q(\registers[12][17] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][18]$_SDFFCE_PN0P_  (.D(_0203_),
    .DE(net112),
    .Q(\registers[12][18] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][19]$_SDFFCE_PN0P_  (.D(_0204_),
    .DE(net112),
    .Q(\registers[12][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][1]$_SDFFCE_PN0P_  (.D(_0205_),
    .DE(net112),
    .Q(\registers[12][1] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][20]$_SDFFCE_PN0P_  (.D(_0206_),
    .DE(net112),
    .Q(\registers[12][20] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][21]$_SDFFCE_PN0P_  (.D(_0207_),
    .DE(net112),
    .Q(\registers[12][21] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][22]$_SDFFCE_PN0P_  (.D(_0208_),
    .DE(net112),
    .Q(\registers[12][22] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][23]$_SDFFCE_PN0P_  (.D(_0209_),
    .DE(net112),
    .Q(\registers[12][23] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][24]$_SDFFCE_PN0P_  (.D(_0210_),
    .DE(net112),
    .Q(\registers[12][24] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][25]$_SDFFCE_PN0P_  (.D(_0211_),
    .DE(net112),
    .Q(\registers[12][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][26]$_SDFFCE_PN0P_  (.D(_0212_),
    .DE(net112),
    .Q(\registers[12][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][27]$_SDFFCE_PN0P_  (.D(_0213_),
    .DE(net112),
    .Q(\registers[12][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][28]$_SDFFCE_PN0P_  (.D(_0214_),
    .DE(_0028_),
    .Q(\registers[12][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][29]$_SDFFCE_PN0P_  (.D(_0215_),
    .DE(_0028_),
    .Q(\registers[12][29] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][2]$_SDFFCE_PN0P_  (.D(_0216_),
    .DE(_0028_),
    .Q(\registers[12][2] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][30]$_SDFFCE_PN0P_  (.D(_0217_),
    .DE(_0028_),
    .Q(\registers[12][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][31]$_SDFFCE_PN0P_  (.D(_0218_),
    .DE(_0028_),
    .Q(\registers[12][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][3]$_SDFFCE_PN0P_  (.D(_0219_),
    .DE(_0028_),
    .Q(\registers[12][3] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][4]$_SDFFCE_PN0P_  (.D(_0220_),
    .DE(_0028_),
    .Q(\registers[12][4] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][5]$_SDFFCE_PN0P_  (.D(_0221_),
    .DE(_0028_),
    .Q(\registers[12][5] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][6]$_SDFFCE_PN0P_  (.D(_0222_),
    .DE(_0028_),
    .Q(\registers[12][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][7]$_SDFFCE_PN0P_  (.D(_0223_),
    .DE(_0028_),
    .Q(\registers[12][7] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][8]$_SDFFCE_PN0P_  (.D(_0224_),
    .DE(_0028_),
    .Q(\registers[12][8] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[12][9]$_SDFFCE_PN0P_  (.D(_0225_),
    .DE(_0028_),
    .Q(\registers[12][9] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][0]$_SDFFCE_PN0P_  (.D(_0226_),
    .DE(net133),
    .Q(\registers[13][0] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][10]$_SDFFCE_PN0P_  (.D(_0227_),
    .DE(net133),
    .Q(\registers[13][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][11]$_SDFFCE_PN0P_  (.D(_0228_),
    .DE(net133),
    .Q(\registers[13][11] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][12]$_SDFFCE_PN0P_  (.D(_0229_),
    .DE(net133),
    .Q(\registers[13][12] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][13]$_SDFFCE_PN0P_  (.D(_0230_),
    .DE(net133),
    .Q(\registers[13][13] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][14]$_SDFFCE_PN0P_  (.D(_0231_),
    .DE(net133),
    .Q(\registers[13][14] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][15]$_SDFFCE_PN0P_  (.D(_0232_),
    .DE(net133),
    .Q(\registers[13][15] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][16]$_SDFFCE_PN0P_  (.D(_0233_),
    .DE(net133),
    .Q(\registers[13][16] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][17]$_SDFFCE_PN0P_  (.D(_0234_),
    .DE(net133),
    .Q(\registers[13][17] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][18]$_SDFFCE_PN0P_  (.D(_0235_),
    .DE(net133),
    .Q(\registers[13][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][19]$_SDFFCE_PN0P_  (.D(_0236_),
    .DE(net133),
    .Q(\registers[13][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][1]$_SDFFCE_PN0P_  (.D(_0237_),
    .DE(net133),
    .Q(\registers[13][1] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][20]$_SDFFCE_PN0P_  (.D(_0238_),
    .DE(net133),
    .Q(\registers[13][20] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][21]$_SDFFCE_PN0P_  (.D(_0239_),
    .DE(net133),
    .Q(\registers[13][21] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][22]$_SDFFCE_PN0P_  (.D(_0240_),
    .DE(net133),
    .Q(\registers[13][22] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][23]$_SDFFCE_PN0P_  (.D(_0241_),
    .DE(net133),
    .Q(\registers[13][23] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][24]$_SDFFCE_PN0P_  (.D(_0242_),
    .DE(net133),
    .Q(\registers[13][24] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][25]$_SDFFCE_PN0P_  (.D(_0243_),
    .DE(net133),
    .Q(\registers[13][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][26]$_SDFFCE_PN0P_  (.D(_0244_),
    .DE(net133),
    .Q(\registers[13][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][27]$_SDFFCE_PN0P_  (.D(_0245_),
    .DE(net133),
    .Q(\registers[13][27] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][28]$_SDFFCE_PN0P_  (.D(_0246_),
    .DE(_0027_),
    .Q(\registers[13][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][29]$_SDFFCE_PN0P_  (.D(_0247_),
    .DE(_0027_),
    .Q(\registers[13][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][2]$_SDFFCE_PN0P_  (.D(_0248_),
    .DE(_0027_),
    .Q(\registers[13][2] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][30]$_SDFFCE_PN0P_  (.D(_0249_),
    .DE(_0027_),
    .Q(\registers[13][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][31]$_SDFFCE_PN0P_  (.D(_0250_),
    .DE(_0027_),
    .Q(\registers[13][31] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][3]$_SDFFCE_PN0P_  (.D(_0251_),
    .DE(_0027_),
    .Q(\registers[13][3] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][4]$_SDFFCE_PN0P_  (.D(_0252_),
    .DE(_0027_),
    .Q(\registers[13][4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][5]$_SDFFCE_PN0P_  (.D(_0253_),
    .DE(_0027_),
    .Q(\registers[13][5] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][6]$_SDFFCE_PN0P_  (.D(_0254_),
    .DE(_0027_),
    .Q(\registers[13][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][7]$_SDFFCE_PN0P_  (.D(_0255_),
    .DE(_0027_),
    .Q(\registers[13][7] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][8]$_SDFFCE_PN0P_  (.D(_0256_),
    .DE(_0027_),
    .Q(\registers[13][8] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[13][9]$_SDFFCE_PN0P_  (.D(_0257_),
    .DE(_0027_),
    .Q(\registers[13][9] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][0]$_SDFFCE_PN0P_  (.D(_0258_),
    .DE(net132),
    .Q(\registers[14][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][10]$_SDFFCE_PN0P_  (.D(_0259_),
    .DE(net132),
    .Q(\registers[14][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][11]$_SDFFCE_PN0P_  (.D(_0260_),
    .DE(net132),
    .Q(\registers[14][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][12]$_SDFFCE_PN0P_  (.D(_0261_),
    .DE(net132),
    .Q(\registers[14][12] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][13]$_SDFFCE_PN0P_  (.D(_0262_),
    .DE(net132),
    .Q(\registers[14][13] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][14]$_SDFFCE_PN0P_  (.D(_0263_),
    .DE(net132),
    .Q(\registers[14][14] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][15]$_SDFFCE_PN0P_  (.D(_0264_),
    .DE(net132),
    .Q(\registers[14][15] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][16]$_SDFFCE_PN0P_  (.D(_0265_),
    .DE(net132),
    .Q(\registers[14][16] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][17]$_SDFFCE_PN0P_  (.D(_0266_),
    .DE(net132),
    .Q(\registers[14][17] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][18]$_SDFFCE_PN0P_  (.D(_0267_),
    .DE(net132),
    .Q(\registers[14][18] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][19]$_SDFFCE_PN0P_  (.D(_0268_),
    .DE(net132),
    .Q(\registers[14][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][1]$_SDFFCE_PN0P_  (.D(_0269_),
    .DE(net132),
    .Q(\registers[14][1] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][20]$_SDFFCE_PN0P_  (.D(_0270_),
    .DE(net132),
    .Q(\registers[14][20] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][21]$_SDFFCE_PN0P_  (.D(_0271_),
    .DE(net132),
    .Q(\registers[14][21] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][22]$_SDFFCE_PN0P_  (.D(_0272_),
    .DE(net132),
    .Q(\registers[14][22] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][23]$_SDFFCE_PN0P_  (.D(_0273_),
    .DE(net132),
    .Q(\registers[14][23] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][24]$_SDFFCE_PN0P_  (.D(_0274_),
    .DE(net132),
    .Q(\registers[14][24] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][25]$_SDFFCE_PN0P_  (.D(_0275_),
    .DE(net132),
    .Q(\registers[14][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][26]$_SDFFCE_PN0P_  (.D(_0276_),
    .DE(net132),
    .Q(\registers[14][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][27]$_SDFFCE_PN0P_  (.D(_0277_),
    .DE(net132),
    .Q(\registers[14][27] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][28]$_SDFFCE_PN0P_  (.D(_0278_),
    .DE(_0026_),
    .Q(\registers[14][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][29]$_SDFFCE_PN0P_  (.D(_0279_),
    .DE(net132),
    .Q(\registers[14][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][2]$_SDFFCE_PN0P_  (.D(_0280_),
    .DE(_0026_),
    .Q(\registers[14][2] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][30]$_SDFFCE_PN0P_  (.D(_0281_),
    .DE(_0026_),
    .Q(\registers[14][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][31]$_SDFFCE_PN0P_  (.D(_0282_),
    .DE(_0026_),
    .Q(\registers[14][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][3]$_SDFFCE_PN0P_  (.D(_0283_),
    .DE(_0026_),
    .Q(\registers[14][3] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][4]$_SDFFCE_PN0P_  (.D(_0284_),
    .DE(_0026_),
    .Q(\registers[14][4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][5]$_SDFFCE_PN0P_  (.D(_0285_),
    .DE(_0026_),
    .Q(\registers[14][5] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][6]$_SDFFCE_PN0P_  (.D(_0286_),
    .DE(_0026_),
    .Q(\registers[14][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][7]$_SDFFCE_PN0P_  (.D(_0287_),
    .DE(_0026_),
    .Q(\registers[14][7] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][8]$_SDFFCE_PN0P_  (.D(_0288_),
    .DE(_0026_),
    .Q(\registers[14][8] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[14][9]$_SDFFCE_PN0P_  (.D(_0289_),
    .DE(_0026_),
    .Q(\registers[14][9] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][0]$_SDFFCE_PN0P_  (.D(_0290_),
    .DE(net120),
    .Q(\registers[15][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][10]$_SDFFCE_PN0P_  (.D(_0291_),
    .DE(net120),
    .Q(\registers[15][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][11]$_SDFFCE_PN0P_  (.D(_0292_),
    .DE(net120),
    .Q(\registers[15][11] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][12]$_SDFFCE_PN0P_  (.D(_0293_),
    .DE(net120),
    .Q(\registers[15][12] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][13]$_SDFFCE_PN0P_  (.D(_0294_),
    .DE(net120),
    .Q(\registers[15][13] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][14]$_SDFFCE_PN0P_  (.D(_0295_),
    .DE(net120),
    .Q(\registers[15][14] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][15]$_SDFFCE_PN0P_  (.D(_0296_),
    .DE(net120),
    .Q(\registers[15][15] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][16]$_SDFFCE_PN0P_  (.D(_0297_),
    .DE(net120),
    .Q(\registers[15][16] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][17]$_SDFFCE_PN0P_  (.D(_0298_),
    .DE(net120),
    .Q(\registers[15][17] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][18]$_SDFFCE_PN0P_  (.D(_0299_),
    .DE(net120),
    .Q(\registers[15][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][19]$_SDFFCE_PN0P_  (.D(_0300_),
    .DE(net120),
    .Q(\registers[15][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][1]$_SDFFCE_PN0P_  (.D(_0301_),
    .DE(net120),
    .Q(\registers[15][1] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][20]$_SDFFCE_PN0P_  (.D(_0302_),
    .DE(net120),
    .Q(\registers[15][20] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][21]$_SDFFCE_PN0P_  (.D(_0303_),
    .DE(net120),
    .Q(\registers[15][21] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][22]$_SDFFCE_PN0P_  (.D(_0304_),
    .DE(net120),
    .Q(\registers[15][22] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][23]$_SDFFCE_PN0P_  (.D(_0305_),
    .DE(net120),
    .Q(\registers[15][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][24]$_SDFFCE_PN0P_  (.D(_0306_),
    .DE(net120),
    .Q(\registers[15][24] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][25]$_SDFFCE_PN0P_  (.D(_0307_),
    .DE(net120),
    .Q(\registers[15][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][26]$_SDFFCE_PN0P_  (.D(_0308_),
    .DE(net120),
    .Q(\registers[15][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][27]$_SDFFCE_PN0P_  (.D(_0309_),
    .DE(net120),
    .Q(\registers[15][27] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][28]$_SDFFCE_PN0P_  (.D(_0310_),
    .DE(_0025_),
    .Q(\registers[15][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][29]$_SDFFCE_PN0P_  (.D(_0311_),
    .DE(net120),
    .Q(\registers[15][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][2]$_SDFFCE_PN0P_  (.D(_0312_),
    .DE(_0025_),
    .Q(\registers[15][2] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][30]$_SDFFCE_PN0P_  (.D(_0313_),
    .DE(_0025_),
    .Q(\registers[15][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][31]$_SDFFCE_PN0P_  (.D(_0314_),
    .DE(_0025_),
    .Q(\registers[15][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][3]$_SDFFCE_PN0P_  (.D(_0315_),
    .DE(_0025_),
    .Q(\registers[15][3] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][4]$_SDFFCE_PN0P_  (.D(_0316_),
    .DE(_0025_),
    .Q(\registers[15][4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][5]$_SDFFCE_PN0P_  (.D(_0317_),
    .DE(_0025_),
    .Q(\registers[15][5] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][6]$_SDFFCE_PN0P_  (.D(_0318_),
    .DE(_0025_),
    .Q(\registers[15][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][7]$_SDFFCE_PN0P_  (.D(_0319_),
    .DE(_0025_),
    .Q(\registers[15][7] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][8]$_SDFFCE_PN0P_  (.D(_0320_),
    .DE(_0025_),
    .Q(\registers[15][8] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[15][9]$_SDFFCE_PN0P_  (.D(_0321_),
    .DE(_0025_),
    .Q(\registers[15][9] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][0]$_SDFFCE_PN0P_  (.D(_0322_),
    .DE(_0024_),
    .Q(\registers[16][0] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][10]$_SDFFCE_PN0P_  (.D(_0323_),
    .DE(_0024_),
    .Q(\registers[16][10] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][11]$_SDFFCE_PN0P_  (.D(_0324_),
    .DE(_0024_),
    .Q(\registers[16][11] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][12]$_SDFFCE_PN0P_  (.D(_0325_),
    .DE(_0024_),
    .Q(\registers[16][12] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][13]$_SDFFCE_PN0P_  (.D(_0326_),
    .DE(_0024_),
    .Q(\registers[16][13] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][14]$_SDFFCE_PN0P_  (.D(_0327_),
    .DE(_0024_),
    .Q(\registers[16][14] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][15]$_SDFFCE_PN0P_  (.D(_0328_),
    .DE(_0024_),
    .Q(\registers[16][15] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][16]$_SDFFCE_PN0P_  (.D(_0329_),
    .DE(_0024_),
    .Q(\registers[16][16] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][17]$_SDFFCE_PN0P_  (.D(_0330_),
    .DE(_0024_),
    .Q(\registers[16][17] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][18]$_SDFFCE_PN0P_  (.D(_0331_),
    .DE(_0024_),
    .Q(\registers[16][18] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][19]$_SDFFCE_PN0P_  (.D(_0332_),
    .DE(_0024_),
    .Q(\registers[16][19] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][1]$_SDFFCE_PN0P_  (.D(_0333_),
    .DE(_0024_),
    .Q(\registers[16][1] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][20]$_SDFFCE_PN0P_  (.D(_0334_),
    .DE(_0024_),
    .Q(\registers[16][20] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][21]$_SDFFCE_PN0P_  (.D(_0335_),
    .DE(_0024_),
    .Q(\registers[16][21] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][22]$_SDFFCE_PN0P_  (.D(_0336_),
    .DE(_0024_),
    .Q(\registers[16][22] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][23]$_SDFFCE_PN0P_  (.D(_0337_),
    .DE(_0024_),
    .Q(\registers[16][23] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][24]$_SDFFCE_PN0P_  (.D(_0338_),
    .DE(_0024_),
    .Q(\registers[16][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][25]$_SDFFCE_PN0P_  (.D(_0339_),
    .DE(_0024_),
    .Q(\registers[16][25] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][26]$_SDFFCE_PN0P_  (.D(_0340_),
    .DE(_0024_),
    .Q(\registers[16][26] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][27]$_SDFFCE_PN0P_  (.D(_0341_),
    .DE(_0024_),
    .Q(\registers[16][27] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][28]$_SDFFCE_PN0P_  (.D(_0342_),
    .DE(_0024_),
    .Q(\registers[16][28] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][29]$_SDFFCE_PN0P_  (.D(_0343_),
    .DE(_0024_),
    .Q(\registers[16][29] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][2]$_SDFFCE_PN0P_  (.D(_0344_),
    .DE(_0024_),
    .Q(\registers[16][2] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][30]$_SDFFCE_PN0P_  (.D(_0345_),
    .DE(_0024_),
    .Q(\registers[16][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][31]$_SDFFCE_PN0P_  (.D(_0346_),
    .DE(_0024_),
    .Q(\registers[16][31] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][3]$_SDFFCE_PN0P_  (.D(_0347_),
    .DE(_0024_),
    .Q(\registers[16][3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][4]$_SDFFCE_PN0P_  (.D(_0348_),
    .DE(_0024_),
    .Q(\registers[16][4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][5]$_SDFFCE_PN0P_  (.D(_0349_),
    .DE(_0024_),
    .Q(\registers[16][5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][6]$_SDFFCE_PN0P_  (.D(_0350_),
    .DE(_0024_),
    .Q(\registers[16][6] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][7]$_SDFFCE_PN0P_  (.D(_0351_),
    .DE(_0024_),
    .Q(\registers[16][7] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][8]$_SDFFCE_PN0P_  (.D(_0352_),
    .DE(_0024_),
    .Q(\registers[16][8] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[16][9]$_SDFFCE_PN0P_  (.D(_0353_),
    .DE(_0024_),
    .Q(\registers[16][9] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][0]$_SDFFCE_PN0P_  (.D(_0354_),
    .DE(_0023_),
    .Q(\registers[17][0] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][10]$_SDFFCE_PN0P_  (.D(_0355_),
    .DE(_0023_),
    .Q(\registers[17][10] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][11]$_SDFFCE_PN0P_  (.D(_0356_),
    .DE(_0023_),
    .Q(\registers[17][11] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][12]$_SDFFCE_PN0P_  (.D(_0357_),
    .DE(_0023_),
    .Q(\registers[17][12] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][13]$_SDFFCE_PN0P_  (.D(_0358_),
    .DE(_0023_),
    .Q(\registers[17][13] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][14]$_SDFFCE_PN0P_  (.D(_0359_),
    .DE(_0023_),
    .Q(\registers[17][14] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][15]$_SDFFCE_PN0P_  (.D(_0360_),
    .DE(_0023_),
    .Q(\registers[17][15] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][16]$_SDFFCE_PN0P_  (.D(_0361_),
    .DE(_0023_),
    .Q(\registers[17][16] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][17]$_SDFFCE_PN0P_  (.D(_0362_),
    .DE(_0023_),
    .Q(\registers[17][17] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][18]$_SDFFCE_PN0P_  (.D(_0363_),
    .DE(_0023_),
    .Q(\registers[17][18] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][19]$_SDFFCE_PN0P_  (.D(_0364_),
    .DE(_0023_),
    .Q(\registers[17][19] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][1]$_SDFFCE_PN0P_  (.D(_0365_),
    .DE(_0023_),
    .Q(\registers[17][1] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][20]$_SDFFCE_PN0P_  (.D(_0366_),
    .DE(_0023_),
    .Q(\registers[17][20] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][21]$_SDFFCE_PN0P_  (.D(_0367_),
    .DE(_0023_),
    .Q(\registers[17][21] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][22]$_SDFFCE_PN0P_  (.D(_0368_),
    .DE(_0023_),
    .Q(\registers[17][22] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][23]$_SDFFCE_PN0P_  (.D(_0369_),
    .DE(_0023_),
    .Q(\registers[17][23] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][24]$_SDFFCE_PN0P_  (.D(_0370_),
    .DE(_0023_),
    .Q(\registers[17][24] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][25]$_SDFFCE_PN0P_  (.D(_0371_),
    .DE(_0023_),
    .Q(\registers[17][25] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][26]$_SDFFCE_PN0P_  (.D(_0372_),
    .DE(_0023_),
    .Q(\registers[17][26] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][27]$_SDFFCE_PN0P_  (.D(_0373_),
    .DE(_0023_),
    .Q(\registers[17][27] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][28]$_SDFFCE_PN0P_  (.D(_0374_),
    .DE(_0023_),
    .Q(\registers[17][28] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][29]$_SDFFCE_PN0P_  (.D(_0375_),
    .DE(_0023_),
    .Q(\registers[17][29] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][2]$_SDFFCE_PN0P_  (.D(_0376_),
    .DE(_0023_),
    .Q(\registers[17][2] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][30]$_SDFFCE_PN0P_  (.D(_0377_),
    .DE(_0023_),
    .Q(\registers[17][30] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][31]$_SDFFCE_PN0P_  (.D(_0378_),
    .DE(_0023_),
    .Q(\registers[17][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][3]$_SDFFCE_PN0P_  (.D(_0379_),
    .DE(_0023_),
    .Q(\registers[17][3] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][4]$_SDFFCE_PN0P_  (.D(_0380_),
    .DE(_0023_),
    .Q(\registers[17][4] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][5]$_SDFFCE_PN0P_  (.D(_0381_),
    .DE(_0023_),
    .Q(\registers[17][5] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][6]$_SDFFCE_PN0P_  (.D(_0382_),
    .DE(_0023_),
    .Q(\registers[17][6] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][7]$_SDFFCE_PN0P_  (.D(_0383_),
    .DE(_0023_),
    .Q(\registers[17][7] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][8]$_SDFFCE_PN0P_  (.D(_0384_),
    .DE(_0023_),
    .Q(\registers[17][8] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[17][9]$_SDFFCE_PN0P_  (.D(_0385_),
    .DE(_0023_),
    .Q(\registers[17][9] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][0]$_SDFFCE_PN0P_  (.D(_0386_),
    .DE(_0022_),
    .Q(\registers[18][0] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][10]$_SDFFCE_PN0P_  (.D(_0387_),
    .DE(_0022_),
    .Q(\registers[18][10] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][11]$_SDFFCE_PN0P_  (.D(_0388_),
    .DE(_0022_),
    .Q(\registers[18][11] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][12]$_SDFFCE_PN0P_  (.D(_0389_),
    .DE(_0022_),
    .Q(\registers[18][12] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][13]$_SDFFCE_PN0P_  (.D(_0390_),
    .DE(_0022_),
    .Q(\registers[18][13] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][14]$_SDFFCE_PN0P_  (.D(_0391_),
    .DE(_0022_),
    .Q(\registers[18][14] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][15]$_SDFFCE_PN0P_  (.D(_0392_),
    .DE(_0022_),
    .Q(\registers[18][15] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][16]$_SDFFCE_PN0P_  (.D(_0393_),
    .DE(_0022_),
    .Q(\registers[18][16] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][17]$_SDFFCE_PN0P_  (.D(_0394_),
    .DE(_0022_),
    .Q(\registers[18][17] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][18]$_SDFFCE_PN0P_  (.D(_0395_),
    .DE(_0022_),
    .Q(\registers[18][18] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][19]$_SDFFCE_PN0P_  (.D(_0396_),
    .DE(_0022_),
    .Q(\registers[18][19] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][1]$_SDFFCE_PN0P_  (.D(_0397_),
    .DE(_0022_),
    .Q(\registers[18][1] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][20]$_SDFFCE_PN0P_  (.D(_0398_),
    .DE(_0022_),
    .Q(\registers[18][20] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][21]$_SDFFCE_PN0P_  (.D(_0399_),
    .DE(_0022_),
    .Q(\registers[18][21] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][22]$_SDFFCE_PN0P_  (.D(_0400_),
    .DE(_0022_),
    .Q(\registers[18][22] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][23]$_SDFFCE_PN0P_  (.D(_0401_),
    .DE(_0022_),
    .Q(\registers[18][23] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][24]$_SDFFCE_PN0P_  (.D(_0402_),
    .DE(_0022_),
    .Q(\registers[18][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][25]$_SDFFCE_PN0P_  (.D(_0403_),
    .DE(_0022_),
    .Q(\registers[18][25] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][26]$_SDFFCE_PN0P_  (.D(_0404_),
    .DE(_0022_),
    .Q(\registers[18][26] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][27]$_SDFFCE_PN0P_  (.D(_0405_),
    .DE(_0022_),
    .Q(\registers[18][27] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][28]$_SDFFCE_PN0P_  (.D(_0406_),
    .DE(_0022_),
    .Q(\registers[18][28] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][29]$_SDFFCE_PN0P_  (.D(_0407_),
    .DE(_0022_),
    .Q(\registers[18][29] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][2]$_SDFFCE_PN0P_  (.D(_0408_),
    .DE(_0022_),
    .Q(\registers[18][2] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][30]$_SDFFCE_PN0P_  (.D(_0409_),
    .DE(_0022_),
    .Q(\registers[18][30] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][31]$_SDFFCE_PN0P_  (.D(_0410_),
    .DE(_0022_),
    .Q(\registers[18][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][3]$_SDFFCE_PN0P_  (.D(_0411_),
    .DE(_0022_),
    .Q(\registers[18][3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][4]$_SDFFCE_PN0P_  (.D(_0412_),
    .DE(_0022_),
    .Q(\registers[18][4] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][5]$_SDFFCE_PN0P_  (.D(_0413_),
    .DE(_0022_),
    .Q(\registers[18][5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][6]$_SDFFCE_PN0P_  (.D(_0414_),
    .DE(_0022_),
    .Q(\registers[18][6] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][7]$_SDFFCE_PN0P_  (.D(_0415_),
    .DE(_0022_),
    .Q(\registers[18][7] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][8]$_SDFFCE_PN0P_  (.D(_0416_),
    .DE(_0022_),
    .Q(\registers[18][8] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[18][9]$_SDFFCE_PN0P_  (.D(_0417_),
    .DE(_0022_),
    .Q(\registers[18][9] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][0]$_SDFFCE_PN0P_  (.D(_0418_),
    .DE(_0021_),
    .Q(\registers[19][0] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][10]$_SDFFCE_PN0P_  (.D(_0419_),
    .DE(_0021_),
    .Q(\registers[19][10] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][11]$_SDFFCE_PN0P_  (.D(_0420_),
    .DE(_0021_),
    .Q(\registers[19][11] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][12]$_SDFFCE_PN0P_  (.D(_0421_),
    .DE(_0021_),
    .Q(\registers[19][12] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][13]$_SDFFCE_PN0P_  (.D(_0422_),
    .DE(_0021_),
    .Q(\registers[19][13] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][14]$_SDFFCE_PN0P_  (.D(_0423_),
    .DE(_0021_),
    .Q(\registers[19][14] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][15]$_SDFFCE_PN0P_  (.D(_0424_),
    .DE(_0021_),
    .Q(\registers[19][15] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][16]$_SDFFCE_PN0P_  (.D(_0425_),
    .DE(_0021_),
    .Q(\registers[19][16] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][17]$_SDFFCE_PN0P_  (.D(_0426_),
    .DE(_0021_),
    .Q(\registers[19][17] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][18]$_SDFFCE_PN0P_  (.D(_0427_),
    .DE(_0021_),
    .Q(\registers[19][18] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][19]$_SDFFCE_PN0P_  (.D(_0428_),
    .DE(_0021_),
    .Q(\registers[19][19] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][1]$_SDFFCE_PN0P_  (.D(_0429_),
    .DE(_0021_),
    .Q(\registers[19][1] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][20]$_SDFFCE_PN0P_  (.D(_0430_),
    .DE(_0021_),
    .Q(\registers[19][20] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][21]$_SDFFCE_PN0P_  (.D(_0431_),
    .DE(_0021_),
    .Q(\registers[19][21] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][22]$_SDFFCE_PN0P_  (.D(_0432_),
    .DE(_0021_),
    .Q(\registers[19][22] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][23]$_SDFFCE_PN0P_  (.D(_0433_),
    .DE(_0021_),
    .Q(\registers[19][23] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][24]$_SDFFCE_PN0P_  (.D(_0434_),
    .DE(_0021_),
    .Q(\registers[19][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][25]$_SDFFCE_PN0P_  (.D(_0435_),
    .DE(_0021_),
    .Q(\registers[19][25] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][26]$_SDFFCE_PN0P_  (.D(_0436_),
    .DE(_0021_),
    .Q(\registers[19][26] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][27]$_SDFFCE_PN0P_  (.D(_0437_),
    .DE(_0021_),
    .Q(\registers[19][27] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][28]$_SDFFCE_PN0P_  (.D(_0438_),
    .DE(_0021_),
    .Q(\registers[19][28] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][29]$_SDFFCE_PN0P_  (.D(_0439_),
    .DE(_0021_),
    .Q(\registers[19][29] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][2]$_SDFFCE_PN0P_  (.D(_0440_),
    .DE(_0021_),
    .Q(\registers[19][2] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][30]$_SDFFCE_PN0P_  (.D(_0441_),
    .DE(_0021_),
    .Q(\registers[19][30] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][31]$_SDFFCE_PN0P_  (.D(_0442_),
    .DE(_0021_),
    .Q(\registers[19][31] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][3]$_SDFFCE_PN0P_  (.D(_0443_),
    .DE(_0021_),
    .Q(\registers[19][3] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][4]$_SDFFCE_PN0P_  (.D(_0444_),
    .DE(_0021_),
    .Q(\registers[19][4] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][5]$_SDFFCE_PN0P_  (.D(_0445_),
    .DE(_0021_),
    .Q(\registers[19][5] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][6]$_SDFFCE_PN0P_  (.D(_0446_),
    .DE(_0021_),
    .Q(\registers[19][6] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][7]$_SDFFCE_PN0P_  (.D(_0447_),
    .DE(_0021_),
    .Q(\registers[19][7] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][8]$_SDFFCE_PN0P_  (.D(_0448_),
    .DE(_0021_),
    .Q(\registers[19][8] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[19][9]$_SDFFCE_PN0P_  (.D(_0449_),
    .DE(_0021_),
    .Q(\registers[19][9] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][0]$_SDFFCE_PN0P_  (.D(_0450_),
    .DE(_0020_),
    .Q(\registers[1][0] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][10]$_SDFFCE_PN0P_  (.D(_0451_),
    .DE(_0020_),
    .Q(\registers[1][10] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][11]$_SDFFCE_PN0P_  (.D(_0452_),
    .DE(_0020_),
    .Q(\registers[1][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][12]$_SDFFCE_PN0P_  (.D(_0453_),
    .DE(_0020_),
    .Q(\registers[1][12] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][13]$_SDFFCE_PN0P_  (.D(_0454_),
    .DE(_0020_),
    .Q(\registers[1][13] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][14]$_SDFFCE_PN0P_  (.D(_0455_),
    .DE(_0020_),
    .Q(\registers[1][14] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][15]$_SDFFCE_PN0P_  (.D(_0456_),
    .DE(_0020_),
    .Q(\registers[1][15] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][16]$_SDFFCE_PN0P_  (.D(_0457_),
    .DE(_0020_),
    .Q(\registers[1][16] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][17]$_SDFFCE_PN0P_  (.D(_0458_),
    .DE(net131),
    .Q(\registers[1][17] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][18]$_SDFFCE_PN0P_  (.D(_0459_),
    .DE(_0020_),
    .Q(\registers[1][18] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][19]$_SDFFCE_PN0P_  (.D(_0460_),
    .DE(net131),
    .Q(\registers[1][19] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][1]$_SDFFCE_PN0P_  (.D(_0461_),
    .DE(net131),
    .Q(\registers[1][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][20]$_SDFFCE_PN0P_  (.D(_0462_),
    .DE(net131),
    .Q(\registers[1][20] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][21]$_SDFFCE_PN0P_  (.D(_0463_),
    .DE(net131),
    .Q(\registers[1][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][22]$_SDFFCE_PN0P_  (.D(_0464_),
    .DE(net131),
    .Q(\registers[1][22] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][23]$_SDFFCE_PN0P_  (.D(_0465_),
    .DE(net131),
    .Q(\registers[1][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][24]$_SDFFCE_PN0P_  (.D(_0466_),
    .DE(net131),
    .Q(\registers[1][24] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][25]$_SDFFCE_PN0P_  (.D(_0467_),
    .DE(net131),
    .Q(\registers[1][25] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][26]$_SDFFCE_PN0P_  (.D(_0468_),
    .DE(net131),
    .Q(\registers[1][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][27]$_SDFFCE_PN0P_  (.D(_0469_),
    .DE(net131),
    .Q(\registers[1][27] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][28]$_SDFFCE_PN0P_  (.D(_0470_),
    .DE(_0020_),
    .Q(\registers[1][28] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][29]$_SDFFCE_PN0P_  (.D(_0471_),
    .DE(net131),
    .Q(\registers[1][29] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][2]$_SDFFCE_PN0P_  (.D(_0472_),
    .DE(net131),
    .Q(\registers[1][2] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][30]$_SDFFCE_PN0P_  (.D(_0473_),
    .DE(net131),
    .Q(\registers[1][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][31]$_SDFFCE_PN0P_  (.D(_0474_),
    .DE(_0020_),
    .Q(\registers[1][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][3]$_SDFFCE_PN0P_  (.D(_0475_),
    .DE(_0020_),
    .Q(\registers[1][3] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][4]$_SDFFCE_PN0P_  (.D(_0476_),
    .DE(_0020_),
    .Q(\registers[1][4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][5]$_SDFFCE_PN0P_  (.D(_0477_),
    .DE(_0020_),
    .Q(\registers[1][5] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][6]$_SDFFCE_PN0P_  (.D(_0478_),
    .DE(_0020_),
    .Q(\registers[1][6] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][7]$_SDFFCE_PN0P_  (.D(_0479_),
    .DE(_0020_),
    .Q(\registers[1][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][8]$_SDFFCE_PN0P_  (.D(_0480_),
    .DE(_0020_),
    .Q(\registers[1][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[1][9]$_SDFFCE_PN0P_  (.D(_0481_),
    .DE(net131),
    .Q(\registers[1][9] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][0]$_SDFFCE_PN0P_  (.D(_0482_),
    .DE(_0019_),
    .Q(\registers[20][0] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][10]$_SDFFCE_PN0P_  (.D(_0483_),
    .DE(_0019_),
    .Q(\registers[20][10] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][11]$_SDFFCE_PN0P_  (.D(_0484_),
    .DE(_0019_),
    .Q(\registers[20][11] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][12]$_SDFFCE_PN0P_  (.D(_0485_),
    .DE(_0019_),
    .Q(\registers[20][12] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][13]$_SDFFCE_PN0P_  (.D(_0486_),
    .DE(_0019_),
    .Q(\registers[20][13] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][14]$_SDFFCE_PN0P_  (.D(_0487_),
    .DE(_0019_),
    .Q(\registers[20][14] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][15]$_SDFFCE_PN0P_  (.D(_0488_),
    .DE(_0019_),
    .Q(\registers[20][15] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][16]$_SDFFCE_PN0P_  (.D(_0489_),
    .DE(_0019_),
    .Q(\registers[20][16] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][17]$_SDFFCE_PN0P_  (.D(_0490_),
    .DE(_0019_),
    .Q(\registers[20][17] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][18]$_SDFFCE_PN0P_  (.D(_0491_),
    .DE(_0019_),
    .Q(\registers[20][18] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][19]$_SDFFCE_PN0P_  (.D(_0492_),
    .DE(_0019_),
    .Q(\registers[20][19] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][1]$_SDFFCE_PN0P_  (.D(_0493_),
    .DE(_0019_),
    .Q(\registers[20][1] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][20]$_SDFFCE_PN0P_  (.D(_0494_),
    .DE(_0019_),
    .Q(\registers[20][20] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][21]$_SDFFCE_PN0P_  (.D(_0495_),
    .DE(_0019_),
    .Q(\registers[20][21] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][22]$_SDFFCE_PN0P_  (.D(_0496_),
    .DE(_0019_),
    .Q(\registers[20][22] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][23]$_SDFFCE_PN0P_  (.D(_0497_),
    .DE(_0019_),
    .Q(\registers[20][23] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][24]$_SDFFCE_PN0P_  (.D(_0498_),
    .DE(_0019_),
    .Q(\registers[20][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][25]$_SDFFCE_PN0P_  (.D(_0499_),
    .DE(_0019_),
    .Q(\registers[20][25] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][26]$_SDFFCE_PN0P_  (.D(_0500_),
    .DE(_0019_),
    .Q(\registers[20][26] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][27]$_SDFFCE_PN0P_  (.D(_0501_),
    .DE(_0019_),
    .Q(\registers[20][27] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][28]$_SDFFCE_PN0P_  (.D(_0502_),
    .DE(_0019_),
    .Q(\registers[20][28] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][29]$_SDFFCE_PN0P_  (.D(_0503_),
    .DE(_0019_),
    .Q(\registers[20][29] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][2]$_SDFFCE_PN0P_  (.D(_0504_),
    .DE(_0019_),
    .Q(\registers[20][2] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][30]$_SDFFCE_PN0P_  (.D(_0505_),
    .DE(_0019_),
    .Q(\registers[20][30] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][31]$_SDFFCE_PN0P_  (.D(_0506_),
    .DE(_0019_),
    .Q(\registers[20][31] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][3]$_SDFFCE_PN0P_  (.D(_0507_),
    .DE(_0019_),
    .Q(\registers[20][3] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][4]$_SDFFCE_PN0P_  (.D(_0508_),
    .DE(_0019_),
    .Q(\registers[20][4] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][5]$_SDFFCE_PN0P_  (.D(_0509_),
    .DE(_0019_),
    .Q(\registers[20][5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][6]$_SDFFCE_PN0P_  (.D(_0510_),
    .DE(_0019_),
    .Q(\registers[20][6] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][7]$_SDFFCE_PN0P_  (.D(_0511_),
    .DE(_0019_),
    .Q(\registers[20][7] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][8]$_SDFFCE_PN0P_  (.D(_0512_),
    .DE(_0019_),
    .Q(\registers[20][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[20][9]$_SDFFCE_PN0P_  (.D(_0513_),
    .DE(_0019_),
    .Q(\registers[20][9] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][0]$_SDFFCE_PN0P_  (.D(_0514_),
    .DE(_0018_),
    .Q(\registers[21][0] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][10]$_SDFFCE_PN0P_  (.D(_0515_),
    .DE(_0018_),
    .Q(\registers[21][10] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][11]$_SDFFCE_PN0P_  (.D(_0516_),
    .DE(_0018_),
    .Q(\registers[21][11] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][12]$_SDFFCE_PN0P_  (.D(_0517_),
    .DE(_0018_),
    .Q(\registers[21][12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][13]$_SDFFCE_PN0P_  (.D(_0518_),
    .DE(_0018_),
    .Q(\registers[21][13] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][14]$_SDFFCE_PN0P_  (.D(_0519_),
    .DE(_0018_),
    .Q(\registers[21][14] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][15]$_SDFFCE_PN0P_  (.D(_0520_),
    .DE(_0018_),
    .Q(\registers[21][15] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][16]$_SDFFCE_PN0P_  (.D(_0521_),
    .DE(_0018_),
    .Q(\registers[21][16] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][17]$_SDFFCE_PN0P_  (.D(_0522_),
    .DE(_0018_),
    .Q(\registers[21][17] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][18]$_SDFFCE_PN0P_  (.D(_0523_),
    .DE(_0018_),
    .Q(\registers[21][18] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][19]$_SDFFCE_PN0P_  (.D(_0524_),
    .DE(_0018_),
    .Q(\registers[21][19] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][1]$_SDFFCE_PN0P_  (.D(_0525_),
    .DE(_0018_),
    .Q(\registers[21][1] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][20]$_SDFFCE_PN0P_  (.D(_0526_),
    .DE(_0018_),
    .Q(\registers[21][20] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][21]$_SDFFCE_PN0P_  (.D(_0527_),
    .DE(_0018_),
    .Q(\registers[21][21] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][22]$_SDFFCE_PN0P_  (.D(_0528_),
    .DE(_0018_),
    .Q(\registers[21][22] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][23]$_SDFFCE_PN0P_  (.D(_0529_),
    .DE(_0018_),
    .Q(\registers[21][23] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][24]$_SDFFCE_PN0P_  (.D(_0530_),
    .DE(_0018_),
    .Q(\registers[21][24] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][25]$_SDFFCE_PN0P_  (.D(_0531_),
    .DE(_0018_),
    .Q(\registers[21][25] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][26]$_SDFFCE_PN0P_  (.D(_0532_),
    .DE(_0018_),
    .Q(\registers[21][26] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][27]$_SDFFCE_PN0P_  (.D(_0533_),
    .DE(_0018_),
    .Q(\registers[21][27] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][28]$_SDFFCE_PN0P_  (.D(_0534_),
    .DE(_0018_),
    .Q(\registers[21][28] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][29]$_SDFFCE_PN0P_  (.D(_0535_),
    .DE(_0018_),
    .Q(\registers[21][29] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][2]$_SDFFCE_PN0P_  (.D(_0536_),
    .DE(_0018_),
    .Q(\registers[21][2] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][30]$_SDFFCE_PN0P_  (.D(_0537_),
    .DE(_0018_),
    .Q(\registers[21][30] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][31]$_SDFFCE_PN0P_  (.D(_0538_),
    .DE(_0018_),
    .Q(\registers[21][31] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][3]$_SDFFCE_PN0P_  (.D(_0539_),
    .DE(_0018_),
    .Q(\registers[21][3] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][4]$_SDFFCE_PN0P_  (.D(_0540_),
    .DE(_0018_),
    .Q(\registers[21][4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][5]$_SDFFCE_PN0P_  (.D(_0541_),
    .DE(_0018_),
    .Q(\registers[21][5] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][6]$_SDFFCE_PN0P_  (.D(_0542_),
    .DE(_0018_),
    .Q(\registers[21][6] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][7]$_SDFFCE_PN0P_  (.D(_0543_),
    .DE(_0018_),
    .Q(\registers[21][7] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][8]$_SDFFCE_PN0P_  (.D(_0544_),
    .DE(_0018_),
    .Q(\registers[21][8] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[21][9]$_SDFFCE_PN0P_  (.D(_0545_),
    .DE(_0018_),
    .Q(\registers[21][9] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][0]$_SDFFCE_PN0P_  (.D(_0546_),
    .DE(_0017_),
    .Q(\registers[22][0] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][10]$_SDFFCE_PN0P_  (.D(_0547_),
    .DE(_0017_),
    .Q(\registers[22][10] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][11]$_SDFFCE_PN0P_  (.D(_0548_),
    .DE(_0017_),
    .Q(\registers[22][11] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][12]$_SDFFCE_PN0P_  (.D(_0549_),
    .DE(_0017_),
    .Q(\registers[22][12] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][13]$_SDFFCE_PN0P_  (.D(_0550_),
    .DE(_0017_),
    .Q(\registers[22][13] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][14]$_SDFFCE_PN0P_  (.D(_0551_),
    .DE(_0017_),
    .Q(\registers[22][14] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][15]$_SDFFCE_PN0P_  (.D(_0552_),
    .DE(_0017_),
    .Q(\registers[22][15] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][16]$_SDFFCE_PN0P_  (.D(_0553_),
    .DE(_0017_),
    .Q(\registers[22][16] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][17]$_SDFFCE_PN0P_  (.D(_0554_),
    .DE(_0017_),
    .Q(\registers[22][17] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][18]$_SDFFCE_PN0P_  (.D(_0555_),
    .DE(_0017_),
    .Q(\registers[22][18] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][19]$_SDFFCE_PN0P_  (.D(_0556_),
    .DE(_0017_),
    .Q(\registers[22][19] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][1]$_SDFFCE_PN0P_  (.D(_0557_),
    .DE(_0017_),
    .Q(\registers[22][1] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][20]$_SDFFCE_PN0P_  (.D(_0558_),
    .DE(_0017_),
    .Q(\registers[22][20] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][21]$_SDFFCE_PN0P_  (.D(_0559_),
    .DE(_0017_),
    .Q(\registers[22][21] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][22]$_SDFFCE_PN0P_  (.D(_0560_),
    .DE(_0017_),
    .Q(\registers[22][22] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][23]$_SDFFCE_PN0P_  (.D(_0561_),
    .DE(_0017_),
    .Q(\registers[22][23] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][24]$_SDFFCE_PN0P_  (.D(_0562_),
    .DE(_0017_),
    .Q(\registers[22][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][25]$_SDFFCE_PN0P_  (.D(_0563_),
    .DE(_0017_),
    .Q(\registers[22][25] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][26]$_SDFFCE_PN0P_  (.D(_0564_),
    .DE(_0017_),
    .Q(\registers[22][26] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][27]$_SDFFCE_PN0P_  (.D(_0565_),
    .DE(_0017_),
    .Q(\registers[22][27] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][28]$_SDFFCE_PN0P_  (.D(_0566_),
    .DE(_0017_),
    .Q(\registers[22][28] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][29]$_SDFFCE_PN0P_  (.D(_0567_),
    .DE(_0017_),
    .Q(\registers[22][29] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][2]$_SDFFCE_PN0P_  (.D(_0568_),
    .DE(_0017_),
    .Q(\registers[22][2] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][30]$_SDFFCE_PN0P_  (.D(_0569_),
    .DE(_0017_),
    .Q(\registers[22][30] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][31]$_SDFFCE_PN0P_  (.D(_0570_),
    .DE(_0017_),
    .Q(\registers[22][31] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][3]$_SDFFCE_PN0P_  (.D(_0571_),
    .DE(_0017_),
    .Q(\registers[22][3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][4]$_SDFFCE_PN0P_  (.D(_0572_),
    .DE(_0017_),
    .Q(\registers[22][4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][5]$_SDFFCE_PN0P_  (.D(_0573_),
    .DE(_0017_),
    .Q(\registers[22][5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][6]$_SDFFCE_PN0P_  (.D(_0574_),
    .DE(_0017_),
    .Q(\registers[22][6] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][7]$_SDFFCE_PN0P_  (.D(_0575_),
    .DE(_0017_),
    .Q(\registers[22][7] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][8]$_SDFFCE_PN0P_  (.D(_0576_),
    .DE(_0017_),
    .Q(\registers[22][8] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[22][9]$_SDFFCE_PN0P_  (.D(_0577_),
    .DE(_0017_),
    .Q(\registers[22][9] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][0]$_SDFFCE_PN0P_  (.D(_0578_),
    .DE(_0016_),
    .Q(\registers[23][0] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][10]$_SDFFCE_PN0P_  (.D(_0579_),
    .DE(_0016_),
    .Q(\registers[23][10] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][11]$_SDFFCE_PN0P_  (.D(_0580_),
    .DE(_0016_),
    .Q(\registers[23][11] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][12]$_SDFFCE_PN0P_  (.D(_0581_),
    .DE(_0016_),
    .Q(\registers[23][12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][13]$_SDFFCE_PN0P_  (.D(_0582_),
    .DE(_0016_),
    .Q(\registers[23][13] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][14]$_SDFFCE_PN0P_  (.D(_0583_),
    .DE(_0016_),
    .Q(\registers[23][14] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][15]$_SDFFCE_PN0P_  (.D(_0584_),
    .DE(_0016_),
    .Q(\registers[23][15] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][16]$_SDFFCE_PN0P_  (.D(_0585_),
    .DE(_0016_),
    .Q(\registers[23][16] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][17]$_SDFFCE_PN0P_  (.D(_0586_),
    .DE(_0016_),
    .Q(\registers[23][17] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][18]$_SDFFCE_PN0P_  (.D(_0587_),
    .DE(_0016_),
    .Q(\registers[23][18] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][19]$_SDFFCE_PN0P_  (.D(_0588_),
    .DE(_0016_),
    .Q(\registers[23][19] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][1]$_SDFFCE_PN0P_  (.D(_0589_),
    .DE(_0016_),
    .Q(\registers[23][1] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][20]$_SDFFCE_PN0P_  (.D(_0590_),
    .DE(_0016_),
    .Q(\registers[23][20] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][21]$_SDFFCE_PN0P_  (.D(_0591_),
    .DE(_0016_),
    .Q(\registers[23][21] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][22]$_SDFFCE_PN0P_  (.D(_0592_),
    .DE(_0016_),
    .Q(\registers[23][22] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][23]$_SDFFCE_PN0P_  (.D(_0593_),
    .DE(_0016_),
    .Q(\registers[23][23] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][24]$_SDFFCE_PN0P_  (.D(_0594_),
    .DE(_0016_),
    .Q(\registers[23][24] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][25]$_SDFFCE_PN0P_  (.D(_0595_),
    .DE(_0016_),
    .Q(\registers[23][25] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][26]$_SDFFCE_PN0P_  (.D(_0596_),
    .DE(_0016_),
    .Q(\registers[23][26] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][27]$_SDFFCE_PN0P_  (.D(_0597_),
    .DE(_0016_),
    .Q(\registers[23][27] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][28]$_SDFFCE_PN0P_  (.D(_0598_),
    .DE(_0016_),
    .Q(\registers[23][28] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][29]$_SDFFCE_PN0P_  (.D(_0599_),
    .DE(_0016_),
    .Q(\registers[23][29] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][2]$_SDFFCE_PN0P_  (.D(_0600_),
    .DE(_0016_),
    .Q(\registers[23][2] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][30]$_SDFFCE_PN0P_  (.D(_0601_),
    .DE(_0016_),
    .Q(\registers[23][30] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][31]$_SDFFCE_PN0P_  (.D(_0602_),
    .DE(_0016_),
    .Q(\registers[23][31] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][3]$_SDFFCE_PN0P_  (.D(_0603_),
    .DE(_0016_),
    .Q(\registers[23][3] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][4]$_SDFFCE_PN0P_  (.D(_0604_),
    .DE(_0016_),
    .Q(\registers[23][4] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][5]$_SDFFCE_PN0P_  (.D(_0605_),
    .DE(_0016_),
    .Q(\registers[23][5] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][6]$_SDFFCE_PN0P_  (.D(_0606_),
    .DE(_0016_),
    .Q(\registers[23][6] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][7]$_SDFFCE_PN0P_  (.D(_0607_),
    .DE(_0016_),
    .Q(\registers[23][7] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][8]$_SDFFCE_PN0P_  (.D(_0608_),
    .DE(_0016_),
    .Q(\registers[23][8] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[23][9]$_SDFFCE_PN0P_  (.D(_0609_),
    .DE(_0016_),
    .Q(\registers[23][9] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][0]$_SDFFCE_PN0P_  (.D(_0610_),
    .DE(_0015_),
    .Q(\registers[24][0] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][10]$_SDFFCE_PN0P_  (.D(_0611_),
    .DE(_0015_),
    .Q(\registers[24][10] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][11]$_SDFFCE_PN0P_  (.D(_0612_),
    .DE(_0015_),
    .Q(\registers[24][11] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][12]$_SDFFCE_PN0P_  (.D(_0613_),
    .DE(_0015_),
    .Q(\registers[24][12] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][13]$_SDFFCE_PN0P_  (.D(_0614_),
    .DE(_0015_),
    .Q(\registers[24][13] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][14]$_SDFFCE_PN0P_  (.D(_0615_),
    .DE(_0015_),
    .Q(\registers[24][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][15]$_SDFFCE_PN0P_  (.D(_0616_),
    .DE(_0015_),
    .Q(\registers[24][15] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][16]$_SDFFCE_PN0P_  (.D(_0617_),
    .DE(_0015_),
    .Q(\registers[24][16] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][17]$_SDFFCE_PN0P_  (.D(_0618_),
    .DE(_0015_),
    .Q(\registers[24][17] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][18]$_SDFFCE_PN0P_  (.D(_0619_),
    .DE(_0015_),
    .Q(\registers[24][18] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][19]$_SDFFCE_PN0P_  (.D(_0620_),
    .DE(_0015_),
    .Q(\registers[24][19] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][1]$_SDFFCE_PN0P_  (.D(_0621_),
    .DE(_0015_),
    .Q(\registers[24][1] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][20]$_SDFFCE_PN0P_  (.D(_0622_),
    .DE(_0015_),
    .Q(\registers[24][20] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][21]$_SDFFCE_PN0P_  (.D(_0623_),
    .DE(_0015_),
    .Q(\registers[24][21] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][22]$_SDFFCE_PN0P_  (.D(_0624_),
    .DE(_0015_),
    .Q(\registers[24][22] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][23]$_SDFFCE_PN0P_  (.D(_0625_),
    .DE(net111),
    .Q(\registers[24][23] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][24]$_SDFFCE_PN0P_  (.D(_0626_),
    .DE(net111),
    .Q(\registers[24][24] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][25]$_SDFFCE_PN0P_  (.D(_0627_),
    .DE(net111),
    .Q(\registers[24][25] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][26]$_SDFFCE_PN0P_  (.D(_0628_),
    .DE(net111),
    .Q(\registers[24][26] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][27]$_SDFFCE_PN0P_  (.D(_0629_),
    .DE(net111),
    .Q(\registers[24][27] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][28]$_SDFFCE_PN0P_  (.D(_0630_),
    .DE(net111),
    .Q(\registers[24][28] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][29]$_SDFFCE_PN0P_  (.D(_0631_),
    .DE(net111),
    .Q(\registers[24][29] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][2]$_SDFFCE_PN0P_  (.D(_0632_),
    .DE(net111),
    .Q(\registers[24][2] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][30]$_SDFFCE_PN0P_  (.D(_0633_),
    .DE(net111),
    .Q(\registers[24][30] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][31]$_SDFFCE_PN0P_  (.D(_0634_),
    .DE(net111),
    .Q(\registers[24][31] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][3]$_SDFFCE_PN0P_  (.D(_0635_),
    .DE(net111),
    .Q(\registers[24][3] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][4]$_SDFFCE_PN0P_  (.D(_0636_),
    .DE(net111),
    .Q(\registers[24][4] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][5]$_SDFFCE_PN0P_  (.D(_0637_),
    .DE(net111),
    .Q(\registers[24][5] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][6]$_SDFFCE_PN0P_  (.D(_0638_),
    .DE(net111),
    .Q(\registers[24][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][7]$_SDFFCE_PN0P_  (.D(_0639_),
    .DE(net111),
    .Q(\registers[24][7] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][8]$_SDFFCE_PN0P_  (.D(_0640_),
    .DE(net111),
    .Q(\registers[24][8] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[24][9]$_SDFFCE_PN0P_  (.D(_0641_),
    .DE(net111),
    .Q(\registers[24][9] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][0]$_SDFFCE_PN0P_  (.D(_0642_),
    .DE(net130),
    .Q(\registers[25][0] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][10]$_SDFFCE_PN0P_  (.D(_0643_),
    .DE(net130),
    .Q(\registers[25][10] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][11]$_SDFFCE_PN0P_  (.D(_0644_),
    .DE(net130),
    .Q(\registers[25][11] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][12]$_SDFFCE_PN0P_  (.D(_0645_),
    .DE(net130),
    .Q(\registers[25][12] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][13]$_SDFFCE_PN0P_  (.D(_0646_),
    .DE(net130),
    .Q(\registers[25][13] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][14]$_SDFFCE_PN0P_  (.D(_0647_),
    .DE(net130),
    .Q(\registers[25][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][15]$_SDFFCE_PN0P_  (.D(_0648_),
    .DE(net130),
    .Q(\registers[25][15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][16]$_SDFFCE_PN0P_  (.D(_0649_),
    .DE(net130),
    .Q(\registers[25][16] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][17]$_SDFFCE_PN0P_  (.D(_0650_),
    .DE(net130),
    .Q(\registers[25][17] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][18]$_SDFFCE_PN0P_  (.D(_0651_),
    .DE(net130),
    .Q(\registers[25][18] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][19]$_SDFFCE_PN0P_  (.D(_0652_),
    .DE(net130),
    .Q(\registers[25][19] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][1]$_SDFFCE_PN0P_  (.D(_0653_),
    .DE(net130),
    .Q(\registers[25][1] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][20]$_SDFFCE_PN0P_  (.D(_0654_),
    .DE(net130),
    .Q(\registers[25][20] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][21]$_SDFFCE_PN0P_  (.D(_0655_),
    .DE(net130),
    .Q(\registers[25][21] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][22]$_SDFFCE_PN0P_  (.D(_0656_),
    .DE(net130),
    .Q(\registers[25][22] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][23]$_SDFFCE_PN0P_  (.D(_0657_),
    .DE(_0014_),
    .Q(\registers[25][23] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][24]$_SDFFCE_PN0P_  (.D(_0658_),
    .DE(net130),
    .Q(\registers[25][24] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][25]$_SDFFCE_PN0P_  (.D(_0659_),
    .DE(net130),
    .Q(\registers[25][25] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][26]$_SDFFCE_PN0P_  (.D(_0660_),
    .DE(_0014_),
    .Q(\registers[25][26] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][27]$_SDFFCE_PN0P_  (.D(_0661_),
    .DE(net130),
    .Q(\registers[25][27] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][28]$_SDFFCE_PN0P_  (.D(_0662_),
    .DE(net130),
    .Q(\registers[25][28] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][29]$_SDFFCE_PN0P_  (.D(_0663_),
    .DE(net130),
    .Q(\registers[25][29] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][2]$_SDFFCE_PN0P_  (.D(_0664_),
    .DE(_0014_),
    .Q(\registers[25][2] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][30]$_SDFFCE_PN0P_  (.D(_0665_),
    .DE(_0014_),
    .Q(\registers[25][30] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][31]$_SDFFCE_PN0P_  (.D(_0666_),
    .DE(_0014_),
    .Q(\registers[25][31] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][3]$_SDFFCE_PN0P_  (.D(_0667_),
    .DE(_0014_),
    .Q(\registers[25][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][4]$_SDFFCE_PN0P_  (.D(_0668_),
    .DE(_0014_),
    .Q(\registers[25][4] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][5]$_SDFFCE_PN0P_  (.D(_0669_),
    .DE(_0014_),
    .Q(\registers[25][5] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][6]$_SDFFCE_PN0P_  (.D(_0670_),
    .DE(_0014_),
    .Q(\registers[25][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][7]$_SDFFCE_PN0P_  (.D(_0671_),
    .DE(_0014_),
    .Q(\registers[25][7] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][8]$_SDFFCE_PN0P_  (.D(_0672_),
    .DE(_0014_),
    .Q(\registers[25][8] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[25][9]$_SDFFCE_PN0P_  (.D(_0673_),
    .DE(_0014_),
    .Q(\registers[25][9] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][0]$_SDFFCE_PN0P_  (.D(_0674_),
    .DE(_0013_),
    .Q(\registers[26][0] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][10]$_SDFFCE_PN0P_  (.D(_0675_),
    .DE(_0013_),
    .Q(\registers[26][10] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][11]$_SDFFCE_PN0P_  (.D(_0676_),
    .DE(_0013_),
    .Q(\registers[26][11] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][12]$_SDFFCE_PN0P_  (.D(_0677_),
    .DE(_0013_),
    .Q(\registers[26][12] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][13]$_SDFFCE_PN0P_  (.D(_0678_),
    .DE(_0013_),
    .Q(\registers[26][13] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][14]$_SDFFCE_PN0P_  (.D(_0679_),
    .DE(_0013_),
    .Q(\registers[26][14] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][15]$_SDFFCE_PN0P_  (.D(_0680_),
    .DE(_0013_),
    .Q(\registers[26][15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][16]$_SDFFCE_PN0P_  (.D(_0681_),
    .DE(_0013_),
    .Q(\registers[26][16] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][17]$_SDFFCE_PN0P_  (.D(_0682_),
    .DE(_0013_),
    .Q(\registers[26][17] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][18]$_SDFFCE_PN0P_  (.D(_0683_),
    .DE(_0013_),
    .Q(\registers[26][18] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][19]$_SDFFCE_PN0P_  (.D(_0684_),
    .DE(_0013_),
    .Q(\registers[26][19] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][1]$_SDFFCE_PN0P_  (.D(_0685_),
    .DE(_0013_),
    .Q(\registers[26][1] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][20]$_SDFFCE_PN0P_  (.D(_0686_),
    .DE(_0013_),
    .Q(\registers[26][20] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][21]$_SDFFCE_PN0P_  (.D(_0687_),
    .DE(_0013_),
    .Q(\registers[26][21] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][22]$_SDFFCE_PN0P_  (.D(_0688_),
    .DE(_0013_),
    .Q(\registers[26][22] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][23]$_SDFFCE_PN0P_  (.D(_0689_),
    .DE(net129),
    .Q(\registers[26][23] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][24]$_SDFFCE_PN0P_  (.D(_0690_),
    .DE(net129),
    .Q(\registers[26][24] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][25]$_SDFFCE_PN0P_  (.D(_0691_),
    .DE(net129),
    .Q(\registers[26][25] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][26]$_SDFFCE_PN0P_  (.D(_0692_),
    .DE(net129),
    .Q(\registers[26][26] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][27]$_SDFFCE_PN0P_  (.D(_0693_),
    .DE(net129),
    .Q(\registers[26][27] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][28]$_SDFFCE_PN0P_  (.D(_0694_),
    .DE(net129),
    .Q(\registers[26][28] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][29]$_SDFFCE_PN0P_  (.D(_0695_),
    .DE(net129),
    .Q(\registers[26][29] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][2]$_SDFFCE_PN0P_  (.D(_0696_),
    .DE(net129),
    .Q(\registers[26][2] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][30]$_SDFFCE_PN0P_  (.D(_0697_),
    .DE(net129),
    .Q(\registers[26][30] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][31]$_SDFFCE_PN0P_  (.D(_0698_),
    .DE(net129),
    .Q(\registers[26][31] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][3]$_SDFFCE_PN0P_  (.D(_0699_),
    .DE(net129),
    .Q(\registers[26][3] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][4]$_SDFFCE_PN0P_  (.D(_0700_),
    .DE(net129),
    .Q(\registers[26][4] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][5]$_SDFFCE_PN0P_  (.D(_0701_),
    .DE(net129),
    .Q(\registers[26][5] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][6]$_SDFFCE_PN0P_  (.D(_0702_),
    .DE(net129),
    .Q(\registers[26][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][7]$_SDFFCE_PN0P_  (.D(_0703_),
    .DE(net129),
    .Q(\registers[26][7] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][8]$_SDFFCE_PN0P_  (.D(_0704_),
    .DE(net129),
    .Q(\registers[26][8] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[26][9]$_SDFFCE_PN0P_  (.D(_0705_),
    .DE(net129),
    .Q(\registers[26][9] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][0]$_SDFFCE_PN0P_  (.D(_0706_),
    .DE(net118),
    .Q(\registers[27][0] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][10]$_SDFFCE_PN0P_  (.D(_0707_),
    .DE(_0012_),
    .Q(\registers[27][10] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][11]$_SDFFCE_PN0P_  (.D(_0708_),
    .DE(_0012_),
    .Q(\registers[27][11] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][12]$_SDFFCE_PN0P_  (.D(_0709_),
    .DE(net118),
    .Q(\registers[27][12] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][13]$_SDFFCE_PN0P_  (.D(_0710_),
    .DE(_0012_),
    .Q(\registers[27][13] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][14]$_SDFFCE_PN0P_  (.D(_0711_),
    .DE(net118),
    .Q(\registers[27][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][15]$_SDFFCE_PN0P_  (.D(_0712_),
    .DE(_0012_),
    .Q(\registers[27][15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][16]$_SDFFCE_PN0P_  (.D(_0713_),
    .DE(_0012_),
    .Q(\registers[27][16] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][17]$_SDFFCE_PN0P_  (.D(_0714_),
    .DE(_0012_),
    .Q(\registers[27][17] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][18]$_SDFFCE_PN0P_  (.D(_0715_),
    .DE(_0012_),
    .Q(\registers[27][18] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][19]$_SDFFCE_PN0P_  (.D(_0716_),
    .DE(net118),
    .Q(\registers[27][19] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][1]$_SDFFCE_PN0P_  (.D(_0717_),
    .DE(net118),
    .Q(\registers[27][1] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][20]$_SDFFCE_PN0P_  (.D(_0718_),
    .DE(net118),
    .Q(\registers[27][20] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][21]$_SDFFCE_PN0P_  (.D(_0719_),
    .DE(net118),
    .Q(\registers[27][21] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][22]$_SDFFCE_PN0P_  (.D(_0720_),
    .DE(net118),
    .Q(\registers[27][22] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][23]$_SDFFCE_PN0P_  (.D(_0721_),
    .DE(net119),
    .Q(\registers[27][23] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][24]$_SDFFCE_PN0P_  (.D(_0722_),
    .DE(net118),
    .Q(\registers[27][24] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][25]$_SDFFCE_PN0P_  (.D(_0723_),
    .DE(net118),
    .Q(\registers[27][25] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][26]$_SDFFCE_PN0P_  (.D(_0724_),
    .DE(net119),
    .Q(\registers[27][26] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][27]$_SDFFCE_PN0P_  (.D(_0725_),
    .DE(net118),
    .Q(\registers[27][27] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][28]$_SDFFCE_PN0P_  (.D(_0726_),
    .DE(net118),
    .Q(\registers[27][28] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][29]$_SDFFCE_PN0P_  (.D(_0727_),
    .DE(net118),
    .Q(\registers[27][29] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][2]$_SDFFCE_PN0P_  (.D(_0728_),
    .DE(net119),
    .Q(\registers[27][2] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][30]$_SDFFCE_PN0P_  (.D(_0729_),
    .DE(net119),
    .Q(\registers[27][30] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][31]$_SDFFCE_PN0P_  (.D(_0730_),
    .DE(net119),
    .Q(\registers[27][31] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][3]$_SDFFCE_PN0P_  (.D(_0731_),
    .DE(net119),
    .Q(\registers[27][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][4]$_SDFFCE_PN0P_  (.D(_0732_),
    .DE(net119),
    .Q(\registers[27][4] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][5]$_SDFFCE_PN0P_  (.D(_0733_),
    .DE(net119),
    .Q(\registers[27][5] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][6]$_SDFFCE_PN0P_  (.D(_0734_),
    .DE(net119),
    .Q(\registers[27][6] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][7]$_SDFFCE_PN0P_  (.D(_0735_),
    .DE(net119),
    .Q(\registers[27][7] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][8]$_SDFFCE_PN0P_  (.D(_0736_),
    .DE(net119),
    .Q(\registers[27][8] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[27][9]$_SDFFCE_PN0P_  (.D(_0737_),
    .DE(net119),
    .Q(\registers[27][9] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][0]$_SDFFCE_PN0P_  (.D(_0738_),
    .DE(_0011_),
    .Q(\registers[28][0] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][10]$_SDFFCE_PN0P_  (.D(_0739_),
    .DE(_0011_),
    .Q(\registers[28][10] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][11]$_SDFFCE_PN0P_  (.D(_0740_),
    .DE(_0011_),
    .Q(\registers[28][11] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][12]$_SDFFCE_PN0P_  (.D(_0741_),
    .DE(_0011_),
    .Q(\registers[28][12] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][13]$_SDFFCE_PN0P_  (.D(_0742_),
    .DE(_0011_),
    .Q(\registers[28][13] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][14]$_SDFFCE_PN0P_  (.D(_0743_),
    .DE(_0011_),
    .Q(\registers[28][14] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][15]$_SDFFCE_PN0P_  (.D(_0744_),
    .DE(_0011_),
    .Q(\registers[28][15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][16]$_SDFFCE_PN0P_  (.D(_0745_),
    .DE(_0011_),
    .Q(\registers[28][16] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][17]$_SDFFCE_PN0P_  (.D(_0746_),
    .DE(_0011_),
    .Q(\registers[28][17] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][18]$_SDFFCE_PN0P_  (.D(_0747_),
    .DE(_0011_),
    .Q(\registers[28][18] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][19]$_SDFFCE_PN0P_  (.D(_0748_),
    .DE(_0011_),
    .Q(\registers[28][19] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][1]$_SDFFCE_PN0P_  (.D(_0749_),
    .DE(_0011_),
    .Q(\registers[28][1] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][20]$_SDFFCE_PN0P_  (.D(_0750_),
    .DE(net169),
    .Q(\registers[28][20] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][21]$_SDFFCE_PN0P_  (.D(_0751_),
    .DE(_0011_),
    .Q(\registers[28][21] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][22]$_SDFFCE_PN0P_  (.D(_0752_),
    .DE(net169),
    .Q(\registers[28][22] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][23]$_SDFFCE_PN0P_  (.D(_0753_),
    .DE(net169),
    .Q(\registers[28][23] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][24]$_SDFFCE_PN0P_  (.D(_0754_),
    .DE(net169),
    .Q(\registers[28][24] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][25]$_SDFFCE_PN0P_  (.D(_0755_),
    .DE(net169),
    .Q(\registers[28][25] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][26]$_SDFFCE_PN0P_  (.D(_0756_),
    .DE(net169),
    .Q(\registers[28][26] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][27]$_SDFFCE_PN0P_  (.D(_0757_),
    .DE(net169),
    .Q(\registers[28][27] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][28]$_SDFFCE_PN0P_  (.D(_0758_),
    .DE(net169),
    .Q(\registers[28][28] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][29]$_SDFFCE_PN0P_  (.D(_0759_),
    .DE(net169),
    .Q(\registers[28][29] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][2]$_SDFFCE_PN0P_  (.D(_0760_),
    .DE(net169),
    .Q(\registers[28][2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][30]$_SDFFCE_PN0P_  (.D(_0761_),
    .DE(net169),
    .Q(\registers[28][30] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][31]$_SDFFCE_PN0P_  (.D(_0762_),
    .DE(net169),
    .Q(\registers[28][31] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][3]$_SDFFCE_PN0P_  (.D(_0763_),
    .DE(net169),
    .Q(\registers[28][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][4]$_SDFFCE_PN0P_  (.D(_0764_),
    .DE(net169),
    .Q(\registers[28][4] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][5]$_SDFFCE_PN0P_  (.D(_0765_),
    .DE(net169),
    .Q(\registers[28][5] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][6]$_SDFFCE_PN0P_  (.D(_0766_),
    .DE(net169),
    .Q(\registers[28][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][7]$_SDFFCE_PN0P_  (.D(_0767_),
    .DE(net169),
    .Q(\registers[28][7] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][8]$_SDFFCE_PN0P_  (.D(_0768_),
    .DE(net169),
    .Q(\registers[28][8] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[28][9]$_SDFFCE_PN0P_  (.D(_0769_),
    .DE(net169),
    .Q(\registers[28][9] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][0]$_SDFFCE_PN0P_  (.D(_0770_),
    .DE(net128),
    .Q(\registers[29][0] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][10]$_SDFFCE_PN0P_  (.D(_0771_),
    .DE(net128),
    .Q(\registers[29][10] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][11]$_SDFFCE_PN0P_  (.D(_0772_),
    .DE(net128),
    .Q(\registers[29][11] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][12]$_SDFFCE_PN0P_  (.D(_0773_),
    .DE(net128),
    .Q(\registers[29][12] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][13]$_SDFFCE_PN0P_  (.D(_0774_),
    .DE(net128),
    .Q(\registers[29][13] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][14]$_SDFFCE_PN0P_  (.D(_0775_),
    .DE(net128),
    .Q(\registers[29][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][15]$_SDFFCE_PN0P_  (.D(_0776_),
    .DE(net128),
    .Q(\registers[29][15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][16]$_SDFFCE_PN0P_  (.D(_0777_),
    .DE(net128),
    .Q(\registers[29][16] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][17]$_SDFFCE_PN0P_  (.D(_0778_),
    .DE(net128),
    .Q(\registers[29][17] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][18]$_SDFFCE_PN0P_  (.D(_0779_),
    .DE(net128),
    .Q(\registers[29][18] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][19]$_SDFFCE_PN0P_  (.D(_0780_),
    .DE(net128),
    .Q(\registers[29][19] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][1]$_SDFFCE_PN0P_  (.D(_0781_),
    .DE(net128),
    .Q(\registers[29][1] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][20]$_SDFFCE_PN0P_  (.D(_0782_),
    .DE(net128),
    .Q(\registers[29][20] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][21]$_SDFFCE_PN0P_  (.D(_0783_),
    .DE(net128),
    .Q(\registers[29][21] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][22]$_SDFFCE_PN0P_  (.D(_0784_),
    .DE(net128),
    .Q(\registers[29][22] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][23]$_SDFFCE_PN0P_  (.D(_0785_),
    .DE(_0010_),
    .Q(\registers[29][23] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][24]$_SDFFCE_PN0P_  (.D(_0786_),
    .DE(net128),
    .Q(\registers[29][24] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][25]$_SDFFCE_PN0P_  (.D(_0787_),
    .DE(net128),
    .Q(\registers[29][25] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][26]$_SDFFCE_PN0P_  (.D(_0788_),
    .DE(_0010_),
    .Q(\registers[29][26] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][27]$_SDFFCE_PN0P_  (.D(_0789_),
    .DE(net128),
    .Q(\registers[29][27] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][28]$_SDFFCE_PN0P_  (.D(_0790_),
    .DE(net128),
    .Q(\registers[29][28] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][29]$_SDFFCE_PN0P_  (.D(_0791_),
    .DE(net128),
    .Q(\registers[29][29] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][2]$_SDFFCE_PN0P_  (.D(_0792_),
    .DE(_0010_),
    .Q(\registers[29][2] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][30]$_SDFFCE_PN0P_  (.D(_0793_),
    .DE(_0010_),
    .Q(\registers[29][30] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][31]$_SDFFCE_PN0P_  (.D(_0794_),
    .DE(_0010_),
    .Q(\registers[29][31] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][3]$_SDFFCE_PN0P_  (.D(_0795_),
    .DE(_0010_),
    .Q(\registers[29][3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][4]$_SDFFCE_PN0P_  (.D(_0796_),
    .DE(_0010_),
    .Q(\registers[29][4] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][5]$_SDFFCE_PN0P_  (.D(_0797_),
    .DE(_0010_),
    .Q(\registers[29][5] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][6]$_SDFFCE_PN0P_  (.D(_0798_),
    .DE(_0010_),
    .Q(\registers[29][6] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][7]$_SDFFCE_PN0P_  (.D(_0799_),
    .DE(_0010_),
    .Q(\registers[29][7] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][8]$_SDFFCE_PN0P_  (.D(_0800_),
    .DE(_0010_),
    .Q(\registers[29][8] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[29][9]$_SDFFCE_PN0P_  (.D(_0801_),
    .DE(_0010_),
    .Q(\registers[29][9] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][0]$_SDFFCE_PN0P_  (.D(_0802_),
    .DE(_0009_),
    .Q(\registers[2][0] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][10]$_SDFFCE_PN0P_  (.D(_0803_),
    .DE(_0009_),
    .Q(\registers[2][10] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][11]$_SDFFCE_PN0P_  (.D(_0804_),
    .DE(_0009_),
    .Q(\registers[2][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][12]$_SDFFCE_PN0P_  (.D(_0805_),
    .DE(_0009_),
    .Q(\registers[2][12] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][13]$_SDFFCE_PN0P_  (.D(_0806_),
    .DE(_0009_),
    .Q(\registers[2][13] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][14]$_SDFFCE_PN0P_  (.D(_0807_),
    .DE(_0009_),
    .Q(\registers[2][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][15]$_SDFFCE_PN0P_  (.D(_0808_),
    .DE(_0009_),
    .Q(\registers[2][15] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][16]$_SDFFCE_PN0P_  (.D(_0809_),
    .DE(_0009_),
    .Q(\registers[2][16] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][17]$_SDFFCE_PN0P_  (.D(_0810_),
    .DE(_0009_),
    .Q(\registers[2][17] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][18]$_SDFFCE_PN0P_  (.D(_0811_),
    .DE(_0009_),
    .Q(\registers[2][18] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][19]$_SDFFCE_PN0P_  (.D(_0812_),
    .DE(_0009_),
    .Q(\registers[2][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][1]$_SDFFCE_PN0P_  (.D(_0813_),
    .DE(_0009_),
    .Q(\registers[2][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][20]$_SDFFCE_PN0P_  (.D(_0814_),
    .DE(net127),
    .Q(\registers[2][20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][21]$_SDFFCE_PN0P_  (.D(_0815_),
    .DE(net127),
    .Q(\registers[2][21] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][22]$_SDFFCE_PN0P_  (.D(_0816_),
    .DE(net127),
    .Q(\registers[2][22] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][23]$_SDFFCE_PN0P_  (.D(_0817_),
    .DE(net127),
    .Q(\registers[2][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][24]$_SDFFCE_PN0P_  (.D(_0818_),
    .DE(net127),
    .Q(\registers[2][24] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][25]$_SDFFCE_PN0P_  (.D(_0819_),
    .DE(net127),
    .Q(\registers[2][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][26]$_SDFFCE_PN0P_  (.D(_0820_),
    .DE(net127),
    .Q(\registers[2][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][27]$_SDFFCE_PN0P_  (.D(_0821_),
    .DE(net127),
    .Q(\registers[2][27] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][28]$_SDFFCE_PN0P_  (.D(_0822_),
    .DE(net127),
    .Q(\registers[2][28] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][29]$_SDFFCE_PN0P_  (.D(_0823_),
    .DE(net127),
    .Q(\registers[2][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][2]$_SDFFCE_PN0P_  (.D(_0824_),
    .DE(net127),
    .Q(\registers[2][2] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][30]$_SDFFCE_PN0P_  (.D(_0825_),
    .DE(net127),
    .Q(\registers[2][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][31]$_SDFFCE_PN0P_  (.D(_0826_),
    .DE(net127),
    .Q(\registers[2][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][3]$_SDFFCE_PN0P_  (.D(_0827_),
    .DE(net127),
    .Q(\registers[2][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][4]$_SDFFCE_PN0P_  (.D(_0828_),
    .DE(net127),
    .Q(\registers[2][4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][5]$_SDFFCE_PN0P_  (.D(_0829_),
    .DE(net127),
    .Q(\registers[2][5] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][6]$_SDFFCE_PN0P_  (.D(_0830_),
    .DE(net127),
    .Q(\registers[2][6] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][7]$_SDFFCE_PN0P_  (.D(_0831_),
    .DE(net127),
    .Q(\registers[2][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][8]$_SDFFCE_PN0P_  (.D(_0832_),
    .DE(net127),
    .Q(\registers[2][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[2][9]$_SDFFCE_PN0P_  (.D(_0833_),
    .DE(net127),
    .Q(\registers[2][9] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][0]$_SDFFCE_PN0P_  (.D(_0834_),
    .DE(_0008_),
    .Q(\registers[30][0] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][10]$_SDFFCE_PN0P_  (.D(_0835_),
    .DE(_0008_),
    .Q(\registers[30][10] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][11]$_SDFFCE_PN0P_  (.D(_0836_),
    .DE(_0008_),
    .Q(\registers[30][11] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][12]$_SDFFCE_PN0P_  (.D(_0837_),
    .DE(_0008_),
    .Q(\registers[30][12] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][13]$_SDFFCE_PN0P_  (.D(_0838_),
    .DE(_0008_),
    .Q(\registers[30][13] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][14]$_SDFFCE_PN0P_  (.D(_0839_),
    .DE(_0008_),
    .Q(\registers[30][14] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][15]$_SDFFCE_PN0P_  (.D(_0840_),
    .DE(_0008_),
    .Q(\registers[30][15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][16]$_SDFFCE_PN0P_  (.D(_0841_),
    .DE(_0008_),
    .Q(\registers[30][16] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][17]$_SDFFCE_PN0P_  (.D(_0842_),
    .DE(_0008_),
    .Q(\registers[30][17] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][18]$_SDFFCE_PN0P_  (.D(_0843_),
    .DE(_0008_),
    .Q(\registers[30][18] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][19]$_SDFFCE_PN0P_  (.D(_0844_),
    .DE(_0008_),
    .Q(\registers[30][19] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][1]$_SDFFCE_PN0P_  (.D(_0845_),
    .DE(_0008_),
    .Q(\registers[30][1] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][20]$_SDFFCE_PN0P_  (.D(_0846_),
    .DE(_0008_),
    .Q(\registers[30][20] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][21]$_SDFFCE_PN0P_  (.D(_0847_),
    .DE(_0008_),
    .Q(\registers[30][21] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][22]$_SDFFCE_PN0P_  (.D(_0848_),
    .DE(_0008_),
    .Q(\registers[30][22] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][23]$_SDFFCE_PN0P_  (.D(_0849_),
    .DE(_0008_),
    .Q(\registers[30][23] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][24]$_SDFFCE_PN0P_  (.D(_0850_),
    .DE(_0008_),
    .Q(\registers[30][24] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][25]$_SDFFCE_PN0P_  (.D(_0851_),
    .DE(_0008_),
    .Q(\registers[30][25] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][26]$_SDFFCE_PN0P_  (.D(_0852_),
    .DE(_0008_),
    .Q(\registers[30][26] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][27]$_SDFFCE_PN0P_  (.D(_0853_),
    .DE(_0008_),
    .Q(\registers[30][27] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][28]$_SDFFCE_PN0P_  (.D(_0854_),
    .DE(_0008_),
    .Q(\registers[30][28] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][29]$_SDFFCE_PN0P_  (.D(_0855_),
    .DE(_0008_),
    .Q(\registers[30][29] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][2]$_SDFFCE_PN0P_  (.D(_0856_),
    .DE(_0008_),
    .Q(\registers[30][2] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][30]$_SDFFCE_PN0P_  (.D(_0857_),
    .DE(_0008_),
    .Q(\registers[30][30] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][31]$_SDFFCE_PN0P_  (.D(_0858_),
    .DE(_0008_),
    .Q(\registers[30][31] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][3]$_SDFFCE_PN0P_  (.D(_0859_),
    .DE(_0008_),
    .Q(\registers[30][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][4]$_SDFFCE_PN0P_  (.D(_0860_),
    .DE(_0008_),
    .Q(\registers[30][4] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][5]$_SDFFCE_PN0P_  (.D(_0861_),
    .DE(_0008_),
    .Q(\registers[30][5] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][6]$_SDFFCE_PN0P_  (.D(_0862_),
    .DE(_0008_),
    .Q(\registers[30][6] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][7]$_SDFFCE_PN0P_  (.D(_0863_),
    .DE(_0008_),
    .Q(\registers[30][7] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][8]$_SDFFCE_PN0P_  (.D(_0864_),
    .DE(_0008_),
    .Q(\registers[30][8] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[30][9]$_SDFFCE_PN0P_  (.D(_0865_),
    .DE(_0008_),
    .Q(\registers[30][9] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][0]$_SDFFCE_PN0P_  (.D(_0866_),
    .DE(net117),
    .Q(\registers[31][0] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][10]$_SDFFCE_PN0P_  (.D(_0867_),
    .DE(_0007_),
    .Q(\registers[31][10] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][11]$_SDFFCE_PN0P_  (.D(_0868_),
    .DE(_0007_),
    .Q(\registers[31][11] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][12]$_SDFFCE_PN0P_  (.D(_0869_),
    .DE(net117),
    .Q(\registers[31][12] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][13]$_SDFFCE_PN0P_  (.D(_0870_),
    .DE(_0007_),
    .Q(\registers[31][13] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][14]$_SDFFCE_PN0P_  (.D(_0871_),
    .DE(net117),
    .Q(\registers[31][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][15]$_SDFFCE_PN0P_  (.D(_0872_),
    .DE(_0007_),
    .Q(\registers[31][15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][16]$_SDFFCE_PN0P_  (.D(_0873_),
    .DE(_0007_),
    .Q(\registers[31][16] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][17]$_SDFFCE_PN0P_  (.D(_0874_),
    .DE(_0007_),
    .Q(\registers[31][17] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][18]$_SDFFCE_PN0P_  (.D(_0875_),
    .DE(_0007_),
    .Q(\registers[31][18] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][19]$_SDFFCE_PN0P_  (.D(_0876_),
    .DE(net117),
    .Q(\registers[31][19] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][1]$_SDFFCE_PN0P_  (.D(_0877_),
    .DE(_0007_),
    .Q(\registers[31][1] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][20]$_SDFFCE_PN0P_  (.D(_0878_),
    .DE(net117),
    .Q(\registers[31][20] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][21]$_SDFFCE_PN0P_  (.D(_0879_),
    .DE(net117),
    .Q(\registers[31][21] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][22]$_SDFFCE_PN0P_  (.D(_0880_),
    .DE(net117),
    .Q(\registers[31][22] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][23]$_SDFFCE_PN0P_  (.D(_0881_),
    .DE(net116),
    .Q(\registers[31][23] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][24]$_SDFFCE_PN0P_  (.D(_0882_),
    .DE(net117),
    .Q(\registers[31][24] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][25]$_SDFFCE_PN0P_  (.D(_0883_),
    .DE(net117),
    .Q(\registers[31][25] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][26]$_SDFFCE_PN0P_  (.D(_0884_),
    .DE(net116),
    .Q(\registers[31][26] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][27]$_SDFFCE_PN0P_  (.D(_0885_),
    .DE(net117),
    .Q(\registers[31][27] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][28]$_SDFFCE_PN0P_  (.D(_0886_),
    .DE(net117),
    .Q(\registers[31][28] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][29]$_SDFFCE_PN0P_  (.D(_0887_),
    .DE(net117),
    .Q(\registers[31][29] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][2]$_SDFFCE_PN0P_  (.D(_0888_),
    .DE(net116),
    .Q(\registers[31][2] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][30]$_SDFFCE_PN0P_  (.D(_0889_),
    .DE(net116),
    .Q(\registers[31][30] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][31]$_SDFFCE_PN0P_  (.D(_0890_),
    .DE(net116),
    .Q(\registers[31][31] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][3]$_SDFFCE_PN0P_  (.D(_0891_),
    .DE(net116),
    .Q(\registers[31][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][4]$_SDFFCE_PN0P_  (.D(_0892_),
    .DE(net116),
    .Q(\registers[31][4] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][5]$_SDFFCE_PN0P_  (.D(_0893_),
    .DE(net116),
    .Q(\registers[31][5] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][6]$_SDFFCE_PN0P_  (.D(_0894_),
    .DE(net116),
    .Q(\registers[31][6] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][7]$_SDFFCE_PN0P_  (.D(_0895_),
    .DE(net116),
    .Q(\registers[31][7] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][8]$_SDFFCE_PN0P_  (.D(_0896_),
    .DE(net116),
    .Q(\registers[31][8] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[31][9]$_SDFFCE_PN0P_  (.D(_0897_),
    .DE(net116),
    .Q(\registers[31][9] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][0]$_SDFFCE_PN0P_  (.D(_0898_),
    .DE(_0006_),
    .Q(\registers[3][0] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][10]$_SDFFCE_PN0P_  (.D(_0899_),
    .DE(_0006_),
    .Q(\registers[3][10] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][11]$_SDFFCE_PN0P_  (.D(_0900_),
    .DE(_0006_),
    .Q(\registers[3][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][12]$_SDFFCE_PN0P_  (.D(_0901_),
    .DE(_0006_),
    .Q(\registers[3][12] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][13]$_SDFFCE_PN0P_  (.D(_0902_),
    .DE(_0006_),
    .Q(\registers[3][13] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][14]$_SDFFCE_PN0P_  (.D(_0903_),
    .DE(_0006_),
    .Q(\registers[3][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][15]$_SDFFCE_PN0P_  (.D(_0904_),
    .DE(_0006_),
    .Q(\registers[3][15] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][16]$_SDFFCE_PN0P_  (.D(_0905_),
    .DE(_0006_),
    .Q(\registers[3][16] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][17]$_SDFFCE_PN0P_  (.D(_0906_),
    .DE(net115),
    .Q(\registers[3][17] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][18]$_SDFFCE_PN0P_  (.D(_0907_),
    .DE(_0006_),
    .Q(\registers[3][18] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][19]$_SDFFCE_PN0P_  (.D(_0908_),
    .DE(net115),
    .Q(\registers[3][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][1]$_SDFFCE_PN0P_  (.D(_0909_),
    .DE(net115),
    .Q(\registers[3][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][20]$_SDFFCE_PN0P_  (.D(_0910_),
    .DE(net115),
    .Q(\registers[3][20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][21]$_SDFFCE_PN0P_  (.D(_0911_),
    .DE(net115),
    .Q(\registers[3][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][22]$_SDFFCE_PN0P_  (.D(_0912_),
    .DE(net115),
    .Q(\registers[3][22] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][23]$_SDFFCE_PN0P_  (.D(_0913_),
    .DE(net115),
    .Q(\registers[3][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][24]$_SDFFCE_PN0P_  (.D(_0914_),
    .DE(net115),
    .Q(\registers[3][24] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][25]$_SDFFCE_PN0P_  (.D(_0915_),
    .DE(net115),
    .Q(\registers[3][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][26]$_SDFFCE_PN0P_  (.D(_0916_),
    .DE(net115),
    .Q(\registers[3][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][27]$_SDFFCE_PN0P_  (.D(_0917_),
    .DE(net115),
    .Q(\registers[3][27] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][28]$_SDFFCE_PN0P_  (.D(_0918_),
    .DE(net115),
    .Q(\registers[3][28] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][29]$_SDFFCE_PN0P_  (.D(_0919_),
    .DE(net115),
    .Q(\registers[3][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][2]$_SDFFCE_PN0P_  (.D(_0920_),
    .DE(net115),
    .Q(\registers[3][2] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][30]$_SDFFCE_PN0P_  (.D(_0921_),
    .DE(net115),
    .Q(\registers[3][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][31]$_SDFFCE_PN0P_  (.D(_0922_),
    .DE(_0006_),
    .Q(\registers[3][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][3]$_SDFFCE_PN0P_  (.D(_0923_),
    .DE(_0006_),
    .Q(\registers[3][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][4]$_SDFFCE_PN0P_  (.D(_0924_),
    .DE(_0006_),
    .Q(\registers[3][4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][5]$_SDFFCE_PN0P_  (.D(_0925_),
    .DE(_0006_),
    .Q(\registers[3][5] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][6]$_SDFFCE_PN0P_  (.D(_0926_),
    .DE(_0006_),
    .Q(\registers[3][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][7]$_SDFFCE_PN0P_  (.D(_0927_),
    .DE(_0006_),
    .Q(\registers[3][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][8]$_SDFFCE_PN0P_  (.D(_0928_),
    .DE(_0006_),
    .Q(\registers[3][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[3][9]$_SDFFCE_PN0P_  (.D(_0929_),
    .DE(net115),
    .Q(\registers[3][9] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][0]$_SDFFCE_PN0P_  (.D(_0930_),
    .DE(_0005_),
    .Q(\registers[4][0] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][10]$_SDFFCE_PN0P_  (.D(_0931_),
    .DE(_0005_),
    .Q(\registers[4][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][11]$_SDFFCE_PN0P_  (.D(_0932_),
    .DE(_0005_),
    .Q(\registers[4][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][12]$_SDFFCE_PN0P_  (.D(_0933_),
    .DE(_0005_),
    .Q(\registers[4][12] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][13]$_SDFFCE_PN0P_  (.D(_0934_),
    .DE(_0005_),
    .Q(\registers[4][13] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][14]$_SDFFCE_PN0P_  (.D(_0935_),
    .DE(_0005_),
    .Q(\registers[4][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][15]$_SDFFCE_PN0P_  (.D(_0936_),
    .DE(_0005_),
    .Q(\registers[4][15] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][16]$_SDFFCE_PN0P_  (.D(_0937_),
    .DE(_0005_),
    .Q(\registers[4][16] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][17]$_SDFFCE_PN0P_  (.D(_0938_),
    .DE(net109),
    .Q(\registers[4][17] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][18]$_SDFFCE_PN0P_  (.D(_0939_),
    .DE(_0005_),
    .Q(\registers[4][18] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][19]$_SDFFCE_PN0P_  (.D(_0940_),
    .DE(net109),
    .Q(\registers[4][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][1]$_SDFFCE_PN0P_  (.D(_0941_),
    .DE(net109),
    .Q(\registers[4][1] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][20]$_SDFFCE_PN0P_  (.D(_0942_),
    .DE(net109),
    .Q(\registers[4][20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][21]$_SDFFCE_PN0P_  (.D(_0943_),
    .DE(net109),
    .Q(\registers[4][21] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][22]$_SDFFCE_PN0P_  (.D(_0944_),
    .DE(net109),
    .Q(\registers[4][22] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][23]$_SDFFCE_PN0P_  (.D(_0945_),
    .DE(net109),
    .Q(\registers[4][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][24]$_SDFFCE_PN0P_  (.D(_0946_),
    .DE(net109),
    .Q(\registers[4][24] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][25]$_SDFFCE_PN0P_  (.D(_0947_),
    .DE(net109),
    .Q(\registers[4][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][26]$_SDFFCE_PN0P_  (.D(_0948_),
    .DE(net110),
    .Q(\registers[4][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][27]$_SDFFCE_PN0P_  (.D(_0949_),
    .DE(net109),
    .Q(\registers[4][27] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][28]$_SDFFCE_PN0P_  (.D(_0950_),
    .DE(net110),
    .Q(\registers[4][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][29]$_SDFFCE_PN0P_  (.D(_0951_),
    .DE(net109),
    .Q(\registers[4][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][2]$_SDFFCE_PN0P_  (.D(_0952_),
    .DE(net109),
    .Q(\registers[4][2] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][30]$_SDFFCE_PN0P_  (.D(_0953_),
    .DE(net109),
    .Q(\registers[4][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][31]$_SDFFCE_PN0P_  (.D(_0954_),
    .DE(net110),
    .Q(\registers[4][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][3]$_SDFFCE_PN0P_  (.D(_0955_),
    .DE(net110),
    .Q(\registers[4][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][4]$_SDFFCE_PN0P_  (.D(_0956_),
    .DE(net110),
    .Q(\registers[4][4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][5]$_SDFFCE_PN0P_  (.D(_0957_),
    .DE(net110),
    .Q(\registers[4][5] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][6]$_SDFFCE_PN0P_  (.D(_0958_),
    .DE(net110),
    .Q(\registers[4][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][7]$_SDFFCE_PN0P_  (.D(_0959_),
    .DE(net110),
    .Q(\registers[4][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][8]$_SDFFCE_PN0P_  (.D(_0960_),
    .DE(net110),
    .Q(\registers[4][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[4][9]$_SDFFCE_PN0P_  (.D(_0961_),
    .DE(net110),
    .Q(\registers[4][9] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][0]$_SDFFCE_PN0P_  (.D(_0962_),
    .DE(_0004_),
    .Q(\registers[5][0] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][10]$_SDFFCE_PN0P_  (.D(_0963_),
    .DE(_0004_),
    .Q(\registers[5][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][11]$_SDFFCE_PN0P_  (.D(_0964_),
    .DE(_0004_),
    .Q(\registers[5][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][12]$_SDFFCE_PN0P_  (.D(_0965_),
    .DE(_0004_),
    .Q(\registers[5][12] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][13]$_SDFFCE_PN0P_  (.D(_0966_),
    .DE(_0004_),
    .Q(\registers[5][13] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][14]$_SDFFCE_PN0P_  (.D(_0967_),
    .DE(_0004_),
    .Q(\registers[5][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][15]$_SDFFCE_PN0P_  (.D(_0968_),
    .DE(_0004_),
    .Q(\registers[5][15] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][16]$_SDFFCE_PN0P_  (.D(_0969_),
    .DE(_0004_),
    .Q(\registers[5][16] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][17]$_SDFFCE_PN0P_  (.D(_0970_),
    .DE(net125),
    .Q(\registers[5][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][18]$_SDFFCE_PN0P_  (.D(_0971_),
    .DE(_0004_),
    .Q(\registers[5][18] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][19]$_SDFFCE_PN0P_  (.D(_0972_),
    .DE(net125),
    .Q(\registers[5][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][1]$_SDFFCE_PN0P_  (.D(_0973_),
    .DE(net125),
    .Q(\registers[5][1] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][20]$_SDFFCE_PN0P_  (.D(_0974_),
    .DE(net125),
    .Q(\registers[5][20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][21]$_SDFFCE_PN0P_  (.D(_0975_),
    .DE(net125),
    .Q(\registers[5][21] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][22]$_SDFFCE_PN0P_  (.D(_0976_),
    .DE(net125),
    .Q(\registers[5][22] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][23]$_SDFFCE_PN0P_  (.D(_0977_),
    .DE(net125),
    .Q(\registers[5][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][24]$_SDFFCE_PN0P_  (.D(_0978_),
    .DE(net125),
    .Q(\registers[5][24] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][25]$_SDFFCE_PN0P_  (.D(_0979_),
    .DE(net125),
    .Q(\registers[5][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][26]$_SDFFCE_PN0P_  (.D(_0980_),
    .DE(net126),
    .Q(\registers[5][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][27]$_SDFFCE_PN0P_  (.D(_0981_),
    .DE(net125),
    .Q(\registers[5][27] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][28]$_SDFFCE_PN0P_  (.D(_0982_),
    .DE(net126),
    .Q(\registers[5][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][29]$_SDFFCE_PN0P_  (.D(_0983_),
    .DE(net125),
    .Q(\registers[5][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][2]$_SDFFCE_PN0P_  (.D(_0984_),
    .DE(net125),
    .Q(\registers[5][2] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][30]$_SDFFCE_PN0P_  (.D(_0985_),
    .DE(net125),
    .Q(\registers[5][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][31]$_SDFFCE_PN0P_  (.D(_0986_),
    .DE(net126),
    .Q(\registers[5][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][3]$_SDFFCE_PN0P_  (.D(_0987_),
    .DE(net126),
    .Q(\registers[5][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][4]$_SDFFCE_PN0P_  (.D(_0988_),
    .DE(net126),
    .Q(\registers[5][4] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][5]$_SDFFCE_PN0P_  (.D(_0989_),
    .DE(net126),
    .Q(\registers[5][5] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][6]$_SDFFCE_PN0P_  (.D(_0990_),
    .DE(net126),
    .Q(\registers[5][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][7]$_SDFFCE_PN0P_  (.D(_0991_),
    .DE(net126),
    .Q(\registers[5][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][8]$_SDFFCE_PN0P_  (.D(_0992_),
    .DE(net126),
    .Q(\registers[5][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[5][9]$_SDFFCE_PN0P_  (.D(_0993_),
    .DE(net126),
    .Q(\registers[5][9] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][0]$_SDFFCE_PN0P_  (.D(_0994_),
    .DE(_0003_),
    .Q(\registers[6][0] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][10]$_SDFFCE_PN0P_  (.D(_0995_),
    .DE(_0003_),
    .Q(\registers[6][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][11]$_SDFFCE_PN0P_  (.D(_0996_),
    .DE(_0003_),
    .Q(\registers[6][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][12]$_SDFFCE_PN0P_  (.D(_0997_),
    .DE(_0003_),
    .Q(\registers[6][12] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][13]$_SDFFCE_PN0P_  (.D(_0998_),
    .DE(_0003_),
    .Q(\registers[6][13] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][14]$_SDFFCE_PN0P_  (.D(_0999_),
    .DE(_0003_),
    .Q(\registers[6][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][15]$_SDFFCE_PN0P_  (.D(_1000_),
    .DE(_0003_),
    .Q(\registers[6][15] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][16]$_SDFFCE_PN0P_  (.D(_1001_),
    .DE(_0003_),
    .Q(\registers[6][16] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][17]$_SDFFCE_PN0P_  (.D(_1002_),
    .DE(_0003_),
    .Q(\registers[6][17] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][18]$_SDFFCE_PN0P_  (.D(_1003_),
    .DE(_0003_),
    .Q(\registers[6][18] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][19]$_SDFFCE_PN0P_  (.D(_1004_),
    .DE(net123),
    .Q(\registers[6][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][1]$_SDFFCE_PN0P_  (.D(_1005_),
    .DE(net123),
    .Q(\registers[6][1] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][20]$_SDFFCE_PN0P_  (.D(_1006_),
    .DE(net123),
    .Q(\registers[6][20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][21]$_SDFFCE_PN0P_  (.D(_1007_),
    .DE(net123),
    .Q(\registers[6][21] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][22]$_SDFFCE_PN0P_  (.D(_1008_),
    .DE(net123),
    .Q(\registers[6][22] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][23]$_SDFFCE_PN0P_  (.D(_1009_),
    .DE(net123),
    .Q(\registers[6][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][24]$_SDFFCE_PN0P_  (.D(_1010_),
    .DE(net123),
    .Q(\registers[6][24] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][25]$_SDFFCE_PN0P_  (.D(_1011_),
    .DE(net123),
    .Q(\registers[6][25] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][26]$_SDFFCE_PN0P_  (.D(_1012_),
    .DE(net123),
    .Q(\registers[6][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][27]$_SDFFCE_PN0P_  (.D(_1013_),
    .DE(net123),
    .Q(\registers[6][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][28]$_SDFFCE_PN0P_  (.D(_1014_),
    .DE(net123),
    .Q(\registers[6][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][29]$_SDFFCE_PN0P_  (.D(_1015_),
    .DE(net123),
    .Q(\registers[6][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][2]$_SDFFCE_PN0P_  (.D(_1016_),
    .DE(net123),
    .Q(\registers[6][2] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][30]$_SDFFCE_PN0P_  (.D(_1017_),
    .DE(net123),
    .Q(\registers[6][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][31]$_SDFFCE_PN0P_  (.D(_1018_),
    .DE(net124),
    .Q(\registers[6][31] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][3]$_SDFFCE_PN0P_  (.D(_1019_),
    .DE(net124),
    .Q(\registers[6][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][4]$_SDFFCE_PN0P_  (.D(_1020_),
    .DE(net124),
    .Q(\registers[6][4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][5]$_SDFFCE_PN0P_  (.D(_1021_),
    .DE(net124),
    .Q(\registers[6][5] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][6]$_SDFFCE_PN0P_  (.D(_1022_),
    .DE(net124),
    .Q(\registers[6][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][7]$_SDFFCE_PN0P_  (.D(_1023_),
    .DE(net124),
    .Q(\registers[6][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][8]$_SDFFCE_PN0P_  (.D(_1024_),
    .DE(net124),
    .Q(\registers[6][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[6][9]$_SDFFCE_PN0P_  (.D(_1025_),
    .DE(net124),
    .Q(\registers[6][9] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][0]$_SDFFCE_PN0P_  (.D(_1026_),
    .DE(_0002_),
    .Q(\registers[7][0] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][10]$_SDFFCE_PN0P_  (.D(_1027_),
    .DE(_0002_),
    .Q(\registers[7][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][11]$_SDFFCE_PN0P_  (.D(_1028_),
    .DE(_0002_),
    .Q(\registers[7][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][12]$_SDFFCE_PN0P_  (.D(_1029_),
    .DE(_0002_),
    .Q(\registers[7][12] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][13]$_SDFFCE_PN0P_  (.D(_1030_),
    .DE(_0002_),
    .Q(\registers[7][13] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][14]$_SDFFCE_PN0P_  (.D(_1031_),
    .DE(_0002_),
    .Q(\registers[7][14] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][15]$_SDFFCE_PN0P_  (.D(_1032_),
    .DE(_0002_),
    .Q(\registers[7][15] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][16]$_SDFFCE_PN0P_  (.D(_1033_),
    .DE(_0002_),
    .Q(\registers[7][16] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][17]$_SDFFCE_PN0P_  (.D(_1034_),
    .DE(net114),
    .Q(\registers[7][17] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][18]$_SDFFCE_PN0P_  (.D(_1035_),
    .DE(_0002_),
    .Q(\registers[7][18] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][19]$_SDFFCE_PN0P_  (.D(_1036_),
    .DE(net114),
    .Q(\registers[7][19] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][1]$_SDFFCE_PN0P_  (.D(_1037_),
    .DE(net114),
    .Q(\registers[7][1] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][20]$_SDFFCE_PN0P_  (.D(_1038_),
    .DE(net114),
    .Q(\registers[7][20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][21]$_SDFFCE_PN0P_  (.D(_1039_),
    .DE(net114),
    .Q(\registers[7][21] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][22]$_SDFFCE_PN0P_  (.D(_1040_),
    .DE(net114),
    .Q(\registers[7][22] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][23]$_SDFFCE_PN0P_  (.D(_1041_),
    .DE(net114),
    .Q(\registers[7][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][24]$_SDFFCE_PN0P_  (.D(_1042_),
    .DE(net114),
    .Q(\registers[7][24] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][25]$_SDFFCE_PN0P_  (.D(_1043_),
    .DE(net114),
    .Q(\registers[7][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][26]$_SDFFCE_PN0P_  (.D(_1044_),
    .DE(net114),
    .Q(\registers[7][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][27]$_SDFFCE_PN0P_  (.D(_1045_),
    .DE(net114),
    .Q(\registers[7][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][28]$_SDFFCE_PN0P_  (.D(_1046_),
    .DE(net114),
    .Q(\registers[7][28] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][29]$_SDFFCE_PN0P_  (.D(_1047_),
    .DE(net114),
    .Q(\registers[7][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][2]$_SDFFCE_PN0P_  (.D(_1048_),
    .DE(net114),
    .Q(\registers[7][2] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][30]$_SDFFCE_PN0P_  (.D(_1049_),
    .DE(net114),
    .Q(\registers[7][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][31]$_SDFFCE_PN0P_  (.D(_1050_),
    .DE(_0002_),
    .Q(\registers[7][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][3]$_SDFFCE_PN0P_  (.D(_1051_),
    .DE(_0002_),
    .Q(\registers[7][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][4]$_SDFFCE_PN0P_  (.D(_1052_),
    .DE(_0002_),
    .Q(\registers[7][4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][5]$_SDFFCE_PN0P_  (.D(_1053_),
    .DE(_0002_),
    .Q(\registers[7][5] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][6]$_SDFFCE_PN0P_  (.D(_1054_),
    .DE(_0002_),
    .Q(\registers[7][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][7]$_SDFFCE_PN0P_  (.D(_1055_),
    .DE(_0002_),
    .Q(\registers[7][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][8]$_SDFFCE_PN0P_  (.D(_1056_),
    .DE(_0002_),
    .Q(\registers[7][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[7][9]$_SDFFCE_PN0P_  (.D(_1057_),
    .DE(_0002_),
    .Q(\registers[7][9] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][0]$_SDFFCE_PN0P_  (.D(_1058_),
    .DE(_0001_),
    .Q(\registers[8][0] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][10]$_SDFFCE_PN0P_  (.D(_1059_),
    .DE(_0001_),
    .Q(\registers[8][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][11]$_SDFFCE_PN0P_  (.D(_1060_),
    .DE(_0001_),
    .Q(\registers[8][11] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][12]$_SDFFCE_PN0P_  (.D(_1061_),
    .DE(_0001_),
    .Q(\registers[8][12] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][13]$_SDFFCE_PN0P_  (.D(_1062_),
    .DE(_0001_),
    .Q(\registers[8][13] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][14]$_SDFFCE_PN0P_  (.D(_1063_),
    .DE(_0001_),
    .Q(\registers[8][14] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][15]$_SDFFCE_PN0P_  (.D(_1064_),
    .DE(_0001_),
    .Q(\registers[8][15] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][16]$_SDFFCE_PN0P_  (.D(_1065_),
    .DE(_0001_),
    .Q(\registers[8][16] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][17]$_SDFFCE_PN0P_  (.D(_1066_),
    .DE(_0001_),
    .Q(\registers[8][17] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][18]$_SDFFCE_PN0P_  (.D(_1067_),
    .DE(_0001_),
    .Q(\registers[8][18] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][19]$_SDFFCE_PN0P_  (.D(_1068_),
    .DE(_0001_),
    .Q(\registers[8][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][1]$_SDFFCE_PN0P_  (.D(_1069_),
    .DE(_0001_),
    .Q(\registers[8][1] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][20]$_SDFFCE_PN0P_  (.D(_1070_),
    .DE(_0001_),
    .Q(\registers[8][20] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][21]$_SDFFCE_PN0P_  (.D(_1071_),
    .DE(_0001_),
    .Q(\registers[8][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][22]$_SDFFCE_PN0P_  (.D(_1072_),
    .DE(_0001_),
    .Q(\registers[8][22] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][23]$_SDFFCE_PN0P_  (.D(_1073_),
    .DE(_0001_),
    .Q(\registers[8][23] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][24]$_SDFFCE_PN0P_  (.D(_1074_),
    .DE(_0001_),
    .Q(\registers[8][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][25]$_SDFFCE_PN0P_  (.D(_1075_),
    .DE(net108),
    .Q(\registers[8][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][26]$_SDFFCE_PN0P_  (.D(_1076_),
    .DE(net108),
    .Q(\registers[8][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][27]$_SDFFCE_PN0P_  (.D(_1077_),
    .DE(net108),
    .Q(\registers[8][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][28]$_SDFFCE_PN0P_  (.D(_1078_),
    .DE(net108),
    .Q(\registers[8][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][29]$_SDFFCE_PN0P_  (.D(_1079_),
    .DE(net108),
    .Q(\registers[8][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][2]$_SDFFCE_PN0P_  (.D(_1080_),
    .DE(net108),
    .Q(\registers[8][2] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][30]$_SDFFCE_PN0P_  (.D(_1081_),
    .DE(net108),
    .Q(\registers[8][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][31]$_SDFFCE_PN0P_  (.D(_1082_),
    .DE(net108),
    .Q(\registers[8][31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][3]$_SDFFCE_PN0P_  (.D(_1083_),
    .DE(net108),
    .Q(\registers[8][3] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][4]$_SDFFCE_PN0P_  (.D(_1084_),
    .DE(net108),
    .Q(\registers[8][4] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][5]$_SDFFCE_PN0P_  (.D(_1085_),
    .DE(net108),
    .Q(\registers[8][5] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][6]$_SDFFCE_PN0P_  (.D(_1086_),
    .DE(net108),
    .Q(\registers[8][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][7]$_SDFFCE_PN0P_  (.D(_1087_),
    .DE(net108),
    .Q(\registers[8][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][8]$_SDFFCE_PN0P_  (.D(_1088_),
    .DE(net108),
    .Q(\registers[8][8] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[8][9]$_SDFFCE_PN0P_  (.D(_1089_),
    .DE(net108),
    .Q(\registers[8][9] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][0]$_SDFFCE_PN0P_  (.D(_1090_),
    .DE(_0000_),
    .Q(\registers[9][0] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][10]$_SDFFCE_PN0P_  (.D(_1091_),
    .DE(net122),
    .Q(\registers[9][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][11]$_SDFFCE_PN0P_  (.D(_1092_),
    .DE(net122),
    .Q(\registers[9][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][12]$_SDFFCE_PN0P_  (.D(_1093_),
    .DE(net122),
    .Q(\registers[9][12] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][13]$_SDFFCE_PN0P_  (.D(_1094_),
    .DE(net122),
    .Q(\registers[9][13] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][14]$_SDFFCE_PN0P_  (.D(_1095_),
    .DE(net122),
    .Q(\registers[9][14] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][15]$_SDFFCE_PN0P_  (.D(_1096_),
    .DE(net122),
    .Q(\registers[9][15] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][16]$_SDFFCE_PN0P_  (.D(_1097_),
    .DE(net122),
    .Q(\registers[9][16] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][17]$_SDFFCE_PN0P_  (.D(_1098_),
    .DE(net122),
    .Q(\registers[9][17] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][18]$_SDFFCE_PN0P_  (.D(_1099_),
    .DE(net122),
    .Q(\registers[9][18] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][19]$_SDFFCE_PN0P_  (.D(_1100_),
    .DE(net122),
    .Q(\registers[9][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][1]$_SDFFCE_PN0P_  (.D(_1101_),
    .DE(net122),
    .Q(\registers[9][1] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][20]$_SDFFCE_PN0P_  (.D(_1102_),
    .DE(net122),
    .Q(\registers[9][20] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][21]$_SDFFCE_PN0P_  (.D(_1103_),
    .DE(net122),
    .Q(\registers[9][21] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][22]$_SDFFCE_PN0P_  (.D(_1104_),
    .DE(net122),
    .Q(\registers[9][22] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][23]$_SDFFCE_PN0P_  (.D(_1105_),
    .DE(net122),
    .Q(\registers[9][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][24]$_SDFFCE_PN0P_  (.D(_1106_),
    .DE(net122),
    .Q(\registers[9][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][25]$_SDFFCE_PN0P_  (.D(_1107_),
    .DE(net122),
    .Q(\registers[9][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][26]$_SDFFCE_PN0P_  (.D(_1108_),
    .DE(net122),
    .Q(\registers[9][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][27]$_SDFFCE_PN0P_  (.D(_1109_),
    .DE(net122),
    .Q(\registers[9][27] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][28]$_SDFFCE_PN0P_  (.D(_1110_),
    .DE(net122),
    .Q(\registers[9][28] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][29]$_SDFFCE_PN0P_  (.D(_1111_),
    .DE(net122),
    .Q(\registers[9][29] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][2]$_SDFFCE_PN0P_  (.D(_1112_),
    .DE(net122),
    .Q(\registers[9][2] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][30]$_SDFFCE_PN0P_  (.D(_1113_),
    .DE(_0000_),
    .Q(\registers[9][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][31]$_SDFFCE_PN0P_  (.D(_1114_),
    .DE(_0000_),
    .Q(\registers[9][31] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][3]$_SDFFCE_PN0P_  (.D(_1115_),
    .DE(_0000_),
    .Q(\registers[9][3] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][4]$_SDFFCE_PN0P_  (.D(_1116_),
    .DE(_0000_),
    .Q(\registers[9][4] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][5]$_SDFFCE_PN0P_  (.D(_1117_),
    .DE(_0000_),
    .Q(\registers[9][5] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][6]$_SDFFCE_PN0P_  (.D(_1118_),
    .DE(_0000_),
    .Q(\registers[9][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][7]$_SDFFCE_PN0P_  (.D(_1119_),
    .DE(_0000_),
    .Q(\registers[9][7] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][8]$_SDFFCE_PN0P_  (.D(_1120_),
    .DE(_0000_),
    .Q(\registers[9][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \registers[9][9]$_SDFFCE_PN0P_  (.D(_1121_),
    .DE(_0000_),
    .Q(\registers[9][9] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1367 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(read_addr1[3]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(read_addr2[3]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(read_en1),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(read_en2),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(rst_n),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(write_addr[0]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(write_addr[1]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_8 input8 (.A(write_addr[2]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(write_addr[3]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(write_addr[4]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(net153),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(net152),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(net154),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(net165),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(net155),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(net147),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(net145),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(net158),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(net156),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(net164),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(net151),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(net140),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(net148),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(net137),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(net138),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(net135),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(net149),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(net139),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(net150),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(net142),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(net161),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(net136),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(net160),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(net143),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(net141),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(net163),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(net146),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(net144),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(net166),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input40 (.A(net162),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(net157),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(net159),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(write_en),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net44),
    .X(read_data1[0]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net45),
    .X(read_data1[10]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net46),
    .X(read_data1[11]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net47),
    .X(read_data1[12]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net48),
    .X(read_data1[13]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net49),
    .X(read_data1[14]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net50),
    .X(read_data1[15]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net51),
    .X(read_data1[16]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net52),
    .X(read_data1[17]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(read_data1[18]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(read_data1[19]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(read_data1[1]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(read_data1[20]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(read_data1[21]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(read_data1[22]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(read_data1[23]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(read_data1[24]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(read_data1[25]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(read_data1[26]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(read_data1[27]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .X(read_data1[28]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .X(read_data1[29]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(read_data1[2]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(read_data1[30]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(read_data1[31]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(read_data1[3]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(read_data1[4]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(read_data1[5]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(read_data1[6]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(read_data1[7]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(read_data1[8]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(read_data1[9]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(read_data2[0]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(read_data2[10]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(read_data2[11]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(read_data2[12]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(read_data2[13]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(read_data2[14]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(read_data2[15]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(read_data2[16]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(read_data2[17]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .X(read_data2[18]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .X(read_data2[19]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(read_data2[1]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(read_data2[20]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(read_data2[21]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .X(read_data2[22]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .X(read_data2[23]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(read_data2[24]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .X(read_data2[25]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .X(read_data2[26]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(read_data2[27]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .X(read_data2[28]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .X(read_data2[29]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .X(read_data2[2]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net99),
    .X(read_data2[30]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net100),
    .X(read_data2[31]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net101),
    .X(read_data2[3]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net102),
    .X(read_data2[4]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net103),
    .X(read_data2[5]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net104),
    .X(read_data2[6]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net105),
    .X(read_data2[7]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net106),
    .X(read_data2[8]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net107),
    .X(read_data2[9]));
 sky130_fd_sc_hd__buf_16 max_cap108 (.A(_0001_),
    .X(net108));
 sky130_fd_sc_hd__buf_16 load_slew109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_16 load_slew110 (.A(_0005_),
    .X(net110));
 sky130_fd_sc_hd__buf_16 load_slew111 (.A(_0015_),
    .X(net111));
 sky130_fd_sc_hd__buf_16 max_cap112 (.A(_0028_),
    .X(net112));
 sky130_fd_sc_hd__buf_16 load_slew113 (.A(_0031_),
    .X(net113));
 sky130_fd_sc_hd__buf_16 load_slew114 (.A(_0002_),
    .X(net114));
 sky130_fd_sc_hd__buf_16 load_slew115 (.A(_0006_),
    .X(net115));
 sky130_fd_sc_hd__buf_16 load_slew116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_16 load_slew117 (.A(_0007_),
    .X(net117));
 sky130_fd_sc_hd__buf_16 load_slew118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__buf_16 load_slew119 (.A(_0012_),
    .X(net119));
 sky130_fd_sc_hd__buf_12 max_cap120 (.A(_0025_),
    .X(net120));
 sky130_fd_sc_hd__buf_12 max_cap121 (.A(_0029_),
    .X(net121));
 sky130_fd_sc_hd__buf_12 load_slew122 (.A(_0000_),
    .X(net122));
 sky130_fd_sc_hd__buf_16 load_slew123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_16 load_slew124 (.A(_0003_),
    .X(net124));
 sky130_fd_sc_hd__buf_16 load_slew125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_16 load_slew126 (.A(_0004_),
    .X(net126));
 sky130_fd_sc_hd__buf_12 max_cap127 (.A(_0009_),
    .X(net127));
 sky130_fd_sc_hd__buf_12 max_cap128 (.A(_0010_),
    .X(net128));
 sky130_fd_sc_hd__buf_16 max_cap129 (.A(_0013_),
    .X(net129));
 sky130_fd_sc_hd__buf_12 max_cap130 (.A(_0014_),
    .X(net130));
 sky130_fd_sc_hd__buf_16 load_slew131 (.A(_0020_),
    .X(net131));
 sky130_fd_sc_hd__buf_12 max_cap132 (.A(_0026_),
    .X(net132));
 sky130_fd_sc_hd__buf_12 max_cap133 (.A(_0027_),
    .X(net133));
 sky130_fd_sc_hd__buf_16 max_cap134 (.A(_0030_),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload4 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload7 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkinv_1 clkload8 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkinv_1 clkload9 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkinv_1 clkload10 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkinv_1 clkload11 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload12 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__bufinv_16 clkload13 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkinv_1 clkload14 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload15 (.A(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload16 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkinv_1 clkload17 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload18 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinv_1 clkload19 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinv_1 clkload20 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_2 clkload21 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkinv_2 clkload22 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__bufinv_16 clkload23 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__bufinv_16 clkload24 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_2 clkload25 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkinv_1 clkload26 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkinv_1 clkload27 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkinv_1 clkload28 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload29 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkinv_2 clkload30 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkinv_2 clkload31 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__bufinv_16 clkload32 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkinv_1 clkload33 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload34 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkinv_2 clkload35 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkinv_2 clkload36 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkinv_1 clkload37 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkinv_1 clkload38 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkinv_2 clkload39 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__bufinv_16 clkload40 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__bufinv_16 clkload41 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload42 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkinv_1 clkload43 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload44 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload45 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload46 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload47 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload48 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkinv_1 clkload49 (.A(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload50 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload51 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload52 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkinv_1 clkload53 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload54 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinv_2 clkload55 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkinv_2 clkload56 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinv_2 clkload57 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__bufinv_16 clkload58 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_2 clkload59 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkinv_2 clkload60 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__bufinv_16 clkload61 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkinv_2 clkload62 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__inv_6 clkload63 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinv_1 clkload64 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkinv_2 clkload65 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload66 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkinv_1 clkload67 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload68 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload69 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload70 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload71 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload72 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinv_2 clkload73 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkinv_1 clkload74 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload75 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_1 clkload76 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__bufinv_16 clkload77 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__bufinv_16 clkload78 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__bufinv_16 clkload79 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkinv_2 clkload80 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload81 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload82 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkinv_1 clkload83 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkinv_2 clkload84 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkinv_1 clkload85 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload86 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkinv_1 clkload87 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkinv_1 clkload88 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__bufinv_16 clkload89 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__bufinv_16 clkload90 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__bufinv_16 clkload91 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkinv_2 clkload92 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkinv_2 clkload93 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkinv_2 clkload94 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__bufinv_16 clkload95 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkinv_2 clkload96 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload97 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinv_2 clkload98 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__bufinv_16 clkload99 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload100 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__bufinv_16 clkload101 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(write_data[23]),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(write_data[29]),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(write_data[21]),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(write_data[22]),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(write_data[25]),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(write_data[1]),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(write_data[31]),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(write_data[27]),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(write_data[30]),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(write_data[5]),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(write_data[15]),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(write_data[4]),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(write_data[14]),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(write_data[20]),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(write_data[24]),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(write_data[26]),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(write_data[19]),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(write_data[10]),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(write_data[0]),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(write_data[11]),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(write_data[13]),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(write_data[17]),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(write_data[8]),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(write_data[16]),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(write_data[9]),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(write_data[2]),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(write_data[28]),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(write_data[7]),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(write_data[3]),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(write_data[18]),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(write_data[12]),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(write_data[6]),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(read_addr2[4]),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(read_addr1[4]),
    .X(net168));
 sky130_fd_sc_hd__buf_16 max_cap1 (.A(_0011_),
    .X(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0076_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_2357_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_2369_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_2401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_2514_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_2514_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_2348_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_2349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_2430_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_630 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_480 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_542 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_684 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_684 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_695 ();
endmodule
