module barrel_rotator (direction,
    data_in,
    data_out,
    rotate_amount);
 input direction;
 input [7:0] data_in;
 output [7:0] data_out;
 input [2:0] rotate_amount;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 BUF_X2 _148_ (.A(data_in[0]),
    .Z(_071_));
 BUF_X4 _149_ (.A(net1),
    .Z(_072_));
 CLKBUF_X3 _150_ (.A(_072_),
    .Z(_073_));
 BUF_X4 _151_ (.A(_073_),
    .Z(_074_));
 BUF_X4 _152_ (.A(rotate_amount[1]),
    .Z(_075_));
 INV_X4 _153_ (.A(_075_),
    .ZN(_076_));
 BUF_X4 _154_ (.A(rotate_amount[0]),
    .Z(_077_));
 INV_X2 _155_ (.A(_077_),
    .ZN(_078_));
 NAND2_X2 _156_ (.A1(_076_),
    .A2(_078_),
    .ZN(_079_));
 NOR2_X2 _157_ (.A1(_074_),
    .A2(_079_),
    .ZN(_080_));
 NAND2_X1 _158_ (.A1(_071_),
    .A2(_080_),
    .ZN(_081_));
 CLKBUF_X3 _159_ (.A(_075_),
    .Z(_082_));
 INV_X1 _160_ (.A(_072_),
    .ZN(_083_));
 CLKBUF_X3 _161_ (.A(_083_),
    .Z(_084_));
 CLKBUF_X2 _162_ (.A(data_in[6]),
    .Z(_085_));
 BUF_X2 _163_ (.A(data_in[7]),
    .Z(_086_));
 BUF_X8 _164_ (.A(_077_),
    .Z(_087_));
 MUX2_X1 _165_ (.A(_085_),
    .B(_086_),
    .S(_087_),
    .Z(_088_));
 NOR2_X1 _166_ (.A1(_084_),
    .A2(_088_),
    .ZN(_089_));
 BUF_X4 _167_ (.A(_087_),
    .Z(_090_));
 BUF_X2 _168_ (.A(data_in[2]),
    .Z(_091_));
 OR2_X1 _169_ (.A1(_090_),
    .A2(_091_),
    .ZN(_092_));
 BUF_X4 _170_ (.A(data_in[3]),
    .Z(_093_));
 CLKBUF_X3 _171_ (.A(_078_),
    .Z(_094_));
 OAI21_X1 _172_ (.A(_092_),
    .B1(_093_),
    .B2(_094_),
    .ZN(_095_));
 AOI21_X1 _173_ (.A(_089_),
    .B1(_095_),
    .B2(_084_),
    .ZN(_096_));
 CLKBUF_X3 _174_ (.A(_075_),
    .Z(_097_));
 BUF_X2 _175_ (.A(data_in[4]),
    .Z(_098_));
 BUF_X4 _176_ (.A(direction),
    .Z(_099_));
 OAI22_X1 _177_ (.A1(_097_),
    .A2(_074_),
    .B1(_098_),
    .B2(_099_),
    .ZN(_100_));
 NAND2_X1 _178_ (.A1(_094_),
    .A2(_100_),
    .ZN(_101_));
 INV_X4 _179_ (.A(_099_),
    .ZN(_102_));
 BUF_X2 _180_ (.A(data_in[1]),
    .Z(_103_));
 BUF_X2 _181_ (.A(data_in[5]),
    .Z(_104_));
 MUX2_X1 _182_ (.A(_103_),
    .B(_104_),
    .S(_072_),
    .Z(_105_));
 NOR2_X1 _183_ (.A1(_078_),
    .A2(_105_),
    .ZN(_106_));
 OAI21_X1 _184_ (.A(_102_),
    .B1(_106_),
    .B2(_082_),
    .ZN(_107_));
 AOI22_X1 _185_ (.A1(_082_),
    .A2(_096_),
    .B1(_101_),
    .B2(_107_),
    .ZN(_108_));
 NAND2_X1 _186_ (.A1(_073_),
    .A2(_098_),
    .ZN(_109_));
 CLKBUF_X3 _187_ (.A(_087_),
    .Z(_110_));
 MUX2_X2 _188_ (.A(_086_),
    .B(_093_),
    .S(net1),
    .Z(_111_));
 NAND2_X1 _189_ (.A1(_110_),
    .A2(_111_),
    .ZN(_112_));
 OAI221_X1 _190_ (.A(_099_),
    .B1(_079_),
    .B2(_109_),
    .C1(_112_),
    .C2(_097_),
    .ZN(_113_));
 MUX2_X2 _191_ (.A(_104_),
    .B(_103_),
    .S(_072_),
    .Z(_114_));
 NAND2_X1 _192_ (.A1(_110_),
    .A2(_114_),
    .ZN(_115_));
 MUX2_X2 _193_ (.A(_085_),
    .B(_091_),
    .S(_072_),
    .Z(_116_));
 NAND2_X1 _194_ (.A1(_094_),
    .A2(_116_),
    .ZN(_117_));
 NAND2_X1 _195_ (.A1(_115_),
    .A2(_117_),
    .ZN(_118_));
 AOI21_X1 _196_ (.A(_113_),
    .B1(_118_),
    .B2(_082_),
    .ZN(_119_));
 OAI21_X1 _197_ (.A(_081_),
    .B1(_108_),
    .B2(_119_),
    .ZN(net2));
 NOR3_X1 _198_ (.A1(_074_),
    .A2(_103_),
    .A3(_079_),
    .ZN(_120_));
 AOI21_X1 _199_ (.A(_090_),
    .B1(_086_),
    .B2(_072_),
    .ZN(_121_));
 INV_X1 _200_ (.A(_093_),
    .ZN(_122_));
 OAI21_X1 _201_ (.A(_121_),
    .B1(_122_),
    .B2(_073_),
    .ZN(_123_));
 MUX2_X1 _202_ (.A(_098_),
    .B(_071_),
    .S(_072_),
    .Z(_124_));
 OR2_X1 _203_ (.A1(_078_),
    .A2(_124_),
    .ZN(_125_));
 NAND3_X1 _204_ (.A1(_082_),
    .A2(_123_),
    .A3(_125_),
    .ZN(_126_));
 NOR2_X2 _205_ (.A1(_075_),
    .A2(_077_),
    .ZN(_127_));
 OR2_X1 _206_ (.A1(_083_),
    .A2(_104_),
    .ZN(_128_));
 MUX2_X1 _207_ (.A(_091_),
    .B(_085_),
    .S(_072_),
    .Z(_129_));
 NOR2_X2 _208_ (.A1(_075_),
    .A2(_078_),
    .ZN(_130_));
 AOI221_X1 _209_ (.A(_099_),
    .B1(_127_),
    .B2(_128_),
    .C1(_129_),
    .C2(_130_),
    .ZN(_131_));
 AND2_X1 _210_ (.A1(_126_),
    .A2(_131_),
    .ZN(_132_));
 NAND3_X1 _211_ (.A1(_097_),
    .A2(_110_),
    .A3(_116_),
    .ZN(_133_));
 MUX2_X1 _212_ (.A(_071_),
    .B(_098_),
    .S(_072_),
    .Z(_134_));
 NAND3_X1 _213_ (.A1(_076_),
    .A2(_090_),
    .A3(_134_),
    .ZN(_135_));
 NAND3_X1 _214_ (.A1(_075_),
    .A2(_094_),
    .A3(_111_),
    .ZN(_136_));
 NAND4_X1 _215_ (.A1(_099_),
    .A2(_133_),
    .A3(_135_),
    .A4(_136_),
    .ZN(_137_));
 AOI21_X1 _216_ (.A(_137_),
    .B1(_128_),
    .B2(_127_),
    .ZN(_138_));
 NOR3_X1 _217_ (.A1(_120_),
    .A2(_132_),
    .A3(_138_),
    .ZN(net3));
 OAI21_X1 _218_ (.A(_075_),
    .B1(_090_),
    .B2(_134_),
    .ZN(_139_));
 INV_X1 _219_ (.A(_111_),
    .ZN(_140_));
 AOI21_X1 _220_ (.A(_139_),
    .B1(_140_),
    .B2(_110_),
    .ZN(_141_));
 NOR3_X1 _221_ (.A1(_083_),
    .A2(_087_),
    .A3(_085_),
    .ZN(_142_));
 NOR3_X1 _222_ (.A1(_097_),
    .A2(_106_),
    .A3(_142_),
    .ZN(_143_));
 OAI33_X1 _223_ (.A1(_074_),
    .A2(_091_),
    .A3(_079_),
    .B1(_141_),
    .B2(_143_),
    .B3(_102_),
    .ZN(_144_));
 NOR3_X1 _224_ (.A1(_074_),
    .A2(_094_),
    .A3(_093_),
    .ZN(_145_));
 OAI21_X1 _225_ (.A(_076_),
    .B1(_089_),
    .B2(_145_),
    .ZN(_146_));
 MUX2_X1 _226_ (.A(_114_),
    .B(_124_),
    .S(_094_),
    .Z(_147_));
 OAI21_X1 _227_ (.A(_146_),
    .B1(_147_),
    .B2(_076_),
    .ZN(_000_));
 AOI21_X1 _228_ (.A(_144_),
    .B1(_000_),
    .B2(_102_),
    .ZN(net4));
 NOR2_X1 _229_ (.A1(_082_),
    .A2(_121_),
    .ZN(_001_));
 MUX2_X1 _230_ (.A(_114_),
    .B(_116_),
    .S(_110_),
    .Z(_002_));
 AOI22_X2 _231_ (.A1(_125_),
    .A2(_001_),
    .B1(_002_),
    .B2(_082_),
    .ZN(_003_));
 AOI21_X1 _232_ (.A(_099_),
    .B1(_080_),
    .B2(_093_),
    .ZN(_004_));
 AOI21_X1 _233_ (.A(_102_),
    .B1(_080_),
    .B2(_093_),
    .ZN(_005_));
 MUX2_X1 _234_ (.A(_086_),
    .B(_085_),
    .S(_087_),
    .Z(_006_));
 NAND2_X1 _235_ (.A1(_073_),
    .A2(_006_),
    .ZN(_007_));
 NAND3_X1 _236_ (.A1(_084_),
    .A2(_110_),
    .A3(_091_),
    .ZN(_008_));
 AOI21_X1 _237_ (.A(_097_),
    .B1(_007_),
    .B2(_008_),
    .ZN(_009_));
 MUX2_X1 _238_ (.A(_105_),
    .B(_134_),
    .S(_110_),
    .Z(_010_));
 AOI21_X2 _239_ (.A(_009_),
    .B1(_010_),
    .B2(_082_),
    .ZN(_011_));
 AOI22_X2 _240_ (.A1(_003_),
    .A2(_004_),
    .B1(_005_),
    .B2(_011_),
    .ZN(net5));
 OAI21_X1 _241_ (.A(_127_),
    .B1(_071_),
    .B2(_084_),
    .ZN(_012_));
 NAND2_X1 _242_ (.A1(_102_),
    .A2(_012_),
    .ZN(_013_));
 AOI21_X1 _243_ (.A(_082_),
    .B1(_110_),
    .B2(_114_),
    .ZN(_014_));
 INV_X1 _244_ (.A(_014_),
    .ZN(_015_));
 NAND3_X1 _245_ (.A1(_082_),
    .A2(_117_),
    .A3(_112_),
    .ZN(_016_));
 AOI21_X1 _246_ (.A(_013_),
    .B1(_015_),
    .B2(_016_),
    .ZN(_017_));
 NAND3_X1 _247_ (.A1(_097_),
    .A2(_110_),
    .A3(_103_),
    .ZN(_018_));
 OAI21_X1 _248_ (.A(_094_),
    .B1(_091_),
    .B2(_076_),
    .ZN(_019_));
 AOI21_X1 _249_ (.A(_074_),
    .B1(_018_),
    .B2(_019_),
    .ZN(_020_));
 MUX2_X1 _250_ (.A(_085_),
    .B(_104_),
    .S(_087_),
    .Z(_021_));
 NAND3_X1 _251_ (.A1(_097_),
    .A2(_073_),
    .A3(_021_),
    .ZN(_022_));
 NAND2_X1 _252_ (.A1(_099_),
    .A2(_022_),
    .ZN(_023_));
 MUX2_X1 _253_ (.A(_071_),
    .B(_086_),
    .S(_087_),
    .Z(_024_));
 NAND2_X1 _254_ (.A1(_073_),
    .A2(_024_),
    .ZN(_025_));
 NAND3_X1 _255_ (.A1(_084_),
    .A2(_090_),
    .A3(_093_),
    .ZN(_026_));
 AOI21_X1 _256_ (.A(_097_),
    .B1(_025_),
    .B2(_026_),
    .ZN(_027_));
 OAI33_X1 _257_ (.A1(_074_),
    .A2(_098_),
    .A3(_079_),
    .B1(_020_),
    .B2(_023_),
    .B3(_027_),
    .ZN(_028_));
 NOR2_X1 _258_ (.A1(_017_),
    .A2(_028_),
    .ZN(net6));
 OAI21_X1 _259_ (.A(_127_),
    .B1(_103_),
    .B2(_083_),
    .ZN(_029_));
 NAND2_X1 _260_ (.A1(_102_),
    .A2(_029_),
    .ZN(_030_));
 MUX2_X1 _261_ (.A(_111_),
    .B(_134_),
    .S(_087_),
    .Z(_031_));
 AOI221_X2 _262_ (.A(_030_),
    .B1(_031_),
    .B2(_097_),
    .C1(_116_),
    .C2(_130_),
    .ZN(_032_));
 NAND3_X1 _263_ (.A1(_084_),
    .A2(_110_),
    .A3(_098_),
    .ZN(_033_));
 MUX2_X1 _264_ (.A(_103_),
    .B(_071_),
    .S(_087_),
    .Z(_034_));
 NAND2_X1 _265_ (.A1(_073_),
    .A2(_034_),
    .ZN(_035_));
 AOI21_X1 _266_ (.A(_097_),
    .B1(_033_),
    .B2(_035_),
    .ZN(_036_));
 NAND3_X1 _267_ (.A1(_075_),
    .A2(_090_),
    .A3(_091_),
    .ZN(_037_));
 OAI21_X1 _268_ (.A(_094_),
    .B1(_093_),
    .B2(_076_),
    .ZN(_038_));
 AOI21_X1 _269_ (.A(_074_),
    .B1(_037_),
    .B2(_038_),
    .ZN(_039_));
 NAND3_X1 _270_ (.A1(_075_),
    .A2(_073_),
    .A3(_006_),
    .ZN(_040_));
 NAND2_X1 _271_ (.A1(_099_),
    .A2(_040_),
    .ZN(_041_));
 OAI33_X1 _272_ (.A1(_074_),
    .A2(_104_),
    .A3(_079_),
    .B1(_036_),
    .B2(_039_),
    .B3(_041_),
    .ZN(_042_));
 NOR2_X1 _273_ (.A1(_032_),
    .A2(_042_),
    .ZN(net7));
 INV_X1 _274_ (.A(_130_),
    .ZN(_043_));
 MUX2_X1 _275_ (.A(_114_),
    .B(_111_),
    .S(_102_),
    .Z(_044_));
 OAI22_X1 _276_ (.A1(_079_),
    .A2(_116_),
    .B1(_043_),
    .B2(_044_),
    .ZN(_045_));
 MUX2_X1 _277_ (.A(_098_),
    .B(_104_),
    .S(_090_),
    .Z(_046_));
 NAND2_X1 _278_ (.A1(_074_),
    .A2(_046_),
    .ZN(_047_));
 MUX2_X1 _279_ (.A(_071_),
    .B(_103_),
    .S(_090_),
    .Z(_048_));
 NAND2_X1 _280_ (.A1(_084_),
    .A2(_048_),
    .ZN(_049_));
 OAI221_X1 _281_ (.A(_076_),
    .B1(_094_),
    .B2(_111_),
    .C1(_092_),
    .C2(_084_),
    .ZN(_050_));
 NAND3_X1 _282_ (.A1(_047_),
    .A2(_049_),
    .A3(_050_),
    .ZN(_051_));
 NAND2_X1 _283_ (.A1(_102_),
    .A2(_051_),
    .ZN(_052_));
 MUX2_X1 _284_ (.A(_098_),
    .B(_093_),
    .S(_090_),
    .Z(_053_));
 NAND2_X1 _285_ (.A1(_084_),
    .A2(_053_),
    .ZN(_054_));
 OAI221_X1 _286_ (.A(_076_),
    .B1(_094_),
    .B2(_114_),
    .C1(_092_),
    .C2(_084_),
    .ZN(_055_));
 NAND3_X1 _287_ (.A1(_025_),
    .A2(_054_),
    .A3(_055_),
    .ZN(_056_));
 NAND2_X1 _288_ (.A1(_099_),
    .A2(_056_),
    .ZN(_057_));
 AOI21_X1 _289_ (.A(_045_),
    .B1(_052_),
    .B2(_057_),
    .ZN(net8));
 INV_X1 _290_ (.A(_086_),
    .ZN(_058_));
 NAND2_X1 _291_ (.A1(_073_),
    .A2(_122_),
    .ZN(_059_));
 AOI221_X2 _292_ (.A(_102_),
    .B1(_116_),
    .B2(_130_),
    .C1(_059_),
    .C2(_127_),
    .ZN(_060_));
 OR2_X1 _293_ (.A1(_090_),
    .A2(_114_),
    .ZN(_061_));
 NAND3_X1 _294_ (.A1(_082_),
    .A2(_125_),
    .A3(_061_),
    .ZN(_062_));
 MUX2_X1 _295_ (.A(_093_),
    .B(_098_),
    .S(_087_),
    .Z(_063_));
 NOR2_X1 _296_ (.A1(_083_),
    .A2(_063_),
    .ZN(_064_));
 NOR3_X1 _297_ (.A1(_073_),
    .A2(_078_),
    .A3(_071_),
    .ZN(_065_));
 OAI21_X1 _298_ (.A(_076_),
    .B1(_064_),
    .B2(_065_),
    .ZN(_066_));
 MUX2_X1 _299_ (.A(_103_),
    .B(_091_),
    .S(_077_),
    .Z(_067_));
 MUX2_X1 _300_ (.A(_104_),
    .B(_085_),
    .S(_077_),
    .Z(_068_));
 MUX2_X1 _301_ (.A(_067_),
    .B(_068_),
    .S(_072_),
    .Z(_069_));
 OAI21_X1 _302_ (.A(_066_),
    .B1(_069_),
    .B2(_076_),
    .ZN(_070_));
 AOI222_X2 _303_ (.A1(_058_),
    .A2(_080_),
    .B1(_060_),
    .B2(_062_),
    .C1(_070_),
    .C2(_102_),
    .ZN(net9));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_87 ();
 BUF_X1 input1 (.A(rotate_amount[2]),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(data_out[0]));
 BUF_X1 output3 (.A(net3),
    .Z(data_out[1]));
 BUF_X1 output4 (.A(net4),
    .Z(data_out[2]));
 BUF_X1 output5 (.A(net5),
    .Z(data_out[3]));
 BUF_X1 output6 (.A(net6),
    .Z(data_out[4]));
 BUF_X1 output7 (.A(net7),
    .Z(data_out[5]));
 BUF_X1 output8 (.A(net8),
    .Z(data_out[6]));
 BUF_X1 output9 (.A(net9),
    .Z(data_out[7]));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X16 FILLER_0_97 ();
 FILLCELL_X8 FILLER_0_113 ();
 FILLCELL_X1 FILLER_0_121 ();
 FILLCELL_X32 FILLER_0_125 ();
 FILLCELL_X32 FILLER_0_157 ();
 FILLCELL_X32 FILLER_0_189 ();
 FILLCELL_X32 FILLER_0_221 ();
 FILLCELL_X32 FILLER_0_253 ();
 FILLCELL_X32 FILLER_0_285 ();
 FILLCELL_X8 FILLER_0_317 ();
 FILLCELL_X1 FILLER_0_325 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X4 FILLER_1_321 ();
 FILLCELL_X1 FILLER_1_325 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X4 FILLER_2_321 ();
 FILLCELL_X1 FILLER_2_325 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X4 FILLER_3_321 ();
 FILLCELL_X1 FILLER_3_325 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X4 FILLER_4_321 ();
 FILLCELL_X1 FILLER_4_325 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X4 FILLER_5_321 ();
 FILLCELL_X1 FILLER_5_325 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X4 FILLER_6_321 ();
 FILLCELL_X1 FILLER_6_325 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X4 FILLER_7_321 ();
 FILLCELL_X1 FILLER_7_325 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X4 FILLER_8_321 ();
 FILLCELL_X1 FILLER_8_325 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X8 FILLER_9_97 ();
 FILLCELL_X2 FILLER_9_105 ();
 FILLCELL_X1 FILLER_9_107 ();
 FILLCELL_X2 FILLER_9_112 ();
 FILLCELL_X32 FILLER_9_122 ();
 FILLCELL_X32 FILLER_9_154 ();
 FILLCELL_X32 FILLER_9_186 ();
 FILLCELL_X32 FILLER_9_218 ();
 FILLCELL_X32 FILLER_9_250 ();
 FILLCELL_X32 FILLER_9_282 ();
 FILLCELL_X8 FILLER_9_314 ();
 FILLCELL_X4 FILLER_9_322 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X4 FILLER_10_321 ();
 FILLCELL_X1 FILLER_10_325 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X8 FILLER_11_97 ();
 FILLCELL_X4 FILLER_11_105 ();
 FILLCELL_X2 FILLER_11_109 ();
 FILLCELL_X32 FILLER_11_115 ();
 FILLCELL_X32 FILLER_11_147 ();
 FILLCELL_X32 FILLER_11_179 ();
 FILLCELL_X32 FILLER_11_211 ();
 FILLCELL_X32 FILLER_11_243 ();
 FILLCELL_X32 FILLER_11_275 ();
 FILLCELL_X16 FILLER_11_307 ();
 FILLCELL_X2 FILLER_11_323 ();
 FILLCELL_X1 FILLER_11_325 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X4 FILLER_12_321 ();
 FILLCELL_X1 FILLER_12_325 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X4 FILLER_13_321 ();
 FILLCELL_X1 FILLER_13_325 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X4 FILLER_14_104 ();
 FILLCELL_X2 FILLER_14_108 ();
 FILLCELL_X2 FILLER_14_117 ();
 FILLCELL_X4 FILLER_14_126 ();
 FILLCELL_X1 FILLER_14_130 ();
 FILLCELL_X32 FILLER_14_138 ();
 FILLCELL_X32 FILLER_14_170 ();
 FILLCELL_X32 FILLER_14_202 ();
 FILLCELL_X32 FILLER_14_234 ();
 FILLCELL_X32 FILLER_14_266 ();
 FILLCELL_X16 FILLER_14_298 ();
 FILLCELL_X8 FILLER_14_314 ();
 FILLCELL_X4 FILLER_14_322 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X16 FILLER_15_33 ();
 FILLCELL_X8 FILLER_15_49 ();
 FILLCELL_X4 FILLER_15_57 ();
 FILLCELL_X16 FILLER_15_65 ();
 FILLCELL_X2 FILLER_15_81 ();
 FILLCELL_X1 FILLER_15_83 ();
 FILLCELL_X1 FILLER_15_102 ();
 FILLCELL_X1 FILLER_15_106 ();
 FILLCELL_X4 FILLER_15_121 ();
 FILLCELL_X2 FILLER_15_125 ();
 FILLCELL_X4 FILLER_15_130 ();
 FILLCELL_X2 FILLER_15_140 ();
 FILLCELL_X1 FILLER_15_142 ();
 FILLCELL_X8 FILLER_15_164 ();
 FILLCELL_X32 FILLER_15_179 ();
 FILLCELL_X32 FILLER_15_211 ();
 FILLCELL_X32 FILLER_15_243 ();
 FILLCELL_X32 FILLER_15_275 ();
 FILLCELL_X16 FILLER_15_307 ();
 FILLCELL_X2 FILLER_15_323 ();
 FILLCELL_X1 FILLER_15_325 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X8 FILLER_16_33 ();
 FILLCELL_X2 FILLER_16_41 ();
 FILLCELL_X32 FILLER_16_47 ();
 FILLCELL_X4 FILLER_16_79 ();
 FILLCELL_X4 FILLER_16_90 ();
 FILLCELL_X4 FILLER_16_118 ();
 FILLCELL_X2 FILLER_16_122 ();
 FILLCELL_X1 FILLER_16_124 ();
 FILLCELL_X4 FILLER_16_128 ();
 FILLCELL_X2 FILLER_16_132 ();
 FILLCELL_X16 FILLER_16_150 ();
 FILLCELL_X4 FILLER_16_166 ();
 FILLCELL_X1 FILLER_16_170 ();
 FILLCELL_X32 FILLER_16_178 ();
 FILLCELL_X32 FILLER_16_210 ();
 FILLCELL_X32 FILLER_16_242 ();
 FILLCELL_X32 FILLER_16_274 ();
 FILLCELL_X16 FILLER_16_306 ();
 FILLCELL_X4 FILLER_16_322 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X16 FILLER_17_65 ();
 FILLCELL_X8 FILLER_17_81 ();
 FILLCELL_X2 FILLER_17_89 ();
 FILLCELL_X1 FILLER_17_91 ();
 FILLCELL_X4 FILLER_17_95 ();
 FILLCELL_X2 FILLER_17_103 ();
 FILLCELL_X1 FILLER_17_105 ();
 FILLCELL_X1 FILLER_17_111 ();
 FILLCELL_X16 FILLER_17_116 ();
 FILLCELL_X2 FILLER_17_132 ();
 FILLCELL_X1 FILLER_17_134 ();
 FILLCELL_X1 FILLER_17_139 ();
 FILLCELL_X2 FILLER_17_154 ();
 FILLCELL_X4 FILLER_17_168 ();
 FILLCELL_X2 FILLER_17_172 ();
 FILLCELL_X32 FILLER_17_177 ();
 FILLCELL_X32 FILLER_17_209 ();
 FILLCELL_X32 FILLER_17_241 ();
 FILLCELL_X16 FILLER_17_273 ();
 FILLCELL_X1 FILLER_17_289 ();
 FILLCELL_X16 FILLER_17_296 ();
 FILLCELL_X8 FILLER_17_312 ();
 FILLCELL_X4 FILLER_17_320 ();
 FILLCELL_X2 FILLER_17_324 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_9 ();
 FILLCELL_X2 FILLER_18_13 ();
 FILLCELL_X32 FILLER_18_19 ();
 FILLCELL_X16 FILLER_18_51 ();
 FILLCELL_X8 FILLER_18_67 ();
 FILLCELL_X4 FILLER_18_75 ();
 FILLCELL_X2 FILLER_18_79 ();
 FILLCELL_X1 FILLER_18_81 ();
 FILLCELL_X1 FILLER_18_95 ();
 FILLCELL_X16 FILLER_18_105 ();
 FILLCELL_X8 FILLER_18_121 ();
 FILLCELL_X4 FILLER_18_129 ();
 FILLCELL_X2 FILLER_18_145 ();
 FILLCELL_X1 FILLER_18_147 ();
 FILLCELL_X32 FILLER_18_160 ();
 FILLCELL_X32 FILLER_18_192 ();
 FILLCELL_X32 FILLER_18_224 ();
 FILLCELL_X32 FILLER_18_256 ();
 FILLCELL_X32 FILLER_18_288 ();
 FILLCELL_X4 FILLER_18_320 ();
 FILLCELL_X2 FILLER_18_324 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_5 ();
 FILLCELL_X32 FILLER_19_14 ();
 FILLCELL_X32 FILLER_19_46 ();
 FILLCELL_X8 FILLER_19_78 ();
 FILLCELL_X4 FILLER_19_105 ();
 FILLCELL_X32 FILLER_19_120 ();
 FILLCELL_X2 FILLER_19_152 ();
 FILLCELL_X1 FILLER_19_154 ();
 FILLCELL_X4 FILLER_19_157 ();
 FILLCELL_X2 FILLER_19_161 ();
 FILLCELL_X1 FILLER_19_163 ();
 FILLCELL_X32 FILLER_19_167 ();
 FILLCELL_X32 FILLER_19_199 ();
 FILLCELL_X32 FILLER_19_231 ();
 FILLCELL_X32 FILLER_19_263 ();
 FILLCELL_X16 FILLER_19_295 ();
 FILLCELL_X8 FILLER_19_311 ();
 FILLCELL_X4 FILLER_19_319 ();
 FILLCELL_X2 FILLER_19_323 ();
 FILLCELL_X1 FILLER_19_325 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X16 FILLER_20_65 ();
 FILLCELL_X4 FILLER_20_81 ();
 FILLCELL_X1 FILLER_20_85 ();
 FILLCELL_X16 FILLER_20_116 ();
 FILLCELL_X2 FILLER_20_132 ();
 FILLCELL_X16 FILLER_20_138 ();
 FILLCELL_X2 FILLER_20_157 ();
 FILLCELL_X1 FILLER_20_159 ();
 FILLCELL_X32 FILLER_20_177 ();
 FILLCELL_X32 FILLER_20_209 ();
 FILLCELL_X32 FILLER_20_241 ();
 FILLCELL_X32 FILLER_20_273 ();
 FILLCELL_X16 FILLER_20_305 ();
 FILLCELL_X4 FILLER_20_321 ();
 FILLCELL_X1 FILLER_20_325 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_17 ();
 FILLCELL_X2 FILLER_21_21 ();
 FILLCELL_X1 FILLER_21_23 ();
 FILLCELL_X8 FILLER_21_27 ();
 FILLCELL_X32 FILLER_21_38 ();
 FILLCELL_X8 FILLER_21_70 ();
 FILLCELL_X4 FILLER_21_78 ();
 FILLCELL_X2 FILLER_21_82 ();
 FILLCELL_X1 FILLER_21_84 ();
 FILLCELL_X2 FILLER_21_99 ();
 FILLCELL_X4 FILLER_21_105 ();
 FILLCELL_X2 FILLER_21_117 ();
 FILLCELL_X1 FILLER_21_119 ();
 FILLCELL_X8 FILLER_21_124 ();
 FILLCELL_X2 FILLER_21_132 ();
 FILLCELL_X2 FILLER_21_138 ();
 FILLCELL_X8 FILLER_21_145 ();
 FILLCELL_X2 FILLER_21_156 ();
 FILLCELL_X1 FILLER_21_164 ();
 FILLCELL_X4 FILLER_21_169 ();
 FILLCELL_X2 FILLER_21_173 ();
 FILLCELL_X32 FILLER_21_177 ();
 FILLCELL_X32 FILLER_21_209 ();
 FILLCELL_X32 FILLER_21_241 ();
 FILLCELL_X32 FILLER_21_273 ();
 FILLCELL_X16 FILLER_21_305 ();
 FILLCELL_X4 FILLER_21_321 ();
 FILLCELL_X1 FILLER_21_325 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X16 FILLER_22_65 ();
 FILLCELL_X8 FILLER_22_81 ();
 FILLCELL_X2 FILLER_22_99 ();
 FILLCELL_X2 FILLER_22_105 ();
 FILLCELL_X1 FILLER_22_107 ();
 FILLCELL_X4 FILLER_22_119 ();
 FILLCELL_X2 FILLER_22_127 ();
 FILLCELL_X1 FILLER_22_137 ();
 FILLCELL_X1 FILLER_22_143 ();
 FILLCELL_X8 FILLER_22_147 ();
 FILLCELL_X2 FILLER_22_155 ();
 FILLCELL_X4 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_169 ();
 FILLCELL_X32 FILLER_22_201 ();
 FILLCELL_X32 FILLER_22_233 ();
 FILLCELL_X16 FILLER_22_265 ();
 FILLCELL_X4 FILLER_22_281 ();
 FILLCELL_X2 FILLER_22_285 ();
 FILLCELL_X1 FILLER_22_287 ();
 FILLCELL_X32 FILLER_22_291 ();
 FILLCELL_X2 FILLER_22_323 ();
 FILLCELL_X1 FILLER_22_325 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X16 FILLER_23_65 ();
 FILLCELL_X8 FILLER_23_81 ();
 FILLCELL_X4 FILLER_23_89 ();
 FILLCELL_X2 FILLER_23_93 ();
 FILLCELL_X1 FILLER_23_95 ();
 FILLCELL_X2 FILLER_23_100 ();
 FILLCELL_X4 FILLER_23_113 ();
 FILLCELL_X1 FILLER_23_117 ();
 FILLCELL_X16 FILLER_23_129 ();
 FILLCELL_X4 FILLER_23_145 ();
 FILLCELL_X1 FILLER_23_149 ();
 FILLCELL_X4 FILLER_23_154 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X4 FILLER_23_321 ();
 FILLCELL_X1 FILLER_23_325 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X4 FILLER_24_65 ();
 FILLCELL_X2 FILLER_24_69 ();
 FILLCELL_X1 FILLER_24_71 ();
 FILLCELL_X4 FILLER_24_85 ();
 FILLCELL_X4 FILLER_24_96 ();
 FILLCELL_X1 FILLER_24_100 ();
 FILLCELL_X4 FILLER_24_127 ();
 FILLCELL_X2 FILLER_24_131 ();
 FILLCELL_X8 FILLER_24_137 ();
 FILLCELL_X4 FILLER_24_145 ();
 FILLCELL_X2 FILLER_24_149 ();
 FILLCELL_X1 FILLER_24_151 ();
 FILLCELL_X4 FILLER_24_165 ();
 FILLCELL_X32 FILLER_24_173 ();
 FILLCELL_X32 FILLER_24_205 ();
 FILLCELL_X32 FILLER_24_237 ();
 FILLCELL_X32 FILLER_24_269 ();
 FILLCELL_X16 FILLER_24_301 ();
 FILLCELL_X8 FILLER_24_317 ();
 FILLCELL_X1 FILLER_24_325 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X4 FILLER_25_65 ();
 FILLCELL_X2 FILLER_25_69 ();
 FILLCELL_X1 FILLER_25_85 ();
 FILLCELL_X1 FILLER_25_100 ();
 FILLCELL_X2 FILLER_25_126 ();
 FILLCELL_X1 FILLER_25_128 ();
 FILLCELL_X1 FILLER_25_133 ();
 FILLCELL_X1 FILLER_25_138 ();
 FILLCELL_X4 FILLER_25_144 ();
 FILLCELL_X2 FILLER_25_148 ();
 FILLCELL_X4 FILLER_25_153 ();
 FILLCELL_X2 FILLER_25_157 ();
 FILLCELL_X2 FILLER_25_168 ();
 FILLCELL_X1 FILLER_25_170 ();
 FILLCELL_X32 FILLER_25_180 ();
 FILLCELL_X32 FILLER_25_212 ();
 FILLCELL_X32 FILLER_25_244 ();
 FILLCELL_X8 FILLER_25_276 ();
 FILLCELL_X2 FILLER_25_284 ();
 FILLCELL_X1 FILLER_25_286 ();
 FILLCELL_X32 FILLER_25_290 ();
 FILLCELL_X4 FILLER_25_322 ();
 FILLCELL_X8 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_9 ();
 FILLCELL_X32 FILLER_26_18 ();
 FILLCELL_X16 FILLER_26_50 ();
 FILLCELL_X8 FILLER_26_66 ();
 FILLCELL_X2 FILLER_26_74 ();
 FILLCELL_X4 FILLER_26_81 ();
 FILLCELL_X2 FILLER_26_88 ();
 FILLCELL_X1 FILLER_26_90 ();
 FILLCELL_X4 FILLER_26_119 ();
 FILLCELL_X4 FILLER_26_127 ();
 FILLCELL_X2 FILLER_26_131 ();
 FILLCELL_X1 FILLER_26_133 ();
 FILLCELL_X4 FILLER_26_138 ();
 FILLCELL_X2 FILLER_26_142 ();
 FILLCELL_X1 FILLER_26_144 ();
 FILLCELL_X2 FILLER_26_156 ();
 FILLCELL_X32 FILLER_26_171 ();
 FILLCELL_X32 FILLER_26_203 ();
 FILLCELL_X32 FILLER_26_235 ();
 FILLCELL_X32 FILLER_26_267 ();
 FILLCELL_X16 FILLER_26_299 ();
 FILLCELL_X8 FILLER_26_315 ();
 FILLCELL_X2 FILLER_26_323 ();
 FILLCELL_X1 FILLER_26_325 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X16 FILLER_27_97 ();
 FILLCELL_X8 FILLER_27_113 ();
 FILLCELL_X4 FILLER_27_121 ();
 FILLCELL_X16 FILLER_27_129 ();
 FILLCELL_X1 FILLER_27_145 ();
 FILLCELL_X32 FILLER_27_160 ();
 FILLCELL_X32 FILLER_27_192 ();
 FILLCELL_X32 FILLER_27_224 ();
 FILLCELL_X32 FILLER_27_256 ();
 FILLCELL_X32 FILLER_27_288 ();
 FILLCELL_X4 FILLER_27_320 ();
 FILLCELL_X2 FILLER_27_324 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X4 FILLER_28_321 ();
 FILLCELL_X1 FILLER_28_325 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X4 FILLER_29_321 ();
 FILLCELL_X1 FILLER_29_325 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X4 FILLER_30_321 ();
 FILLCELL_X1 FILLER_30_325 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X4 FILLER_31_321 ();
 FILLCELL_X1 FILLER_31_325 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X4 FILLER_32_321 ();
 FILLCELL_X1 FILLER_32_325 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X4 FILLER_33_321 ();
 FILLCELL_X1 FILLER_33_325 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X4 FILLER_34_321 ();
 FILLCELL_X1 FILLER_34_325 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X4 FILLER_35_321 ();
 FILLCELL_X1 FILLER_35_325 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X4 FILLER_36_321 ();
 FILLCELL_X1 FILLER_36_325 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X4 FILLER_37_321 ();
 FILLCELL_X1 FILLER_37_325 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X4 FILLER_38_321 ();
 FILLCELL_X1 FILLER_38_325 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X4 FILLER_39_321 ();
 FILLCELL_X1 FILLER_39_325 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X4 FILLER_40_321 ();
 FILLCELL_X1 FILLER_40_325 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X4 FILLER_41_321 ();
 FILLCELL_X1 FILLER_41_325 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X4 FILLER_42_321 ();
 FILLCELL_X1 FILLER_42_325 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X8 FILLER_43_129 ();
 FILLCELL_X4 FILLER_43_137 ();
 FILLCELL_X16 FILLER_43_144 ();
 FILLCELL_X8 FILLER_43_160 ();
 FILLCELL_X2 FILLER_43_168 ();
 FILLCELL_X1 FILLER_43_170 ();
 FILLCELL_X32 FILLER_43_174 ();
 FILLCELL_X32 FILLER_43_206 ();
 FILLCELL_X32 FILLER_43_238 ();
 FILLCELL_X32 FILLER_43_270 ();
 FILLCELL_X16 FILLER_43_302 ();
 FILLCELL_X8 FILLER_43_318 ();
endmodule
