module sequence_detector_fsm (clk,
    enable,
    load_pattern,
    pattern_detected,
    rst_n,
    serial_in,
    config_pattern);
 input clk;
 input enable;
 input load_pattern;
 output pattern_detected;
 input rst_n;
 input serial_in;
 input [3:0] config_pattern;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire \bit_count[0] ;
 wire \bit_count[1] ;
 wire \bit_count[2] ;
 wire \pattern_reg[0] ;
 wire \pattern_reg[1] ;
 wire \pattern_reg[2] ;
 wire \pattern_reg[3] ;
 wire \shift_reg[0] ;
 wire \shift_reg[1] ;
 wire \shift_reg[2] ;
 wire state;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _064_ (.A(_058_),
    .ZN(_061_));
 BUF_X2 _065_ (.A(load_pattern),
    .Z(_012_));
 INV_X1 _066_ (.A(net5),
    .ZN(_013_));
 NOR2_X2 _067_ (.A1(_012_),
    .A2(_013_),
    .ZN(_014_));
 BUF_X4 _068_ (.A(enable),
    .Z(_015_));
 OAI21_X1 _069_ (.A(_014_),
    .B1(\bit_count[0] ),
    .B2(_015_),
    .ZN(_016_));
 INV_X4 _070_ (.A(_015_),
    .ZN(_017_));
 NOR2_X1 _071_ (.A1(_017_),
    .A2(\bit_count[2] ),
    .ZN(_018_));
 MUX2_X1 _072_ (.A(\bit_count[2] ),
    .B(_018_),
    .S(\bit_count[0] ),
    .Z(_019_));
 CLKBUF_X2 _073_ (.A(state),
    .Z(_020_));
 AOI21_X1 _074_ (.A(_016_),
    .B1(_019_),
    .B2(_020_),
    .ZN(_000_));
 INV_X1 _075_ (.A(_014_),
    .ZN(_021_));
 NAND3_X1 _076_ (.A1(_020_),
    .A2(_059_),
    .A3(_018_),
    .ZN(_022_));
 AND2_X1 _077_ (.A1(_020_),
    .A2(\bit_count[2] ),
    .ZN(_023_));
 OAI21_X1 _078_ (.A(\bit_count[1] ),
    .B1(_023_),
    .B2(_017_),
    .ZN(_024_));
 AOI21_X1 _079_ (.A(_021_),
    .B1(_022_),
    .B2(_024_),
    .ZN(_001_));
 OAI21_X1 _080_ (.A(_014_),
    .B1(_017_),
    .B2(_020_),
    .ZN(_025_));
 AOI21_X1 _081_ (.A(\bit_count[2] ),
    .B1(_063_),
    .B2(_015_),
    .ZN(_026_));
 NOR2_X1 _082_ (.A1(_025_),
    .A2(_026_),
    .ZN(_002_));
 XNOR2_X1 _083_ (.A(\pattern_reg[3] ),
    .B(\shift_reg[2] ),
    .ZN(_027_));
 XNOR2_X1 _084_ (.A(\pattern_reg[0] ),
    .B(net6),
    .ZN(_028_));
 NAND2_X1 _085_ (.A1(_027_),
    .A2(_028_),
    .ZN(_029_));
 NOR2_X1 _086_ (.A1(_017_),
    .A2(_062_),
    .ZN(_030_));
 INV_X1 _087_ (.A(\shift_reg[0] ),
    .ZN(_031_));
 INV_X1 _088_ (.A(\pattern_reg[2] ),
    .ZN(_032_));
 AOI22_X1 _089_ (.A1(\pattern_reg[1] ),
    .A2(_031_),
    .B1(_032_),
    .B2(\shift_reg[1] ),
    .ZN(_033_));
 NAND3_X1 _090_ (.A1(_020_),
    .A2(_030_),
    .A3(_033_),
    .ZN(_034_));
 OAI22_X1 _091_ (.A1(\pattern_reg[1] ),
    .A2(_031_),
    .B1(_032_),
    .B2(\shift_reg[1] ),
    .ZN(_035_));
 NOR4_X1 _092_ (.A1(_021_),
    .A2(_029_),
    .A3(_034_),
    .A4(_035_),
    .ZN(_003_));
 NAND2_X1 _093_ (.A1(_015_),
    .A2(net6),
    .ZN(_036_));
 NAND2_X1 _094_ (.A1(_017_),
    .A2(\shift_reg[0] ),
    .ZN(_037_));
 AOI21_X1 _095_ (.A(_021_),
    .B1(_036_),
    .B2(_037_),
    .ZN(_008_));
 NAND2_X1 _096_ (.A1(_015_),
    .A2(\shift_reg[0] ),
    .ZN(_038_));
 NAND2_X1 _097_ (.A1(_017_),
    .A2(\shift_reg[1] ),
    .ZN(_039_));
 AOI21_X1 _098_ (.A(_021_),
    .B1(_038_),
    .B2(_039_),
    .ZN(_009_));
 NAND2_X1 _099_ (.A1(_015_),
    .A2(\shift_reg[1] ),
    .ZN(_040_));
 NAND2_X1 _100_ (.A1(_017_),
    .A2(\shift_reg[2] ),
    .ZN(_041_));
 AOI21_X1 _101_ (.A(_021_),
    .B1(_040_),
    .B2(_041_),
    .ZN(_010_));
 OAI21_X1 _102_ (.A(_014_),
    .B1(_015_),
    .B2(_020_),
    .ZN(_042_));
 INV_X1 _103_ (.A(_042_),
    .ZN(_011_));
 MUX2_X1 _104_ (.A(\pattern_reg[0] ),
    .B(net1),
    .S(_012_),
    .Z(_043_));
 OR2_X1 _105_ (.A1(_013_),
    .A2(_043_),
    .ZN(_004_));
 MUX2_X1 _106_ (.A(\pattern_reg[1] ),
    .B(net2),
    .S(_012_),
    .Z(_044_));
 OR2_X1 _107_ (.A1(_013_),
    .A2(_044_),
    .ZN(_005_));
 MUX2_X1 _108_ (.A(\pattern_reg[2] ),
    .B(net3),
    .S(_012_),
    .Z(_045_));
 AND2_X1 _109_ (.A1(net5),
    .A2(_045_),
    .ZN(_006_));
 MUX2_X1 _110_ (.A(\pattern_reg[3] ),
    .B(net4),
    .S(_012_),
    .Z(_046_));
 OR2_X1 _111_ (.A1(_013_),
    .A2(_046_),
    .ZN(_007_));
 HA_X1 _112_ (.A(\bit_count[0] ),
    .B(\bit_count[1] ),
    .CO(_058_),
    .S(_059_));
 HA_X1 _113_ (.A(_060_),
    .B(_061_),
    .CO(_062_),
    .S(_063_));
 DFF_X1 \bit_count[0]$_SDFFE_PP0P_  (.D(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\bit_count[0] ),
    .QN(_057_));
 DFF_X1 \bit_count[1]$_SDFFE_PP0P_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\bit_count[1] ),
    .QN(_056_));
 DFF_X1 \bit_count[2]$_SDFFE_PP0P_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\bit_count[2] ),
    .QN(_060_));
 DFF_X1 \pattern_detected$_SDFF_PP0_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net7),
    .QN(_055_));
 DFF_X1 \pattern_reg[0]$_SDFFE_PN1P_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\pattern_reg[0] ),
    .QN(_054_));
 DFF_X1 \pattern_reg[1]$_SDFFE_PN1P_  (.D(_005_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\pattern_reg[1] ),
    .QN(_053_));
 DFF_X1 \pattern_reg[2]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\pattern_reg[2] ),
    .QN(_052_));
 DFF_X1 \pattern_reg[3]$_SDFFE_PN1P_  (.D(_007_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\pattern_reg[3] ),
    .QN(_051_));
 DFF_X1 \shift_reg[0]$_SDFFE_PP0P_  (.D(_008_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\shift_reg[0] ),
    .QN(_050_));
 DFF_X1 \shift_reg[1]$_SDFFE_PP0P_  (.D(_009_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[1] ),
    .QN(_049_));
 DFF_X1 \shift_reg[2]$_SDFFE_PP0P_  (.D(_010_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\shift_reg[2] ),
    .QN(_048_));
 DFF_X1 \state$_SDFFE_PP0P_  (.D(_011_),
    .CK(clknet_1_0__leaf_clk),
    .Q(state),
    .QN(_047_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_111 ();
 BUF_X1 input1 (.A(config_pattern[0]),
    .Z(net1));
 BUF_X1 input2 (.A(config_pattern[1]),
    .Z(net2));
 BUF_X1 input3 (.A(config_pattern[2]),
    .Z(net3));
 BUF_X1 input4 (.A(config_pattern[3]),
    .Z(net4));
 BUF_X1 input5 (.A(rst_n),
    .Z(net5));
 BUF_X1 input6 (.A(serial_in),
    .Z(net6));
 BUF_X1 output7 (.A(net7),
    .Z(pattern_detected));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 INV_X1 clkload0 (.A(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X2 FILLER_0_417 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X2 FILLER_1_417 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X2 FILLER_2_417 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X2 FILLER_3_417 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X2 FILLER_4_417 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X2 FILLER_5_417 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X2 FILLER_6_417 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X2 FILLER_7_417 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X2 FILLER_8_417 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X2 FILLER_9_417 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X2 FILLER_10_417 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X2 FILLER_11_417 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X2 FILLER_12_417 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X2 FILLER_13_417 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X2 FILLER_14_417 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X2 FILLER_15_417 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X2 FILLER_16_417 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X2 FILLER_17_417 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X2 FILLER_18_417 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X2 FILLER_19_417 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X4 FILLER_20_193 ();
 FILLCELL_X2 FILLER_20_197 ();
 FILLCELL_X1 FILLER_20_199 ();
 FILLCELL_X32 FILLER_20_207 ();
 FILLCELL_X32 FILLER_20_239 ();
 FILLCELL_X32 FILLER_20_271 ();
 FILLCELL_X32 FILLER_20_303 ();
 FILLCELL_X32 FILLER_20_335 ();
 FILLCELL_X32 FILLER_20_367 ();
 FILLCELL_X16 FILLER_20_399 ();
 FILLCELL_X4 FILLER_20_415 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X2 FILLER_21_417 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X2 FILLER_22_417 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X2 FILLER_23_417 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X16 FILLER_24_161 ();
 FILLCELL_X8 FILLER_24_177 ();
 FILLCELL_X4 FILLER_24_185 ();
 FILLCELL_X2 FILLER_24_220 ();
 FILLCELL_X32 FILLER_24_224 ();
 FILLCELL_X32 FILLER_24_256 ();
 FILLCELL_X32 FILLER_24_288 ();
 FILLCELL_X32 FILLER_24_320 ();
 FILLCELL_X32 FILLER_24_352 ();
 FILLCELL_X32 FILLER_24_384 ();
 FILLCELL_X2 FILLER_24_416 ();
 FILLCELL_X1 FILLER_24_418 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X2 FILLER_25_161 ();
 FILLCELL_X1 FILLER_25_163 ();
 FILLCELL_X1 FILLER_25_183 ();
 FILLCELL_X1 FILLER_25_192 ();
 FILLCELL_X1 FILLER_25_224 ();
 FILLCELL_X32 FILLER_25_229 ();
 FILLCELL_X32 FILLER_25_261 ();
 FILLCELL_X32 FILLER_25_293 ();
 FILLCELL_X32 FILLER_25_325 ();
 FILLCELL_X32 FILLER_25_357 ();
 FILLCELL_X16 FILLER_25_389 ();
 FILLCELL_X8 FILLER_25_405 ();
 FILLCELL_X4 FILLER_25_413 ();
 FILLCELL_X2 FILLER_25_417 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X16 FILLER_26_161 ();
 FILLCELL_X8 FILLER_26_177 ();
 FILLCELL_X4 FILLER_26_185 ();
 FILLCELL_X1 FILLER_26_189 ();
 FILLCELL_X2 FILLER_26_198 ();
 FILLCELL_X1 FILLER_26_203 ();
 FILLCELL_X2 FILLER_26_219 ();
 FILLCELL_X32 FILLER_26_242 ();
 FILLCELL_X32 FILLER_26_274 ();
 FILLCELL_X32 FILLER_26_306 ();
 FILLCELL_X32 FILLER_26_338 ();
 FILLCELL_X32 FILLER_26_370 ();
 FILLCELL_X16 FILLER_26_402 ();
 FILLCELL_X1 FILLER_26_418 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X8 FILLER_27_193 ();
 FILLCELL_X4 FILLER_27_201 ();
 FILLCELL_X2 FILLER_27_205 ();
 FILLCELL_X1 FILLER_27_207 ();
 FILLCELL_X32 FILLER_27_211 ();
 FILLCELL_X32 FILLER_27_243 ();
 FILLCELL_X32 FILLER_27_275 ();
 FILLCELL_X32 FILLER_27_307 ();
 FILLCELL_X32 FILLER_27_339 ();
 FILLCELL_X32 FILLER_27_371 ();
 FILLCELL_X16 FILLER_27_403 ();
 FILLCELL_X16 FILLER_28_1 ();
 FILLCELL_X1 FILLER_28_17 ();
 FILLCELL_X4 FILLER_28_21 ();
 FILLCELL_X2 FILLER_28_25 ();
 FILLCELL_X1 FILLER_28_27 ();
 FILLCELL_X32 FILLER_28_31 ();
 FILLCELL_X32 FILLER_28_63 ();
 FILLCELL_X32 FILLER_28_95 ();
 FILLCELL_X16 FILLER_28_127 ();
 FILLCELL_X2 FILLER_28_143 ();
 FILLCELL_X32 FILLER_28_151 ();
 FILLCELL_X32 FILLER_28_183 ();
 FILLCELL_X2 FILLER_28_218 ();
 FILLCELL_X1 FILLER_28_220 ();
 FILLCELL_X32 FILLER_28_228 ();
 FILLCELL_X32 FILLER_28_260 ();
 FILLCELL_X32 FILLER_28_292 ();
 FILLCELL_X32 FILLER_28_324 ();
 FILLCELL_X32 FILLER_28_356 ();
 FILLCELL_X16 FILLER_28_388 ();
 FILLCELL_X8 FILLER_28_404 ();
 FILLCELL_X4 FILLER_28_412 ();
 FILLCELL_X2 FILLER_28_416 ();
 FILLCELL_X1 FILLER_28_418 ();
 FILLCELL_X16 FILLER_29_1 ();
 FILLCELL_X8 FILLER_29_17 ();
 FILLCELL_X2 FILLER_29_25 ();
 FILLCELL_X32 FILLER_29_30 ();
 FILLCELL_X32 FILLER_29_62 ();
 FILLCELL_X8 FILLER_29_94 ();
 FILLCELL_X4 FILLER_29_102 ();
 FILLCELL_X2 FILLER_29_106 ();
 FILLCELL_X1 FILLER_29_108 ();
 FILLCELL_X16 FILLER_29_113 ();
 FILLCELL_X8 FILLER_29_129 ();
 FILLCELL_X1 FILLER_29_137 ();
 FILLCELL_X16 FILLER_29_162 ();
 FILLCELL_X2 FILLER_29_178 ();
 FILLCELL_X8 FILLER_29_187 ();
 FILLCELL_X2 FILLER_29_195 ();
 FILLCELL_X2 FILLER_29_199 ();
 FILLCELL_X2 FILLER_29_206 ();
 FILLCELL_X32 FILLER_29_212 ();
 FILLCELL_X32 FILLER_29_244 ();
 FILLCELL_X32 FILLER_29_276 ();
 FILLCELL_X32 FILLER_29_308 ();
 FILLCELL_X32 FILLER_29_340 ();
 FILLCELL_X32 FILLER_29_372 ();
 FILLCELL_X8 FILLER_29_404 ();
 FILLCELL_X4 FILLER_29_412 ();
 FILLCELL_X2 FILLER_29_416 ();
 FILLCELL_X1 FILLER_29_418 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X16 FILLER_30_129 ();
 FILLCELL_X2 FILLER_30_145 ();
 FILLCELL_X1 FILLER_30_158 ();
 FILLCELL_X16 FILLER_30_176 ();
 FILLCELL_X4 FILLER_30_192 ();
 FILLCELL_X32 FILLER_30_212 ();
 FILLCELL_X32 FILLER_30_244 ();
 FILLCELL_X32 FILLER_30_276 ();
 FILLCELL_X32 FILLER_30_308 ();
 FILLCELL_X32 FILLER_30_340 ();
 FILLCELL_X32 FILLER_30_372 ();
 FILLCELL_X8 FILLER_30_404 ();
 FILLCELL_X4 FILLER_30_412 ();
 FILLCELL_X2 FILLER_30_416 ();
 FILLCELL_X1 FILLER_30_418 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X2 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_212 ();
 FILLCELL_X32 FILLER_31_244 ();
 FILLCELL_X32 FILLER_31_276 ();
 FILLCELL_X32 FILLER_31_308 ();
 FILLCELL_X32 FILLER_31_340 ();
 FILLCELL_X32 FILLER_31_372 ();
 FILLCELL_X8 FILLER_31_404 ();
 FILLCELL_X4 FILLER_31_412 ();
 FILLCELL_X2 FILLER_31_416 ();
 FILLCELL_X1 FILLER_31_418 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X8 FILLER_32_161 ();
 FILLCELL_X4 FILLER_32_169 ();
 FILLCELL_X1 FILLER_32_173 ();
 FILLCELL_X2 FILLER_32_179 ();
 FILLCELL_X1 FILLER_32_181 ();
 FILLCELL_X2 FILLER_32_203 ();
 FILLCELL_X1 FILLER_32_205 ();
 FILLCELL_X1 FILLER_32_214 ();
 FILLCELL_X8 FILLER_32_222 ();
 FILLCELL_X4 FILLER_32_230 ();
 FILLCELL_X1 FILLER_32_234 ();
 FILLCELL_X32 FILLER_32_252 ();
 FILLCELL_X32 FILLER_32_284 ();
 FILLCELL_X32 FILLER_32_316 ();
 FILLCELL_X32 FILLER_32_348 ();
 FILLCELL_X1 FILLER_32_380 ();
 FILLCELL_X32 FILLER_32_384 ();
 FILLCELL_X2 FILLER_32_416 ();
 FILLCELL_X1 FILLER_32_418 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X2 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_229 ();
 FILLCELL_X32 FILLER_33_261 ();
 FILLCELL_X32 FILLER_33_293 ();
 FILLCELL_X32 FILLER_33_325 ();
 FILLCELL_X32 FILLER_33_357 ();
 FILLCELL_X16 FILLER_33_389 ();
 FILLCELL_X8 FILLER_33_405 ();
 FILLCELL_X4 FILLER_33_413 ();
 FILLCELL_X2 FILLER_33_417 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X8 FILLER_34_161 ();
 FILLCELL_X4 FILLER_34_169 ();
 FILLCELL_X2 FILLER_34_173 ();
 FILLCELL_X1 FILLER_34_175 ();
 FILLCELL_X1 FILLER_34_199 ();
 FILLCELL_X32 FILLER_34_203 ();
 FILLCELL_X32 FILLER_34_235 ();
 FILLCELL_X32 FILLER_34_267 ();
 FILLCELL_X32 FILLER_34_299 ();
 FILLCELL_X32 FILLER_34_331 ();
 FILLCELL_X32 FILLER_34_363 ();
 FILLCELL_X16 FILLER_34_395 ();
 FILLCELL_X8 FILLER_34_411 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X8 FILLER_35_161 ();
 FILLCELL_X1 FILLER_35_169 ();
 FILLCELL_X8 FILLER_35_185 ();
 FILLCELL_X4 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_203 ();
 FILLCELL_X32 FILLER_35_235 ();
 FILLCELL_X32 FILLER_35_267 ();
 FILLCELL_X32 FILLER_35_299 ();
 FILLCELL_X32 FILLER_35_331 ();
 FILLCELL_X32 FILLER_35_363 ();
 FILLCELL_X16 FILLER_35_395 ();
 FILLCELL_X8 FILLER_35_411 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X4 FILLER_36_161 ();
 FILLCELL_X1 FILLER_36_165 ();
 FILLCELL_X32 FILLER_36_190 ();
 FILLCELL_X32 FILLER_36_222 ();
 FILLCELL_X32 FILLER_36_254 ();
 FILLCELL_X32 FILLER_36_286 ();
 FILLCELL_X32 FILLER_36_318 ();
 FILLCELL_X32 FILLER_36_350 ();
 FILLCELL_X32 FILLER_36_382 ();
 FILLCELL_X4 FILLER_36_414 ();
 FILLCELL_X1 FILLER_36_418 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X2 FILLER_37_417 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X2 FILLER_38_417 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X2 FILLER_39_417 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X2 FILLER_40_417 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X2 FILLER_41_417 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X2 FILLER_42_417 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X2 FILLER_43_417 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X2 FILLER_44_417 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X2 FILLER_45_417 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X2 FILLER_46_417 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X2 FILLER_47_417 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X2 FILLER_48_417 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X2 FILLER_49_417 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X2 FILLER_50_417 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X2 FILLER_51_417 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X2 FILLER_52_417 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X2 FILLER_53_417 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X16 FILLER_54_161 ();
 FILLCELL_X4 FILLER_54_177 ();
 FILLCELL_X16 FILLER_54_184 ();
 FILLCELL_X8 FILLER_54_200 ();
 FILLCELL_X4 FILLER_54_208 ();
 FILLCELL_X32 FILLER_54_215 ();
 FILLCELL_X32 FILLER_54_247 ();
 FILLCELL_X32 FILLER_54_279 ();
 FILLCELL_X32 FILLER_54_311 ();
 FILLCELL_X32 FILLER_54_343 ();
 FILLCELL_X32 FILLER_54_375 ();
 FILLCELL_X8 FILLER_54_407 ();
 FILLCELL_X4 FILLER_54_415 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X16 FILLER_55_161 ();
 FILLCELL_X4 FILLER_55_177 ();
 FILLCELL_X32 FILLER_55_184 ();
 FILLCELL_X32 FILLER_55_216 ();
 FILLCELL_X32 FILLER_55_248 ();
 FILLCELL_X32 FILLER_55_280 ();
 FILLCELL_X32 FILLER_55_312 ();
 FILLCELL_X32 FILLER_55_344 ();
 FILLCELL_X32 FILLER_55_376 ();
 FILLCELL_X8 FILLER_55_408 ();
 FILLCELL_X2 FILLER_55_416 ();
 FILLCELL_X1 FILLER_55_418 ();
endmodule
