module bsg_async_credit_counter (r_clk_i,
    r_credits_avail_o,
    r_dec_credit_i,
    r_infinite_credits_i,
    r_reset_i,
    w_clk_i,
    w_inc_token_i,
    w_reset_i);
 input r_clk_i;
 output r_credits_avail_o;
 input r_dec_credit_i;
 input r_infinite_credits_i;
 input r_reset_i;
 input w_clk_i;
 input w_inc_token_i;
 input w_reset_i;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire _37_;
 wire _38_;
 wire _39_;
 wire _40_;
 wire _41_;
 wire _42_;
 wire _43_;
 wire _44_;
 wire _45_;
 wire _46_;
 wire _47_;
 wire _48_;
 wire _49_;
 wire _50_;
 wire _51_;
 wire _52_;
 wire \bapg.w_ptr_binary_r_o[0] ;
 wire \bapg.w_ptr_binary_r_o[1] ;
 wire \bapg.w_ptr_binary_r_o[2] ;
 wire \bapg.w_ptr_gray_r[0] ;
 wire \bapg.w_ptr_gray_r[1] ;
 wire \bapg.w_ptr_gray_r_rsync_o[0] ;
 wire \bapg.w_ptr_gray_r_rsync_o[1] ;
 wire \bapg.w_ptr_gray_r_rsync_o[2] ;
 wire \bapg.w_ptr_gray_r_rsync_r[0][0] ;
 wire \bapg.w_ptr_gray_r_rsync_r[0][1] ;
 wire \bapg.w_ptr_gray_r_rsync_r[0][2] ;
 wire \bapg.w_ptr_n[0] ;
 wire \bapg.w_ptr_n[1] ;
 wire \r_counter_r[0] ;
 wire \r_counter_r[1] ;
 wire \r_counter_r[2] ;
 wire \r_counter_r_hi_bits_gray[0] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_0_w_clk_i;
 wire clknet_1_0__leaf_w_clk_i;
 wire clknet_1_1__leaf_w_clk_i;

 BUF_X4 _53_ (.A(w_reset_i),
    .Z(_09_));
 BUF_X4 _54_ (.A(net5),
    .Z(_10_));
 NOR2_X1 _55_ (.A1(\bapg.w_ptr_gray_r[0] ),
    .A2(_10_),
    .ZN(_11_));
 INV_X2 _56_ (.A(_10_),
    .ZN(_12_));
 XOR2_X1 _57_ (.A(\bapg.w_ptr_n[0] ),
    .B(\bapg.w_ptr_n[1] ),
    .Z(_13_));
 NOR2_X1 _58_ (.A1(_12_),
    .A2(_13_),
    .ZN(_14_));
 NOR3_X1 _59_ (.A1(_09_),
    .A2(_11_),
    .A3(_14_),
    .ZN(_01_));
 INV_X1 _60_ (.A(_09_),
    .ZN(_15_));
 XNOR2_X1 _61_ (.A(\bapg.w_ptr_n[1] ),
    .B(_51_),
    .ZN(_16_));
 NAND4_X1 _62_ (.A1(_10_),
    .A2(\bapg.w_ptr_binary_r_o[2] ),
    .A3(_15_),
    .A4(_16_),
    .ZN(_17_));
 OR3_X1 _63_ (.A1(_12_),
    .A2(\bapg.w_ptr_binary_r_o[2] ),
    .A3(_09_),
    .ZN(_18_));
 NAND2_X1 _64_ (.A1(_12_),
    .A2(\bapg.w_ptr_gray_r[1] ),
    .ZN(_19_));
 OAI221_X1 _65_ (.A(_17_),
    .B1(_18_),
    .B2(_16_),
    .C1(_09_),
    .C2(_19_),
    .ZN(_02_));
 NAND2_X1 _66_ (.A1(_10_),
    .A2(_51_),
    .ZN(_20_));
 XOR2_X1 _67_ (.A(\bapg.w_ptr_binary_r_o[2] ),
    .B(_20_),
    .Z(_21_));
 NOR2_X1 _68_ (.A1(_09_),
    .A2(_21_),
    .ZN(_03_));
 NAND2_X1 _69_ (.A1(_10_),
    .A2(\bapg.w_ptr_n[0] ),
    .ZN(_22_));
 NAND2_X1 _70_ (.A1(_12_),
    .A2(\bapg.w_ptr_binary_r_o[0] ),
    .ZN(_23_));
 AOI21_X1 _71_ (.A(_09_),
    .B1(_22_),
    .B2(_23_),
    .ZN(_04_));
 NAND2_X1 _72_ (.A1(_10_),
    .A2(\bapg.w_ptr_n[1] ),
    .ZN(_24_));
 NAND2_X1 _73_ (.A1(_12_),
    .A2(\bapg.w_ptr_binary_r_o[1] ),
    .ZN(_25_));
 AOI21_X1 _74_ (.A(_09_),
    .B1(_24_),
    .B2(_25_),
    .ZN(_05_));
 MUX2_X1 _75_ (.A(\r_counter_r[0] ),
    .B(_00_),
    .S(net2),
    .Z(_26_));
 INV_X1 _76_ (.A(_26_),
    .ZN(_27_));
 NOR2_X1 _77_ (.A1(net4),
    .A2(_27_),
    .ZN(_06_));
 MUX2_X1 _78_ (.A(\r_counter_r[1] ),
    .B(\r_counter_r_hi_bits_gray[0] ),
    .S(net2),
    .Z(_28_));
 INV_X1 _79_ (.A(_28_),
    .ZN(_29_));
 NOR2_X1 _80_ (.A1(net4),
    .A2(_29_),
    .ZN(_07_));
 NAND2_X1 _81_ (.A1(_52_),
    .A2(net2),
    .ZN(_30_));
 XNOR2_X1 _82_ (.A(\r_counter_r[2] ),
    .B(_30_),
    .ZN(_31_));
 OR2_X1 _83_ (.A1(net4),
    .A2(_31_),
    .ZN(_08_));
 XOR2_X1 _84_ (.A(\r_counter_r_hi_bits_gray[0] ),
    .B(\bapg.w_ptr_gray_r_rsync_o[0] ),
    .Z(_32_));
 NOR2_X1 _85_ (.A1(net3),
    .A2(_32_),
    .ZN(_33_));
 XOR2_X1 _86_ (.A(\r_counter_r[1] ),
    .B(\bapg.w_ptr_gray_r_rsync_o[1] ),
    .Z(_34_));
 NOR3_X1 _87_ (.A1(\r_counter_r[2] ),
    .A2(\bapg.w_ptr_gray_r_rsync_o[2] ),
    .A3(_34_),
    .ZN(_35_));
 AND3_X1 _88_ (.A1(\r_counter_r[2] ),
    .A2(\bapg.w_ptr_gray_r_rsync_o[2] ),
    .A3(_34_),
    .ZN(_36_));
 OAI21_X1 _89_ (.A(_33_),
    .B1(_35_),
    .B2(_36_),
    .ZN(net6));
 HA_X1 _90_ (.A(net5),
    .B(\bapg.w_ptr_binary_r_o[0] ),
    .CO(_50_),
    .S(\bapg.w_ptr_n[0] ));
 HA_X1 _91_ (.A(\bapg.w_ptr_binary_r_o[1] ),
    .B(_50_),
    .CO(_51_),
    .S(\bapg.w_ptr_n[1] ));
 HA_X1 _92_ (.A(\r_counter_r[0] ),
    .B(\r_counter_r[1] ),
    .CO(_52_),
    .S(\r_counter_r_hi_bits_gray[0] ));
 DFF_X1 \bapg.w_ptr_gray_r[0]$_SDFFE_PP0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_w_clk_i),
    .Q(\bapg.w_ptr_gray_r[0] ),
    .QN(_43_));
 DFF_X1 \bapg.w_ptr_gray_r[1]$_SDFFE_PP0P_  (.D(_02_),
    .CK(clknet_1_1__leaf_w_clk_i),
    .Q(\bapg.w_ptr_gray_r[1] ),
    .QN(_42_));
 DFF_X1 \bapg.w_ptr_gray_r[2]$_SDFFE_PP0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_w_clk_i),
    .Q(\bapg.w_ptr_binary_r_o[2] ),
    .QN(_44_));
 DFF_X1 \bapg.w_ptr_gray_r_rsync_r[0][0]$_DFF_P_  (.D(\bapg.w_ptr_gray_r[0] ),
    .CK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_r[0][0] ),
    .QN(_45_));
 DFF_X1 \bapg.w_ptr_gray_r_rsync_r[0][1]$_DFF_P_  (.D(\bapg.w_ptr_gray_r[1] ),
    .CK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_r[0][1] ),
    .QN(_46_));
 DFF_X1 \bapg.w_ptr_gray_r_rsync_r[0][2]$_DFF_P_  (.D(\bapg.w_ptr_binary_r_o[2] ),
    .CK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_r[0][2] ),
    .QN(_47_));
 DFF_X1 \bapg.w_ptr_gray_r_rsync_r[1][0]$_DFF_P_  (.D(\bapg.w_ptr_gray_r_rsync_r[0][0] ),
    .CK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_o[0] ),
    .QN(_48_));
 DFF_X1 \bapg.w_ptr_gray_r_rsync_r[1][1]$_DFF_P_  (.D(\bapg.w_ptr_gray_r_rsync_r[0][1] ),
    .CK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_o[1] ),
    .QN(_49_));
 DFF_X1 \bapg.w_ptr_gray_r_rsync_r[1][2]$_DFF_P_  (.D(\bapg.w_ptr_gray_r_rsync_r[0][2] ),
    .CK(net1),
    .Q(\bapg.w_ptr_gray_r_rsync_o[2] ),
    .QN(_41_));
 DFF_X1 \bapg.w_ptr_r[0]$_SDFFE_PP0P_  (.D(_04_),
    .CK(clknet_1_0__leaf_w_clk_i),
    .Q(\bapg.w_ptr_binary_r_o[0] ),
    .QN(_40_));
 DFF_X1 \bapg.w_ptr_r[1]$_SDFFE_PP0P_  (.D(_05_),
    .CK(clknet_1_0__leaf_w_clk_i),
    .Q(\bapg.w_ptr_binary_r_o[1] ),
    .QN(_39_));
 DFF_X1 \r_counter_r[0]$_SDFFE_PP0P_  (.D(_06_),
    .CK(net1),
    .Q(\r_counter_r[0] ),
    .QN(_00_));
 DFF_X1 \r_counter_r[1]$_SDFFE_PP0P_  (.D(_07_),
    .CK(net1),
    .Q(\r_counter_r[1] ),
    .QN(_38_));
 DFF_X1 \r_counter_r[2]$_SDFFE_PP1P_  (.D(_08_),
    .CK(net1),
    .Q(\r_counter_r[2] ),
    .QN(_37_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_47 ();
 CLKBUF_X2 input1 (.A(r_clk_i),
    .Z(net1));
 BUF_X1 input2 (.A(r_dec_credit_i),
    .Z(net2));
 BUF_X1 input3 (.A(r_infinite_credits_i),
    .Z(net3));
 BUF_X1 input4 (.A(r_reset_i),
    .Z(net4));
 BUF_X1 input5 (.A(w_inc_token_i),
    .Z(net5));
 BUF_X1 output6 (.A(net6),
    .Z(r_credits_avail_o));
 CLKBUF_X3 clkbuf_0_w_clk_i (.A(w_clk_i),
    .Z(clknet_0_w_clk_i));
 CLKBUF_X3 clkbuf_1_0__f_w_clk_i (.A(clknet_0_w_clk_i),
    .Z(clknet_1_0__leaf_w_clk_i));
 CLKBUF_X3 clkbuf_1_1__f_w_clk_i (.A(clknet_0_w_clk_i),
    .Z(clknet_1_1__leaf_w_clk_i));
 CLKBUF_X1 clkload0 (.A(clknet_1_1__leaf_w_clk_i));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_68 ();
 FILLCELL_X32 FILLER_0_100 ();
 FILLCELL_X32 FILLER_0_132 ();
 FILLCELL_X8 FILLER_0_164 ();
 FILLCELL_X4 FILLER_0_172 ();
 FILLCELL_X1 FILLER_0_176 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X16 FILLER_1_161 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X16 FILLER_2_161 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X16 FILLER_3_161 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X16 FILLER_4_161 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X16 FILLER_5_161 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X16 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_49 ();
 FILLCELL_X2 FILLER_6_57 ();
 FILLCELL_X1 FILLER_6_59 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X16 FILLER_6_161 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X8 FILLER_7_33 ();
 FILLCELL_X2 FILLER_7_75 ();
 FILLCELL_X1 FILLER_7_77 ();
 FILLCELL_X32 FILLER_7_95 ();
 FILLCELL_X16 FILLER_7_127 ();
 FILLCELL_X8 FILLER_7_143 ();
 FILLCELL_X4 FILLER_7_151 ();
 FILLCELL_X2 FILLER_7_155 ();
 FILLCELL_X1 FILLER_7_157 ();
 FILLCELL_X8 FILLER_7_167 ();
 FILLCELL_X2 FILLER_7_175 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X16 FILLER_8_33 ();
 FILLCELL_X4 FILLER_8_49 ();
 FILLCELL_X1 FILLER_8_53 ();
 FILLCELL_X1 FILLER_8_61 ();
 FILLCELL_X2 FILLER_8_71 ();
 FILLCELL_X1 FILLER_8_73 ();
 FILLCELL_X2 FILLER_8_77 ();
 FILLCELL_X1 FILLER_8_79 ();
 FILLCELL_X1 FILLER_8_84 ();
 FILLCELL_X8 FILLER_8_88 ();
 FILLCELL_X4 FILLER_8_96 ();
 FILLCELL_X2 FILLER_8_100 ();
 FILLCELL_X16 FILLER_8_119 ();
 FILLCELL_X2 FILLER_8_135 ();
 FILLCELL_X4 FILLER_8_171 ();
 FILLCELL_X2 FILLER_8_175 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X8 FILLER_9_49 ();
 FILLCELL_X1 FILLER_9_61 ();
 FILLCELL_X4 FILLER_9_75 ();
 FILLCELL_X2 FILLER_9_79 ();
 FILLCELL_X1 FILLER_9_81 ();
 FILLCELL_X32 FILLER_9_85 ();
 FILLCELL_X2 FILLER_9_117 ();
 FILLCELL_X1 FILLER_9_119 ();
 FILLCELL_X8 FILLER_9_137 ();
 FILLCELL_X1 FILLER_9_145 ();
 FILLCELL_X2 FILLER_9_169 ();
 FILLCELL_X1 FILLER_9_171 ();
 FILLCELL_X1 FILLER_9_176 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X8 FILLER_10_33 ();
 FILLCELL_X4 FILLER_10_41 ();
 FILLCELL_X2 FILLER_10_45 ();
 FILLCELL_X1 FILLER_10_67 ();
 FILLCELL_X32 FILLER_10_74 ();
 FILLCELL_X32 FILLER_10_106 ();
 FILLCELL_X4 FILLER_10_138 ();
 FILLCELL_X2 FILLER_10_142 ();
 FILLCELL_X1 FILLER_10_144 ();
 FILLCELL_X2 FILLER_10_156 ();
 FILLCELL_X4 FILLER_10_161 ();
 FILLCELL_X8 FILLER_10_168 ();
 FILLCELL_X1 FILLER_10_176 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X2 FILLER_11_65 ();
 FILLCELL_X1 FILLER_11_67 ();
 FILLCELL_X32 FILLER_11_78 ();
 FILLCELL_X32 FILLER_11_110 ();
 FILLCELL_X8 FILLER_11_142 ();
 FILLCELL_X2 FILLER_11_150 ();
 FILLCELL_X8 FILLER_11_162 ();
 FILLCELL_X4 FILLER_11_170 ();
 FILLCELL_X2 FILLER_11_174 ();
 FILLCELL_X1 FILLER_11_176 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_33 ();
 FILLCELL_X8 FILLER_12_49 ();
 FILLCELL_X2 FILLER_12_57 ();
 FILLCELL_X2 FILLER_12_84 ();
 FILLCELL_X32 FILLER_12_89 ();
 FILLCELL_X8 FILLER_12_121 ();
 FILLCELL_X4 FILLER_12_129 ();
 FILLCELL_X2 FILLER_12_133 ();
 FILLCELL_X1 FILLER_12_135 ();
 FILLCELL_X4 FILLER_12_153 ();
 FILLCELL_X4 FILLER_12_160 ();
 FILLCELL_X1 FILLER_12_164 ();
 FILLCELL_X8 FILLER_12_168 ();
 FILLCELL_X1 FILLER_12_176 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X16 FILLER_13_33 ();
 FILLCELL_X4 FILLER_13_49 ();
 FILLCELL_X2 FILLER_13_53 ();
 FILLCELL_X1 FILLER_13_55 ();
 FILLCELL_X4 FILLER_13_73 ();
 FILLCELL_X1 FILLER_13_77 ();
 FILLCELL_X4 FILLER_13_95 ();
 FILLCELL_X2 FILLER_13_99 ();
 FILLCELL_X1 FILLER_13_101 ();
 FILLCELL_X1 FILLER_13_119 ();
 FILLCELL_X4 FILLER_13_137 ();
 FILLCELL_X2 FILLER_13_141 ();
 FILLCELL_X1 FILLER_13_143 ();
 FILLCELL_X2 FILLER_13_150 ();
 FILLCELL_X4 FILLER_13_160 ();
 FILLCELL_X2 FILLER_13_164 ();
 FILLCELL_X1 FILLER_13_166 ();
 FILLCELL_X4 FILLER_13_170 ();
 FILLCELL_X2 FILLER_13_174 ();
 FILLCELL_X1 FILLER_13_176 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_33 ();
 FILLCELL_X1 FILLER_14_35 ();
 FILLCELL_X32 FILLER_14_43 ();
 FILLCELL_X2 FILLER_14_75 ();
 FILLCELL_X16 FILLER_14_85 ();
 FILLCELL_X4 FILLER_14_101 ();
 FILLCELL_X4 FILLER_14_122 ();
 FILLCELL_X2 FILLER_14_126 ();
 FILLCELL_X4 FILLER_14_145 ();
 FILLCELL_X2 FILLER_14_149 ();
 FILLCELL_X16 FILLER_14_156 ();
 FILLCELL_X4 FILLER_14_172 ();
 FILLCELL_X1 FILLER_14_176 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X16 FILLER_15_161 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X16 FILLER_16_161 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X16 FILLER_17_161 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X16 FILLER_18_161 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X16 FILLER_19_161 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X16 FILLER_20_161 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X16 FILLER_21_161 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X16 FILLER_22_161 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X16 FILLER_23_161 ();
endmodule
