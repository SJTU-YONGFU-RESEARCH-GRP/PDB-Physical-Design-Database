module fifo (clk,
    empty,
    full,
    rd_en,
    rst_n,
    wr_en,
    din,
    dout);
 input clk;
 output empty;
 output full;
 input rd_en;
 input rst_n;
 input wr_en;
 input [7:0] din;
 output [7:0] dout;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net23;
 wire net24;

 sky130_fd_sc_hd__xnor2_1 _261_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .Y(_038_));
 sky130_fd_sc_hd__xnor2_1 _262_ (.A(\rd_ptr[1] ),
    .B(\wr_ptr[1] ),
    .Y(_039_));
 sky130_fd_sc_hd__xnor2_1 _263_ (.A(\rd_ptr[0] ),
    .B(\wr_ptr[0] ),
    .Y(_040_));
 sky130_fd_sc_hd__buf_4 _264_ (.A(\rd_ptr[3] ),
    .X(_041_));
 sky130_fd_sc_hd__clkbuf_4 _265_ (.A(\wr_ptr[3] ),
    .X(_042_));
 sky130_fd_sc_hd__xnor2_1 _266_ (.A(_041_),
    .B(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__clkbuf_4 _267_ (.A(\wr_ptr[2] ),
    .X(_044_));
 sky130_fd_sc_hd__xnor2_1 _268_ (.A(_044_),
    .B(\rd_ptr[2] ),
    .Y(_045_));
 sky130_fd_sc_hd__nand4_2 _269_ (.A(_039_),
    .B(_040_),
    .C(_043_),
    .D(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_1 _270_ (.A(_038_),
    .B(_046_),
    .Y(net22));
 sky130_fd_sc_hd__nand2_8 _271_ (.A(net11),
    .B(_254_),
    .Y(_047_));
 sky130_fd_sc_hd__o21a_1 _272_ (.A1(_038_),
    .A2(_046_),
    .B1(net12),
    .X(_048_));
 sky130_fd_sc_hd__buf_4 _273_ (.A(_048_),
    .X(_049_));
 sky130_fd_sc_hd__nor2_1 _274_ (.A(_044_),
    .B(_042_),
    .Y(_050_));
 sky130_fd_sc_hd__nand2_4 _275_ (.A(_049_),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_4 _276_ (.A(_047_),
    .B(_051_),
    .Y(_015_));
 sky130_fd_sc_hd__nand2_4 _277_ (.A(net11),
    .B(_257_),
    .Y(_052_));
 sky130_fd_sc_hd__nor2_4 _278_ (.A(_051_),
    .B(_052_),
    .Y(_014_));
 sky130_fd_sc_hd__nand2_4 _279_ (.A(net11),
    .B(_255_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_4 _280_ (.A(_051_),
    .B(_053_),
    .Y(_013_));
 sky130_fd_sc_hd__nand2_8 _281_ (.A(net11),
    .B(_259_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_8 _282_ (.A(_051_),
    .B(_054_),
    .Y(_012_));
 sky130_fd_sc_hd__nand3b_4 _283_ (.A_N(_042_),
    .B(_049_),
    .C(_044_),
    .Y(_055_));
 sky130_fd_sc_hd__nor2_8 _284_ (.A(_047_),
    .B(_055_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_4 _285_ (.A(_052_),
    .B(_055_),
    .Y(_010_));
 sky130_fd_sc_hd__nor2_4 _286_ (.A(_053_),
    .B(_055_),
    .Y(_009_));
 sky130_fd_sc_hd__nor2_4 _287_ (.A(_054_),
    .B(_055_),
    .Y(_008_));
 sky130_fd_sc_hd__nand3b_4 _288_ (.A_N(_044_),
    .B(_042_),
    .C(_049_),
    .Y(_056_));
 sky130_fd_sc_hd__nor2_8 _289_ (.A(_047_),
    .B(_056_),
    .Y(_007_));
 sky130_fd_sc_hd__nor2_8 _290_ (.A(_052_),
    .B(_056_),
    .Y(_006_));
 sky130_fd_sc_hd__nor2_8 _291_ (.A(_053_),
    .B(_056_),
    .Y(_005_));
 sky130_fd_sc_hd__nor2_8 _292_ (.A(_054_),
    .B(_056_),
    .Y(_004_));
 sky130_fd_sc_hd__nand3_4 _293_ (.A(_044_),
    .B(_042_),
    .C(_049_),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_8 _294_ (.A(_047_),
    .B(_057_),
    .Y(_003_));
 sky130_fd_sc_hd__nor2_4 _295_ (.A(_052_),
    .B(_057_),
    .Y(_002_));
 sky130_fd_sc_hd__nor2_4 _296_ (.A(_053_),
    .B(_057_),
    .Y(_001_));
 sky130_fd_sc_hd__nor2_4 _297_ (.A(_054_),
    .B(_057_),
    .Y(_000_));
 sky130_fd_sc_hd__xor2_1 _298_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .X(_058_));
 sky130_fd_sc_hd__nor2_1 _299_ (.A(_058_),
    .B(_046_),
    .Y(net21));
 sky130_fd_sc_hd__inv_1 _300_ (.A(\rd_ptr[0] ),
    .Y(_018_));
 sky130_fd_sc_hd__inv_1 _301_ (.A(\wr_ptr[0] ),
    .Y(_016_));
 sky130_fd_sc_hd__inv_1 _302_ (.A(\rd_ptr[1] ),
    .Y(_245_));
 sky130_fd_sc_hd__inv_1 _303_ (.A(\wr_ptr[1] ),
    .Y(_253_));
 sky130_fd_sc_hd__o21ai_1 _304_ (.A1(_058_),
    .A2(_046_),
    .B1(net10),
    .Y(_059_));
 sky130_fd_sc_hd__clkbuf_4 _305_ (.A(_059_),
    .X(_060_));
 sky130_fd_sc_hd__buf_4 _306_ (.A(\rd_ptr[2] ),
    .X(_061_));
 sky130_fd_sc_hd__buf_4 _307_ (.A(_061_),
    .X(_062_));
 sky130_fd_sc_hd__buf_4 _308_ (.A(_062_),
    .X(_063_));
 sky130_fd_sc_hd__buf_6 _309_ (.A(_041_),
    .X(_064_));
 sky130_fd_sc_hd__buf_4 _310_ (.A(_064_),
    .X(_065_));
 sky130_fd_sc_hd__clkbuf_4 _311_ (.A(_251_),
    .X(_066_));
 sky130_fd_sc_hd__clkbuf_4 _312_ (.A(_247_),
    .X(_067_));
 sky130_fd_sc_hd__a22oi_1 _313_ (.A1(_066_),
    .A2(\mem[7][0] ),
    .B1(\mem[6][0] ),
    .B2(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__buf_2 _314_ (.A(_249_),
    .X(_069_));
 sky130_fd_sc_hd__clkbuf_4 _315_ (.A(_069_),
    .X(_070_));
 sky130_fd_sc_hd__nand3_1 _316_ (.A(_065_),
    .B(\mem[13][0] ),
    .C(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__o21ai_0 _317_ (.A1(_065_),
    .A2(_068_),
    .B1(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__buf_6 _318_ (.A(_247_),
    .X(_073_));
 sky130_fd_sc_hd__clkbuf_4 _319_ (.A(_069_),
    .X(_074_));
 sky130_fd_sc_hd__a22oi_1 _320_ (.A1(\mem[10][0] ),
    .A2(_073_),
    .B1(_074_),
    .B2(\mem[9][0] ),
    .Y(_075_));
 sky130_fd_sc_hd__a221oi_1 _321_ (.A1(_066_),
    .A2(\mem[3][0] ),
    .B1(\mem[2][0] ),
    .B2(_073_),
    .C1(_064_),
    .Y(_076_));
 sky130_fd_sc_hd__a211oi_1 _322_ (.A1(_065_),
    .A2(_075_),
    .B1(_076_),
    .C1(_062_),
    .Y(_077_));
 sky130_fd_sc_hd__a21oi_1 _323_ (.A1(_063_),
    .A2(_072_),
    .B1(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__clkbuf_4 _324_ (.A(_246_),
    .X(_079_));
 sky130_fd_sc_hd__mux2_1 _325_ (.A0(\mem[4][0] ),
    .A1(\mem[12][0] ),
    .S(_041_),
    .X(_080_));
 sky130_fd_sc_hd__o21ai_0 _326_ (.A1(_061_),
    .A2(_041_),
    .B1(_246_),
    .Y(_081_));
 sky130_fd_sc_hd__nor3_1 _327_ (.A(_251_),
    .B(_247_),
    .C(_069_),
    .Y(_082_));
 sky130_fd_sc_hd__and2_0 _328_ (.A(_081_),
    .B(_082_),
    .X(_083_));
 sky130_fd_sc_hd__clkbuf_8 _329_ (.A(_064_),
    .X(_084_));
 sky130_fd_sc_hd__clkbuf_4 _330_ (.A(_066_),
    .X(_085_));
 sky130_fd_sc_hd__nand2_1 _331_ (.A(_084_),
    .B(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__mux2i_1 _332_ (.A0(\mem[11][0] ),
    .A1(\mem[15][0] ),
    .S(_062_),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_1 _333_ (.A(_086_),
    .B(_087_),
    .Y(_088_));
 sky130_fd_sc_hd__a311oi_1 _334_ (.A1(_063_),
    .A2(_079_),
    .A3(_080_),
    .B1(_083_),
    .C1(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__nand2_1 _335_ (.A(\mem[1][0] ),
    .B(_070_),
    .Y(_090_));
 sky130_fd_sc_hd__nand3_1 _336_ (.A(_084_),
    .B(\mem[8][0] ),
    .C(_079_),
    .Y(_091_));
 sky130_fd_sc_hd__o21ai_0 _337_ (.A1(_084_),
    .A2(_090_),
    .B1(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__nand2_1 _338_ (.A(\mem[5][0] ),
    .B(_070_),
    .Y(_093_));
 sky130_fd_sc_hd__nand3_1 _339_ (.A(_084_),
    .B(\mem[14][0] ),
    .C(_067_),
    .Y(_094_));
 sky130_fd_sc_hd__o211ai_1 _340_ (.A1(_065_),
    .A2(_093_),
    .B1(_094_),
    .C1(_063_),
    .Y(_095_));
 sky130_fd_sc_hd__o21ai_1 _341_ (.A1(_063_),
    .A2(_092_),
    .B1(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__nand2_2 _342_ (.A(_081_),
    .B(_082_),
    .Y(_097_));
 sky130_fd_sc_hd__clkbuf_4 _343_ (.A(_097_),
    .X(_098_));
 sky130_fd_sc_hd__nor2_1 _344_ (.A(\mem[0][0] ),
    .B(_098_),
    .Y(_099_));
 sky130_fd_sc_hd__a31o_1 _345_ (.A1(_078_),
    .A2(_089_),
    .A3(_096_),
    .B1(_099_),
    .X(_100_));
 sky130_fd_sc_hd__nand2_1 _346_ (.A(net13),
    .B(_060_),
    .Y(_101_));
 sky130_fd_sc_hd__o21ai_0 _347_ (.A1(_060_),
    .A2(_100_),
    .B1(_101_),
    .Y(_020_));
 sky130_fd_sc_hd__buf_4 _348_ (.A(_059_),
    .X(_102_));
 sky130_fd_sc_hd__clkinv_4 _349_ (.A(_061_),
    .Y(_103_));
 sky130_fd_sc_hd__clkbuf_4 _350_ (.A(_064_),
    .X(_104_));
 sky130_fd_sc_hd__a22oi_1 _351_ (.A1(_085_),
    .A2(\mem[3][1] ),
    .B1(\mem[1][1] ),
    .B2(_070_),
    .Y(_105_));
 sky130_fd_sc_hd__clkbuf_4 _352_ (.A(_073_),
    .X(_106_));
 sky130_fd_sc_hd__nand3_1 _353_ (.A(_104_),
    .B(\mem[10][1] ),
    .C(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__o21ai_0 _354_ (.A1(_104_),
    .A2(_105_),
    .B1(_107_),
    .Y(_108_));
 sky130_fd_sc_hd__a22oi_1 _355_ (.A1(\mem[4][1] ),
    .A2(_079_),
    .B1(_106_),
    .B2(\mem[6][1] ),
    .Y(_109_));
 sky130_fd_sc_hd__nand2b_2 _356_ (.A_N(_041_),
    .B(_061_),
    .Y(_110_));
 sky130_fd_sc_hd__nor2_1 _357_ (.A(_109_),
    .B(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__a21oi_1 _358_ (.A1(_103_),
    .A2(_108_),
    .B1(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__nand2b_2 _359_ (.A_N(_061_),
    .B(_041_),
    .Y(_113_));
 sky130_fd_sc_hd__a22oi_1 _360_ (.A1(_085_),
    .A2(\mem[11][1] ),
    .B1(\mem[8][1] ),
    .B2(_079_),
    .Y(_114_));
 sky130_fd_sc_hd__nor2_1 _361_ (.A(_113_),
    .B(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__buf_6 _362_ (.A(_064_),
    .X(_116_));
 sky130_fd_sc_hd__nand2_1 _363_ (.A(_062_),
    .B(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__a22oi_1 _364_ (.A1(\mem[12][1] ),
    .A2(_079_),
    .B1(_106_),
    .B2(\mem[14][1] ),
    .Y(_118_));
 sky130_fd_sc_hd__nand2_2 _365_ (.A(_061_),
    .B(_066_),
    .Y(_119_));
 sky130_fd_sc_hd__mux2i_1 _366_ (.A0(\mem[7][1] ),
    .A1(\mem[15][1] ),
    .S(_084_),
    .Y(_120_));
 sky130_fd_sc_hd__o22ai_1 _367_ (.A1(_117_),
    .A2(_118_),
    .B1(_119_),
    .B2(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__nor3_1 _368_ (.A(_083_),
    .B(_115_),
    .C(_121_),
    .Y(_122_));
 sky130_fd_sc_hd__inv_1 _369_ (.A(\mem[5][1] ),
    .Y(_123_));
 sky130_fd_sc_hd__inv_1 _370_ (.A(\mem[9][1] ),
    .Y(_124_));
 sky130_fd_sc_hd__o22ai_1 _371_ (.A1(_123_),
    .A2(_110_),
    .B1(_113_),
    .B2(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__nand2_1 _372_ (.A(_070_),
    .B(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_1 _373_ (.A(_062_),
    .B(_116_),
    .Y(_127_));
 sky130_fd_sc_hd__and3_1 _374_ (.A(_061_),
    .B(_041_),
    .C(_069_),
    .X(_128_));
 sky130_fd_sc_hd__a32oi_1 _375_ (.A1(\mem[2][1] ),
    .A2(_106_),
    .A3(_127_),
    .B1(_128_),
    .B2(\mem[13][1] ),
    .Y(_129_));
 sky130_fd_sc_hd__nand4_1 _376_ (.A(_112_),
    .B(_122_),
    .C(_126_),
    .D(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__nor2_1 _377_ (.A(\mem[0][1] ),
    .B(_098_),
    .Y(_131_));
 sky130_fd_sc_hd__nor2_1 _378_ (.A(_102_),
    .B(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__a22o_1 _379_ (.A1(net14),
    .A2(_102_),
    .B1(_130_),
    .B2(_132_),
    .X(_021_));
 sky130_fd_sc_hd__clkbuf_4 _380_ (.A(_246_),
    .X(_133_));
 sky130_fd_sc_hd__a222oi_1 _381_ (.A1(\mem[6][2] ),
    .A2(_073_),
    .B1(_069_),
    .B2(\mem[5][2] ),
    .C1(\mem[4][2] ),
    .C2(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__a222oi_1 _382_ (.A1(\mem[14][2] ),
    .A2(_073_),
    .B1(_069_),
    .B2(\mem[13][2] ),
    .C1(\mem[12][2] ),
    .C2(_133_),
    .Y(_135_));
 sky130_fd_sc_hd__mux2i_1 _383_ (.A0(_134_),
    .A1(_135_),
    .S(_084_),
    .Y(_136_));
 sky130_fd_sc_hd__a22oi_2 _384_ (.A1(\mem[8][2] ),
    .A2(_133_),
    .B1(_074_),
    .B2(\mem[9][2] ),
    .Y(_137_));
 sky130_fd_sc_hd__nand2_1 _385_ (.A(_085_),
    .B(\mem[11][2] ),
    .Y(_138_));
 sky130_fd_sc_hd__a21oi_1 _386_ (.A1(\mem[2][2] ),
    .A2(_067_),
    .B1(_116_),
    .Y(_139_));
 sky130_fd_sc_hd__a311oi_4 _387_ (.A1(_065_),
    .A2(_137_),
    .A3(_138_),
    .B1(_139_),
    .C1(_062_),
    .Y(_140_));
 sky130_fd_sc_hd__mux2i_1 _388_ (.A0(\mem[7][2] ),
    .A1(\mem[15][2] ),
    .S(_064_),
    .Y(_141_));
 sky130_fd_sc_hd__o21ai_0 _389_ (.A1(_119_),
    .A2(_141_),
    .B1(_097_),
    .Y(_142_));
 sky130_fd_sc_hd__a22oi_1 _390_ (.A1(_066_),
    .A2(\mem[3][2] ),
    .B1(\mem[1][2] ),
    .B2(_074_),
    .Y(_143_));
 sky130_fd_sc_hd__nand3_1 _391_ (.A(_116_),
    .B(\mem[10][2] ),
    .C(_067_),
    .Y(_144_));
 sky130_fd_sc_hd__o21a_1 _392_ (.A1(_084_),
    .A2(_143_),
    .B1(_144_),
    .X(_145_));
 sky130_fd_sc_hd__nor2_1 _393_ (.A(_063_),
    .B(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__a2111oi_2 _394_ (.A1(_063_),
    .A2(_136_),
    .B1(_140_),
    .C1(_142_),
    .D1(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__nor2_1 _395_ (.A(\mem[0][2] ),
    .B(_098_),
    .Y(_148_));
 sky130_fd_sc_hd__nand2_1 _396_ (.A(net15),
    .B(_060_),
    .Y(_149_));
 sky130_fd_sc_hd__o31ai_1 _397_ (.A1(_060_),
    .A2(_147_),
    .A3(_148_),
    .B1(_149_),
    .Y(_022_));
 sky130_fd_sc_hd__a22oi_1 _398_ (.A1(\mem[12][3] ),
    .A2(_079_),
    .B1(_067_),
    .B2(\mem[14][3] ),
    .Y(_150_));
 sky130_fd_sc_hd__a221oi_1 _399_ (.A1(\mem[6][3] ),
    .A2(_073_),
    .B1(_074_),
    .B2(\mem[5][3] ),
    .C1(_116_),
    .Y(_151_));
 sky130_fd_sc_hd__a211oi_1 _400_ (.A1(_104_),
    .A2(_150_),
    .B1(_151_),
    .C1(_103_),
    .Y(_152_));
 sky130_fd_sc_hd__nand3b_1 _401_ (.A_N(_116_),
    .B(\mem[4][3] ),
    .C(_079_),
    .Y(_153_));
 sky130_fd_sc_hd__a22oi_1 _402_ (.A1(\mem[8][3] ),
    .A2(_246_),
    .B1(_247_),
    .B2(\mem[10][3] ),
    .Y(_154_));
 sky130_fd_sc_hd__nand2_1 _403_ (.A(_066_),
    .B(\mem[11][3] ),
    .Y(_155_));
 sky130_fd_sc_hd__and3_1 _404_ (.A(_064_),
    .B(_154_),
    .C(_155_),
    .X(_156_));
 sky130_fd_sc_hd__or2_0 _405_ (.A(_061_),
    .B(_064_),
    .X(_157_));
 sky130_fd_sc_hd__a221oi_1 _406_ (.A1(_085_),
    .A2(\mem[3][3] ),
    .B1(\mem[1][3] ),
    .B2(_070_),
    .C1(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__a211oi_1 _407_ (.A1(_063_),
    .A2(_153_),
    .B1(_156_),
    .C1(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__nand2_1 _408_ (.A(_104_),
    .B(_070_),
    .Y(_160_));
 sky130_fd_sc_hd__mux2i_1 _409_ (.A0(\mem[9][3] ),
    .A1(\mem[13][3] ),
    .S(_062_),
    .Y(_161_));
 sky130_fd_sc_hd__o21ai_0 _410_ (.A1(_160_),
    .A2(_161_),
    .B1(_097_),
    .Y(_162_));
 sky130_fd_sc_hd__mux2i_1 _411_ (.A0(\mem[7][3] ),
    .A1(\mem[15][3] ),
    .S(_065_),
    .Y(_163_));
 sky130_fd_sc_hd__nand3_1 _412_ (.A(\mem[2][3] ),
    .B(_106_),
    .C(_127_),
    .Y(_164_));
 sky130_fd_sc_hd__o21ai_1 _413_ (.A1(_119_),
    .A2(_163_),
    .B1(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__nor4_1 _414_ (.A(_152_),
    .B(_159_),
    .C(_162_),
    .D(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__nor2_1 _415_ (.A(\mem[0][3] ),
    .B(_098_),
    .Y(_167_));
 sky130_fd_sc_hd__nand2_1 _416_ (.A(net16),
    .B(_060_),
    .Y(_168_));
 sky130_fd_sc_hd__o31ai_1 _417_ (.A1(_102_),
    .A2(_166_),
    .A3(_167_),
    .B1(_168_),
    .Y(_023_));
 sky130_fd_sc_hd__a22oi_2 _418_ (.A1(\mem[4][4] ),
    .A2(_133_),
    .B1(_073_),
    .B2(\mem[6][4] ),
    .Y(_169_));
 sky130_fd_sc_hd__a22oi_2 _419_ (.A1(\mem[12][4] ),
    .A2(_133_),
    .B1(_067_),
    .B2(\mem[14][4] ),
    .Y(_170_));
 sky130_fd_sc_hd__o22ai_2 _420_ (.A1(_110_),
    .A2(_169_),
    .B1(_170_),
    .B2(_117_),
    .Y(_171_));
 sky130_fd_sc_hd__a21o_1 _421_ (.A1(\mem[13][4] ),
    .A2(_128_),
    .B1(_171_),
    .X(_172_));
 sky130_fd_sc_hd__a222oi_1 _422_ (.A1(_085_),
    .A2(\mem[11][4] ),
    .B1(\mem[8][4] ),
    .B2(_079_),
    .C1(_070_),
    .C2(\mem[9][4] ),
    .Y(_173_));
 sky130_fd_sc_hd__mux2i_1 _423_ (.A0(\mem[7][4] ),
    .A1(\mem[15][4] ),
    .S(_084_),
    .Y(_174_));
 sky130_fd_sc_hd__o221ai_1 _424_ (.A1(_113_),
    .A2(_173_),
    .B1(_174_),
    .B2(_119_),
    .C1(_098_),
    .Y(_175_));
 sky130_fd_sc_hd__a22oi_1 _425_ (.A1(_085_),
    .A2(\mem[3][4] ),
    .B1(\mem[1][4] ),
    .B2(_070_),
    .Y(_176_));
 sky130_fd_sc_hd__nand3_1 _426_ (.A(_065_),
    .B(\mem[10][4] ),
    .C(_106_),
    .Y(_177_));
 sky130_fd_sc_hd__o21ai_0 _427_ (.A1(_104_),
    .A2(_176_),
    .B1(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__and3_1 _428_ (.A(_062_),
    .B(\mem[5][4] ),
    .C(_074_),
    .X(_179_));
 sky130_fd_sc_hd__a31oi_1 _429_ (.A1(_103_),
    .A2(\mem[2][4] ),
    .A3(_106_),
    .B1(_179_),
    .Y(_180_));
 sky130_fd_sc_hd__o2bb2ai_1 _430_ (.A1_N(_103_),
    .A2_N(_178_),
    .B1(_180_),
    .B2(_104_),
    .Y(_181_));
 sky130_fd_sc_hd__nor3_1 _431_ (.A(_172_),
    .B(_175_),
    .C(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__nor2_1 _432_ (.A(\mem[0][4] ),
    .B(_098_),
    .Y(_183_));
 sky130_fd_sc_hd__nand2_1 _433_ (.A(net17),
    .B(_060_),
    .Y(_184_));
 sky130_fd_sc_hd__o31ai_1 _434_ (.A1(_102_),
    .A2(_182_),
    .A3(_183_),
    .B1(_184_),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_1 _435_ (.A(_063_),
    .B(\mem[13][5] ),
    .Y(_185_));
 sky130_fd_sc_hd__nand3_1 _436_ (.A(_085_),
    .B(\mem[3][5] ),
    .C(_127_),
    .Y(_186_));
 sky130_fd_sc_hd__o21ai_0 _437_ (.A1(_160_),
    .A2(_185_),
    .B1(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__mux2i_2 _438_ (.A0(\mem[7][5] ),
    .A1(\mem[15][5] ),
    .S(_084_),
    .Y(_188_));
 sky130_fd_sc_hd__nand3_1 _439_ (.A(\mem[2][5] ),
    .B(_106_),
    .C(_127_),
    .Y(_189_));
 sky130_fd_sc_hd__o211ai_1 _440_ (.A1(_119_),
    .A2(_188_),
    .B1(_189_),
    .C1(_098_),
    .Y(_190_));
 sky130_fd_sc_hd__a22oi_1 _441_ (.A1(\mem[12][5] ),
    .A2(_246_),
    .B1(_073_),
    .B2(\mem[14][5] ),
    .Y(_191_));
 sky130_fd_sc_hd__a221oi_1 _442_ (.A1(\mem[6][5] ),
    .A2(_247_),
    .B1(_069_),
    .B2(\mem[5][5] ),
    .C1(_064_),
    .Y(_192_));
 sky130_fd_sc_hd__a21oi_1 _443_ (.A1(_116_),
    .A2(_191_),
    .B1(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__a22oi_1 _444_ (.A1(\mem[10][5] ),
    .A2(_073_),
    .B1(_074_),
    .B2(\mem[9][5] ),
    .Y(_194_));
 sky130_fd_sc_hd__a22oi_1 _445_ (.A1(_066_),
    .A2(\mem[11][5] ),
    .B1(\mem[8][5] ),
    .B2(_133_),
    .Y(_195_));
 sky130_fd_sc_hd__a21oi_1 _446_ (.A1(_194_),
    .A2(_195_),
    .B1(_113_),
    .Y(_196_));
 sky130_fd_sc_hd__nand3_1 _447_ (.A(_062_),
    .B(\mem[4][5] ),
    .C(_079_),
    .Y(_197_));
 sky130_fd_sc_hd__nand3b_1 _448_ (.A_N(_061_),
    .B(\mem[1][5] ),
    .C(_074_),
    .Y(_198_));
 sky130_fd_sc_hd__a21oi_1 _449_ (.A1(_197_),
    .A2(_198_),
    .B1(_065_),
    .Y(_199_));
 sky130_fd_sc_hd__a211o_1 _450_ (.A1(_063_),
    .A2(_193_),
    .B1(_196_),
    .C1(_199_),
    .X(_200_));
 sky130_fd_sc_hd__nor3_1 _451_ (.A(_187_),
    .B(_190_),
    .C(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__nor2_1 _452_ (.A(\mem[0][5] ),
    .B(_098_),
    .Y(_202_));
 sky130_fd_sc_hd__nand2_1 _453_ (.A(net18),
    .B(_060_),
    .Y(_203_));
 sky130_fd_sc_hd__o31ai_1 _454_ (.A1(_102_),
    .A2(_201_),
    .A3(_202_),
    .B1(_203_),
    .Y(_025_));
 sky130_fd_sc_hd__a22oi_2 _455_ (.A1(\mem[12][6] ),
    .A2(_133_),
    .B1(_067_),
    .B2(\mem[14][6] ),
    .Y(_204_));
 sky130_fd_sc_hd__a221oi_1 _456_ (.A1(\mem[6][6] ),
    .A2(_073_),
    .B1(_074_),
    .B2(\mem[5][6] ),
    .C1(_116_),
    .Y(_205_));
 sky130_fd_sc_hd__a211oi_2 _457_ (.A1(_104_),
    .A2(_204_),
    .B1(_205_),
    .C1(_103_),
    .Y(_206_));
 sky130_fd_sc_hd__nand3b_1 _458_ (.A_N(_116_),
    .B(\mem[4][6] ),
    .C(_079_),
    .Y(_207_));
 sky130_fd_sc_hd__a22oi_1 _459_ (.A1(\mem[8][6] ),
    .A2(_246_),
    .B1(_247_),
    .B2(\mem[10][6] ),
    .Y(_208_));
 sky130_fd_sc_hd__nand2_1 _460_ (.A(_066_),
    .B(\mem[11][6] ),
    .Y(_209_));
 sky130_fd_sc_hd__and3_1 _461_ (.A(_064_),
    .B(_208_),
    .C(_209_),
    .X(_210_));
 sky130_fd_sc_hd__a221oi_1 _462_ (.A1(_085_),
    .A2(\mem[3][6] ),
    .B1(\mem[1][6] ),
    .B2(_070_),
    .C1(_157_),
    .Y(_211_));
 sky130_fd_sc_hd__a211oi_1 _463_ (.A1(_063_),
    .A2(_207_),
    .B1(_210_),
    .C1(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__mux2i_1 _464_ (.A0(\mem[9][6] ),
    .A1(\mem[13][6] ),
    .S(_062_),
    .Y(_213_));
 sky130_fd_sc_hd__o21ai_0 _465_ (.A1(_160_),
    .A2(_213_),
    .B1(_097_),
    .Y(_214_));
 sky130_fd_sc_hd__mux2i_1 _466_ (.A0(\mem[7][6] ),
    .A1(\mem[15][6] ),
    .S(_065_),
    .Y(_215_));
 sky130_fd_sc_hd__nand3_1 _467_ (.A(\mem[2][6] ),
    .B(_106_),
    .C(_127_),
    .Y(_216_));
 sky130_fd_sc_hd__o21ai_1 _468_ (.A1(_119_),
    .A2(_215_),
    .B1(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__nor4_1 _469_ (.A(_206_),
    .B(_212_),
    .C(_214_),
    .D(_217_),
    .Y(_218_));
 sky130_fd_sc_hd__nor2_1 _470_ (.A(\mem[0][6] ),
    .B(_098_),
    .Y(_219_));
 sky130_fd_sc_hd__nand2_1 _471_ (.A(net19),
    .B(_060_),
    .Y(_220_));
 sky130_fd_sc_hd__o31ai_1 _472_ (.A1(_102_),
    .A2(_218_),
    .A3(_219_),
    .B1(_220_),
    .Y(_026_));
 sky130_fd_sc_hd__a22oi_1 _473_ (.A1(_066_),
    .A2(\mem[3][7] ),
    .B1(\mem[1][7] ),
    .B2(_074_),
    .Y(_221_));
 sky130_fd_sc_hd__nand3_1 _474_ (.A(_084_),
    .B(\mem[10][7] ),
    .C(_106_),
    .Y(_222_));
 sky130_fd_sc_hd__o21ai_0 _475_ (.A1(_065_),
    .A2(_221_),
    .B1(_222_),
    .Y(_223_));
 sky130_fd_sc_hd__mux2i_1 _476_ (.A0(\mem[7][7] ),
    .A1(\mem[15][7] ),
    .S(_041_),
    .Y(_224_));
 sky130_fd_sc_hd__nor2_1 _477_ (.A(_119_),
    .B(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__a211o_1 _478_ (.A1(\mem[13][7] ),
    .A2(_128_),
    .B1(_225_),
    .C1(_083_),
    .X(_226_));
 sky130_fd_sc_hd__and3_1 _479_ (.A(_061_),
    .B(\mem[5][7] ),
    .C(_069_),
    .X(_227_));
 sky130_fd_sc_hd__a31oi_1 _480_ (.A1(_103_),
    .A2(\mem[2][7] ),
    .A3(_067_),
    .B1(_227_),
    .Y(_228_));
 sky130_fd_sc_hd__a222oi_1 _481_ (.A1(_066_),
    .A2(\mem[11][7] ),
    .B1(\mem[8][7] ),
    .B2(_133_),
    .C1(_074_),
    .C2(\mem[9][7] ),
    .Y(_229_));
 sky130_fd_sc_hd__o22ai_1 _482_ (.A1(_104_),
    .A2(_228_),
    .B1(_229_),
    .B2(_113_),
    .Y(_230_));
 sky130_fd_sc_hd__a22oi_1 _483_ (.A1(\mem[12][7] ),
    .A2(_133_),
    .B1(_067_),
    .B2(\mem[14][7] ),
    .Y(_231_));
 sky130_fd_sc_hd__a221oi_1 _484_ (.A1(\mem[4][7] ),
    .A2(_133_),
    .B1(_067_),
    .B2(\mem[6][7] ),
    .C1(_116_),
    .Y(_232_));
 sky130_fd_sc_hd__a211oi_1 _485_ (.A1(_104_),
    .A2(_231_),
    .B1(_232_),
    .C1(_103_),
    .Y(_233_));
 sky130_fd_sc_hd__a2111oi_2 _486_ (.A1(_103_),
    .A2(_223_),
    .B1(_226_),
    .C1(_230_),
    .D1(_233_),
    .Y(_234_));
 sky130_fd_sc_hd__nor2_1 _487_ (.A(\mem[0][7] ),
    .B(_098_),
    .Y(_235_));
 sky130_fd_sc_hd__nand2_1 _488_ (.A(net20),
    .B(_060_),
    .Y(_236_));
 sky130_fd_sc_hd__o31ai_1 _489_ (.A1(_102_),
    .A2(_234_),
    .A3(_235_),
    .B1(_236_),
    .Y(_027_));
 sky130_fd_sc_hd__xnor2_1 _490_ (.A(\rd_ptr[0] ),
    .B(_060_),
    .Y(_028_));
 sky130_fd_sc_hd__mux2_1 _491_ (.A0(_019_),
    .A1(\rd_ptr[1] ),
    .S(_102_),
    .X(_029_));
 sky130_fd_sc_hd__inv_1 _492_ (.A(_085_),
    .Y(_237_));
 sky130_fd_sc_hd__nor2_1 _493_ (.A(_237_),
    .B(_102_),
    .Y(_238_));
 sky130_fd_sc_hd__xnor2_1 _494_ (.A(_103_),
    .B(_238_),
    .Y(_030_));
 sky130_fd_sc_hd__nor4_1 _495_ (.A(_018_),
    .B(_245_),
    .C(_103_),
    .D(_102_),
    .Y(_239_));
 sky130_fd_sc_hd__xor2_1 _496_ (.A(_104_),
    .B(_239_),
    .X(_031_));
 sky130_fd_sc_hd__or3_1 _497_ (.A(_237_),
    .B(_059_),
    .C(_117_),
    .X(_240_));
 sky130_fd_sc_hd__xnor2_1 _498_ (.A(\rd_ptr[4] ),
    .B(_240_),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_1 _499_ (.A(_016_),
    .B(_049_),
    .Y(_033_));
 sky130_fd_sc_hd__nand2_1 _500_ (.A(_017_),
    .B(_049_),
    .Y(_241_));
 sky130_fd_sc_hd__o21ai_0 _501_ (.A1(_253_),
    .A2(_049_),
    .B1(_241_),
    .Y(_034_));
 sky130_fd_sc_hd__nand2_1 _502_ (.A(_259_),
    .B(_049_),
    .Y(_242_));
 sky130_fd_sc_hd__xnor2_1 _503_ (.A(_044_),
    .B(_242_),
    .Y(_035_));
 sky130_fd_sc_hd__nand4_1 _504_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .C(_044_),
    .D(_049_),
    .Y(_243_));
 sky130_fd_sc_hd__xnor2_1 _505_ (.A(_042_),
    .B(_243_),
    .Y(_036_));
 sky130_fd_sc_hd__nand4_1 _506_ (.A(_044_),
    .B(_042_),
    .C(_259_),
    .D(_049_),
    .Y(_244_));
 sky130_fd_sc_hd__xnor2_1 _507_ (.A(\wr_ptr[4] ),
    .B(_244_),
    .Y(_037_));
 sky130_fd_sc_hd__ha_2 _508_ (.A(_018_),
    .B(_245_),
    .COUT(_246_),
    .SUM(_019_));
 sky130_fd_sc_hd__ha_2 _509_ (.A(_018_),
    .B(\rd_ptr[1] ),
    .COUT(_247_),
    .SUM(_248_));
 sky130_fd_sc_hd__ha_1 _510_ (.A(\rd_ptr[0] ),
    .B(_245_),
    .COUT(_249_),
    .SUM(_250_));
 sky130_fd_sc_hd__ha_1 _511_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .COUT(_251_),
    .SUM(_252_));
 sky130_fd_sc_hd__ha_1 _512_ (.A(_016_),
    .B(_253_),
    .COUT(_254_),
    .SUM(_017_));
 sky130_fd_sc_hd__ha_1 _513_ (.A(_016_),
    .B(\wr_ptr[1] ),
    .COUT(_255_),
    .SUM(_256_));
 sky130_fd_sc_hd__ha_1 _514_ (.A(\wr_ptr[0] ),
    .B(_253_),
    .COUT(_257_),
    .SUM(_258_));
 sky130_fd_sc_hd__ha_2 _515_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .COUT(_259_),
    .SUM(_260_));
 sky130_fd_sc_hd__dfrtp_1 \dout[0]$_DFFE_PN0P_  (.D(_020_),
    .Q(net13),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dout[1]$_DFFE_PN0P_  (.D(_021_),
    .Q(net14),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dout[2]$_DFFE_PN0P_  (.D(_022_),
    .Q(net15),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dout[3]$_DFFE_PN0P_  (.D(_023_),
    .Q(net16),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dout[4]$_DFFE_PN0P_  (.D(_024_),
    .Q(net17),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dout[5]$_DFFE_PN0P_  (.D(_025_),
    .Q(net18),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dout[6]$_DFFE_PN0P_  (.D(_026_),
    .Q(net19),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \dout[7]$_DFFE_PN0P_  (.D(_027_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net2),
    .DE(_015_),
    .Q(\mem[0][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net3),
    .DE(_015_),
    .Q(\mem[0][1] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net4),
    .DE(_015_),
    .Q(\mem[0][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\mem[0][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\mem[0][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\mem[0][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\mem[0][6] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\mem[0][7] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net2),
    .DE(_005_),
    .Q(\mem[10][0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net3),
    .DE(_005_),
    .Q(\mem[10][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net4),
    .DE(_005_),
    .Q(\mem[10][2] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net5),
    .DE(_005_),
    .Q(\mem[10][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net6),
    .DE(_005_),
    .Q(\mem[10][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net7),
    .DE(_005_),
    .Q(\mem[10][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net8),
    .DE(_005_),
    .Q(\mem[10][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net9),
    .DE(_005_),
    .Q(\mem[10][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net2),
    .DE(_004_),
    .Q(\mem[11][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net3),
    .DE(_004_),
    .Q(\mem[11][1] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net4),
    .DE(_004_),
    .Q(\mem[11][2] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net5),
    .DE(_004_),
    .Q(\mem[11][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net6),
    .DE(_004_),
    .Q(\mem[11][4] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net7),
    .DE(_004_),
    .Q(\mem[11][5] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net8),
    .DE(_004_),
    .Q(\mem[11][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net9),
    .DE(_004_),
    .Q(\mem[11][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net2),
    .DE(_003_),
    .Q(\mem[12][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net3),
    .DE(_003_),
    .Q(\mem[12][1] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net4),
    .DE(_003_),
    .Q(\mem[12][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net5),
    .DE(_003_),
    .Q(\mem[12][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net6),
    .DE(_003_),
    .Q(\mem[12][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net7),
    .DE(_003_),
    .Q(\mem[12][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net8),
    .DE(_003_),
    .Q(\mem[12][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net9),
    .DE(_003_),
    .Q(\mem[12][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net2),
    .DE(_002_),
    .Q(\mem[13][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net3),
    .DE(_002_),
    .Q(\mem[13][1] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net4),
    .DE(_002_),
    .Q(\mem[13][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net5),
    .DE(_002_),
    .Q(\mem[13][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net6),
    .DE(_002_),
    .Q(\mem[13][4] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net7),
    .DE(_002_),
    .Q(\mem[13][5] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net8),
    .DE(_002_),
    .Q(\mem[13][6] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net9),
    .DE(_002_),
    .Q(\mem[13][7] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net2),
    .DE(_001_),
    .Q(\mem[14][0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net3),
    .DE(_001_),
    .Q(\mem[14][1] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net4),
    .DE(_001_),
    .Q(\mem[14][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net5),
    .DE(_001_),
    .Q(\mem[14][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net6),
    .DE(_001_),
    .Q(\mem[14][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net7),
    .DE(_001_),
    .Q(\mem[14][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net8),
    .DE(_001_),
    .Q(\mem[14][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net9),
    .DE(_001_),
    .Q(\mem[14][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net2),
    .DE(_000_),
    .Q(\mem[15][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net3),
    .DE(_000_),
    .Q(\mem[15][1] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net4),
    .DE(_000_),
    .Q(\mem[15][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net5),
    .DE(_000_),
    .Q(\mem[15][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net6),
    .DE(_000_),
    .Q(\mem[15][4] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net7),
    .DE(_000_),
    .Q(\mem[15][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net8),
    .DE(_000_),
    .Q(\mem[15][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net9),
    .DE(_000_),
    .Q(\mem[15][7] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net2),
    .DE(_014_),
    .Q(\mem[1][0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net3),
    .DE(_014_),
    .Q(\mem[1][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net4),
    .DE(_014_),
    .Q(\mem[1][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\mem[1][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\mem[1][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\mem[1][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\mem[1][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\mem[1][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net2),
    .DE(_013_),
    .Q(\mem[2][0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net3),
    .DE(_013_),
    .Q(\mem[2][1] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net4),
    .DE(_013_),
    .Q(\mem[2][2] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\mem[2][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\mem[2][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\mem[2][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\mem[2][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\mem[2][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net2),
    .DE(_012_),
    .Q(\mem[3][0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net3),
    .DE(_012_),
    .Q(\mem[3][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net4),
    .DE(_012_),
    .Q(\mem[3][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\mem[3][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\mem[3][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\mem[3][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\mem[3][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\mem[3][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net2),
    .DE(_011_),
    .Q(\mem[4][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net3),
    .DE(_011_),
    .Q(\mem[4][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net4),
    .DE(_011_),
    .Q(\mem[4][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\mem[4][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\mem[4][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\mem[4][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\mem[4][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\mem[4][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net2),
    .DE(_010_),
    .Q(\mem[5][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net3),
    .DE(_010_),
    .Q(\mem[5][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net4),
    .DE(_010_),
    .Q(\mem[5][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net5),
    .DE(_010_),
    .Q(\mem[5][3] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net6),
    .DE(_010_),
    .Q(\mem[5][4] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net7),
    .DE(_010_),
    .Q(\mem[5][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net8),
    .DE(_010_),
    .Q(\mem[5][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net9),
    .DE(_010_),
    .Q(\mem[5][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net2),
    .DE(_009_),
    .Q(\mem[6][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net3),
    .DE(_009_),
    .Q(\mem[6][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net4),
    .DE(_009_),
    .Q(\mem[6][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net5),
    .DE(_009_),
    .Q(\mem[6][3] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net6),
    .DE(_009_),
    .Q(\mem[6][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net7),
    .DE(_009_),
    .Q(\mem[6][5] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net8),
    .DE(_009_),
    .Q(\mem[6][6] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net9),
    .DE(_009_),
    .Q(\mem[6][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net2),
    .DE(_008_),
    .Q(\mem[7][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net3),
    .DE(_008_),
    .Q(\mem[7][1] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net4),
    .DE(_008_),
    .Q(\mem[7][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net5),
    .DE(_008_),
    .Q(\mem[7][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net6),
    .DE(_008_),
    .Q(\mem[7][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net7),
    .DE(_008_),
    .Q(\mem[7][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net8),
    .DE(_008_),
    .Q(\mem[7][6] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net9),
    .DE(_008_),
    .Q(\mem[7][7] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net2),
    .DE(_007_),
    .Q(\mem[8][0] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net3),
    .DE(_007_),
    .Q(\mem[8][1] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net4),
    .DE(_007_),
    .Q(\mem[8][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net5),
    .DE(_007_),
    .Q(\mem[8][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net6),
    .DE(_007_),
    .Q(\mem[8][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net7),
    .DE(_007_),
    .Q(\mem[8][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net8),
    .DE(_007_),
    .Q(\mem[8][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net9),
    .DE(_007_),
    .Q(\mem[8][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net2),
    .DE(_006_),
    .Q(\mem[9][0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net3),
    .DE(_006_),
    .Q(\mem[9][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net4),
    .DE(_006_),
    .Q(\mem[9][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net5),
    .DE(_006_),
    .Q(\mem[9][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net6),
    .DE(_006_),
    .Q(\mem[9][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net7),
    .DE(_006_),
    .Q(\mem[9][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net8),
    .DE(_006_),
    .Q(\mem[9][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net9),
    .DE(_006_),
    .Q(\mem[9][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr[0]$_DFFE_PN0P_  (.D(_028_),
    .Q(\rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[1]$_DFFE_PN0P_  (.D(_029_),
    .Q(\rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[2]$_DFFE_PN0P_  (.D(_030_),
    .Q(\rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[3]$_DFFE_PN0P_  (.D(_031_),
    .Q(\rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[4]$_DFFE_PN0P_  (.D(_032_),
    .Q(\rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[0]$_DFFE_PN0P_  (.D(_033_),
    .Q(\wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[1]$_DFFE_PN0P_  (.D(_034_),
    .Q(\wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[2]$_DFFE_PN0P_  (.D(_035_),
    .Q(\wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[3]$_DFFE_PN0P_  (.D(_036_),
    .Q(\wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[4]$_DFFE_PN0P_  (.D(_037_),
    .Q(\wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__buf_6 hold1 (.A(net11),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_135 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(net24),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input2 (.A(din[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input3 (.A(din[2]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input4 (.A(din[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input5 (.A(din[4]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input6 (.A(din[5]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input7 (.A(din[6]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input8 (.A(din[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(rd_en),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input10 (.A(net23),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(wr_en),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(dout[0]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(dout[1]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(dout[2]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(dout[3]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(dout[4]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(dout[5]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(dout[6]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(dout[7]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(full));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload5 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload6 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload7 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload8 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload9 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(din[0]),
    .X(net24));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_223 ();
endmodule
