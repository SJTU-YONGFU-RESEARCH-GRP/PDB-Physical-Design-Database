module parameterized_self_correcting_counter (clk,
    enable,
    rst_n,
    count);
 input clk;
 input enable;
 input rst_n;
 output [3:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _30_ (.A(net1),
    .ZN(_04_));
 BUF_X2 _31_ (.A(net2),
    .Z(_05_));
 INV_X1 _32_ (.A(_05_),
    .ZN(_06_));
 BUF_X4 _33_ (.A(enable),
    .Z(_07_));
 BUF_X1 _34_ (.A(net5),
    .Z(_08_));
 BUF_X4 _35_ (.A(net3),
    .Z(_09_));
 OAI21_X1 _36_ (.A(_08_),
    .B1(net4),
    .B2(_09_),
    .ZN(_10_));
 NAND3_X1 _37_ (.A1(_06_),
    .A2(_07_),
    .A3(_10_),
    .ZN(_11_));
 INV_X4 _38_ (.A(_07_),
    .ZN(_12_));
 NAND2_X1 _39_ (.A1(_05_),
    .A2(_12_),
    .ZN(_13_));
 AOI21_X1 _40_ (.A(_04_),
    .B1(_11_),
    .B2(_13_),
    .ZN(_00_));
 OAI21_X1 _41_ (.A(_07_),
    .B1(_08_),
    .B2(_05_),
    .ZN(_14_));
 NAND2_X1 _42_ (.A1(_09_),
    .A2(_14_),
    .ZN(_15_));
 OR4_X1 _43_ (.A1(_06_),
    .A2(_09_),
    .A3(_08_),
    .A4(_12_),
    .ZN(_16_));
 AOI21_X1 _44_ (.A(_04_),
    .B1(_15_),
    .B2(_16_),
    .ZN(_01_));
 AND2_X1 _45_ (.A1(_05_),
    .A2(_09_),
    .ZN(_17_));
 OR2_X1 _46_ (.A1(_08_),
    .A2(_17_),
    .ZN(_18_));
 AND2_X1 _47_ (.A1(net4),
    .A2(_07_),
    .ZN(_19_));
 INV_X1 _48_ (.A(_08_),
    .ZN(_20_));
 NAND3_X1 _49_ (.A1(_20_),
    .A2(_07_),
    .A3(_17_),
    .ZN(_21_));
 INV_X1 _50_ (.A(net4),
    .ZN(_22_));
 AOI221_X1 _51_ (.A(_04_),
    .B1(_18_),
    .B2(_19_),
    .C1(_21_),
    .C2(_22_),
    .ZN(_02_));
 NAND3_X1 _52_ (.A1(_20_),
    .A2(_17_),
    .A3(_19_),
    .ZN(_23_));
 NOR3_X1 _53_ (.A1(_05_),
    .A2(_09_),
    .A3(net4),
    .ZN(_24_));
 OAI21_X1 _54_ (.A(_08_),
    .B1(_12_),
    .B2(_24_),
    .ZN(_25_));
 AOI21_X1 _55_ (.A(_04_),
    .B1(_23_),
    .B2(_25_),
    .ZN(_03_));
 DFF_X1 \counter_reg[0]$_SDFFE_PN0P_  (.D(_00_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net2),
    .QN(_29_));
 DFF_X1 \counter_reg[1]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net3),
    .QN(_28_));
 DFF_X1 \counter_reg[2]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net4),
    .QN(_27_));
 DFF_X1 \counter_reg[3]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net5),
    .QN(_26_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_43 ();
 BUF_X1 input1 (.A(rst_n),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(count[0]));
 BUF_X1 output3 (.A(net3),
    .Z(count[1]));
 BUF_X1 output4 (.A(net4),
    .Z(count[2]));
 BUF_X1 output5 (.A(net5),
    .Z(count[3]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_81 ();
 FILLCELL_X1 FILLER_0_85 ();
 FILLCELL_X8 FILLER_0_92 ();
 FILLCELL_X1 FILLER_0_100 ();
 FILLCELL_X32 FILLER_0_104 ();
 FILLCELL_X32 FILLER_0_136 ();
 FILLCELL_X1 FILLER_0_168 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X16 FILLER_1_65 ();
 FILLCELL_X2 FILLER_1_81 ();
 FILLCELL_X1 FILLER_1_83 ();
 FILLCELL_X1 FILLER_1_106 ();
 FILLCELL_X32 FILLER_1_109 ();
 FILLCELL_X16 FILLER_1_141 ();
 FILLCELL_X8 FILLER_1_157 ();
 FILLCELL_X4 FILLER_1_165 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X16 FILLER_2_65 ();
 FILLCELL_X8 FILLER_2_81 ();
 FILLCELL_X8 FILLER_2_92 ();
 FILLCELL_X2 FILLER_2_100 ();
 FILLCELL_X1 FILLER_2_102 ();
 FILLCELL_X32 FILLER_2_111 ();
 FILLCELL_X16 FILLER_2_143 ();
 FILLCELL_X8 FILLER_2_159 ();
 FILLCELL_X2 FILLER_2_167 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X4 FILLER_3_65 ();
 FILLCELL_X2 FILLER_3_69 ();
 FILLCELL_X1 FILLER_3_71 ();
 FILLCELL_X8 FILLER_3_89 ();
 FILLCELL_X2 FILLER_3_97 ();
 FILLCELL_X1 FILLER_3_99 ();
 FILLCELL_X1 FILLER_3_102 ();
 FILLCELL_X32 FILLER_3_111 ();
 FILLCELL_X16 FILLER_3_143 ();
 FILLCELL_X8 FILLER_3_159 ();
 FILLCELL_X2 FILLER_3_167 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X1 FILLER_4_105 ();
 FILLCELL_X32 FILLER_4_110 ();
 FILLCELL_X16 FILLER_4_142 ();
 FILLCELL_X8 FILLER_4_158 ();
 FILLCELL_X2 FILLER_4_166 ();
 FILLCELL_X1 FILLER_4_168 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X16 FILLER_5_65 ();
 FILLCELL_X8 FILLER_5_81 ();
 FILLCELL_X2 FILLER_5_89 ();
 FILLCELL_X1 FILLER_5_91 ();
 FILLCELL_X1 FILLER_5_100 ();
 FILLCELL_X32 FILLER_5_105 ();
 FILLCELL_X32 FILLER_5_137 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X16 FILLER_6_65 ();
 FILLCELL_X8 FILLER_6_81 ();
 FILLCELL_X1 FILLER_6_98 ();
 FILLCELL_X2 FILLER_6_103 ();
 FILLCELL_X1 FILLER_6_105 ();
 FILLCELL_X32 FILLER_6_111 ();
 FILLCELL_X16 FILLER_6_143 ();
 FILLCELL_X8 FILLER_6_159 ();
 FILLCELL_X2 FILLER_6_167 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_65 ();
 FILLCELL_X8 FILLER_7_81 ();
 FILLCELL_X4 FILLER_7_89 ();
 FILLCELL_X4 FILLER_7_107 ();
 FILLCELL_X2 FILLER_7_111 ();
 FILLCELL_X1 FILLER_7_113 ();
 FILLCELL_X32 FILLER_7_121 ();
 FILLCELL_X16 FILLER_7_153 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X8 FILLER_8_65 ();
 FILLCELL_X4 FILLER_8_73 ();
 FILLCELL_X1 FILLER_8_77 ();
 FILLCELL_X1 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_108 ();
 FILLCELL_X16 FILLER_8_140 ();
 FILLCELL_X8 FILLER_8_156 ();
 FILLCELL_X4 FILLER_8_164 ();
 FILLCELL_X1 FILLER_8_168 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X4 FILLER_9_81 ();
 FILLCELL_X1 FILLER_9_85 ();
 FILLCELL_X32 FILLER_9_90 ();
 FILLCELL_X32 FILLER_9_122 ();
 FILLCELL_X8 FILLER_9_154 ();
 FILLCELL_X4 FILLER_9_162 ();
 FILLCELL_X2 FILLER_9_166 ();
 FILLCELL_X1 FILLER_9_168 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X16 FILLER_10_65 ();
 FILLCELL_X4 FILLER_10_81 ();
 FILLCELL_X32 FILLER_10_102 ();
 FILLCELL_X32 FILLER_10_134 ();
 FILLCELL_X2 FILLER_10_166 ();
 FILLCELL_X1 FILLER_10_168 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X16 FILLER_11_65 ();
 FILLCELL_X8 FILLER_11_81 ();
 FILLCELL_X1 FILLER_11_89 ();
 FILLCELL_X2 FILLER_11_95 ();
 FILLCELL_X32 FILLER_11_104 ();
 FILLCELL_X32 FILLER_11_136 ();
 FILLCELL_X1 FILLER_11_168 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X8 FILLER_12_161 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X8 FILLER_13_161 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X8 FILLER_14_161 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X8 FILLER_15_161 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_161 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X8 FILLER_17_161 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X8 FILLER_18_161 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X8 FILLER_19_161 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X8 FILLER_20_161 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X16 FILLER_21_65 ();
 FILLCELL_X2 FILLER_21_81 ();
 FILLCELL_X8 FILLER_21_86 ();
 FILLCELL_X1 FILLER_21_94 ();
 FILLCELL_X32 FILLER_21_98 ();
 FILLCELL_X32 FILLER_21_130 ();
 FILLCELL_X4 FILLER_21_162 ();
 FILLCELL_X2 FILLER_21_166 ();
 FILLCELL_X1 FILLER_21_168 ();
endmodule
