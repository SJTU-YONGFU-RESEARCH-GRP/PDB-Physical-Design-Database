module crossbar_switch (clk,
    rst_n,
    data_in,
    data_out,
    select);
 input clk;
 input rst_n;
 input [31:0] data_in;
 output [31:0] data_out;
 input [7:0] select;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 NAND2_X4 _213_ (.A1(net34),
    .A2(_163_),
    .ZN(_174_));
 MUX2_X1 _214_ (.A(net2),
    .B(net19),
    .S(_168_),
    .Z(_175_));
 INV_X1 _215_ (.A(_175_),
    .ZN(_176_));
 OAI22_X1 _216_ (.A1(_171_),
    .A2(_173_),
    .B1(_174_),
    .B2(_176_),
    .ZN(_001_));
 MUX2_X1 _217_ (.A(net26),
    .B(net11),
    .S(_169_),
    .Z(_177_));
 INV_X1 _218_ (.A(_177_),
    .ZN(_178_));
 MUX2_X1 _219_ (.A(net3),
    .B(net20),
    .S(_169_),
    .Z(_179_));
 INV_X1 _220_ (.A(_179_),
    .ZN(_180_));
 OAI22_X1 _221_ (.A1(_173_),
    .A2(_178_),
    .B1(_180_),
    .B2(_174_),
    .ZN(_002_));
 MUX2_X1 _222_ (.A(net27),
    .B(net13),
    .S(_169_),
    .Z(_032_));
 INV_X1 _223_ (.A(_032_),
    .ZN(_033_));
 MUX2_X1 _224_ (.A(net4),
    .B(net21),
    .S(_169_),
    .Z(_034_));
 INV_X1 _225_ (.A(_034_),
    .ZN(_035_));
 OAI22_X1 _226_ (.A1(_173_),
    .A2(_033_),
    .B1(_035_),
    .B2(_174_),
    .ZN(_003_));
 MUX2_X1 _227_ (.A(net28),
    .B(net14),
    .S(_169_),
    .Z(_036_));
 INV_X1 _228_ (.A(_036_),
    .ZN(_037_));
 MUX2_X1 _229_ (.A(net5),
    .B(net22),
    .S(_168_),
    .Z(_038_));
 INV_X1 _230_ (.A(_038_),
    .ZN(_039_));
 OAI22_X1 _231_ (.A1(_173_),
    .A2(_037_),
    .B1(_039_),
    .B2(_174_),
    .ZN(_004_));
 MUX2_X1 _232_ (.A(net29),
    .B(net15),
    .S(_169_),
    .Z(_040_));
 INV_X1 _233_ (.A(_040_),
    .ZN(_041_));
 MUX2_X1 _234_ (.A(net6),
    .B(net24),
    .S(_168_),
    .Z(_042_));
 INV_X1 _235_ (.A(_042_),
    .ZN(_043_));
 OAI22_X1 _236_ (.A1(_173_),
    .A2(_041_),
    .B1(_043_),
    .B2(_174_),
    .ZN(_005_));
 MUX2_X1 _237_ (.A(net30),
    .B(net16),
    .S(_169_),
    .Z(_044_));
 INV_X1 _238_ (.A(_044_),
    .ZN(_045_));
 MUX2_X1 _239_ (.A(net7),
    .B(net25),
    .S(_168_),
    .Z(_046_));
 INV_X1 _240_ (.A(_046_),
    .ZN(_047_));
 OAI22_X1 _241_ (.A1(_173_),
    .A2(_045_),
    .B1(_047_),
    .B2(_174_),
    .ZN(_006_));
 BUF_X8 _242_ (.A(select[5]),
    .Z(_048_));
 BUF_X8 _243_ (.A(_048_),
    .Z(_049_));
 MUX2_X1 _244_ (.A(net1),
    .B(net8),
    .S(_049_),
    .Z(_050_));
 INV_X1 _245_ (.A(_050_),
    .ZN(_051_));
 INV_X1 _246_ (.A(net35),
    .ZN(_052_));
 NAND2_X4 _247_ (.A1(_052_),
    .A2(_163_),
    .ZN(_053_));
 NAND2_X4 _248_ (.A1(net35),
    .A2(_163_),
    .ZN(_054_));
 MUX2_X1 _249_ (.A(net31),
    .B(net17),
    .S(_048_),
    .Z(_055_));
 INV_X1 _250_ (.A(_055_),
    .ZN(_056_));
 OAI22_X1 _251_ (.A1(_051_),
    .A2(_053_),
    .B1(_054_),
    .B2(_056_),
    .ZN(_007_));
 MUX2_X1 _252_ (.A(net12),
    .B(net9),
    .S(_049_),
    .Z(_057_));
 INV_X1 _253_ (.A(_057_),
    .ZN(_058_));
 MUX2_X1 _254_ (.A(net32),
    .B(net18),
    .S(_049_),
    .Z(_059_));
 INV_X1 _255_ (.A(_059_),
    .ZN(_060_));
 OAI22_X1 _256_ (.A1(_053_),
    .A2(_058_),
    .B1(_060_),
    .B2(_054_),
    .ZN(_008_));
 MUX2_X1 _257_ (.A(net23),
    .B(net10),
    .S(_049_),
    .Z(_061_));
 INV_X1 _258_ (.A(_061_),
    .ZN(_062_));
 MUX2_X1 _259_ (.A(net2),
    .B(net19),
    .S(_049_),
    .Z(_063_));
 INV_X1 _260_ (.A(_063_),
    .ZN(_064_));
 OAI22_X1 _261_ (.A1(_053_),
    .A2(_062_),
    .B1(_064_),
    .B2(_054_),
    .ZN(_009_));
 MUX2_X1 _262_ (.A(net26),
    .B(net11),
    .S(_049_),
    .Z(_065_));
 INV_X1 _263_ (.A(_065_),
    .ZN(_066_));
 MUX2_X1 _264_ (.A(net3),
    .B(net20),
    .S(_048_),
    .Z(_067_));
 INV_X1 _265_ (.A(_067_),
    .ZN(_068_));
 OAI22_X1 _266_ (.A1(_053_),
    .A2(_066_),
    .B1(_068_),
    .B2(_054_),
    .ZN(_010_));
 MUX2_X1 _267_ (.A(net12),
    .B(net9),
    .S(_159_),
    .Z(_069_));
 INV_X1 _268_ (.A(_069_),
    .ZN(_070_));
 MUX2_X1 _269_ (.A(net32),
    .B(net18),
    .S(_159_),
    .Z(_071_));
 INV_X1 _270_ (.A(_071_),
    .ZN(_072_));
 OAI22_X1 _271_ (.A1(_164_),
    .A2(_070_),
    .B1(_072_),
    .B2(_165_),
    .ZN(_011_));
 MUX2_X1 _272_ (.A(net27),
    .B(net13),
    .S(_049_),
    .Z(_073_));
 INV_X1 _273_ (.A(_073_),
    .ZN(_074_));
 MUX2_X1 _274_ (.A(net4),
    .B(net21),
    .S(_048_),
    .Z(_075_));
 INV_X1 _275_ (.A(_075_),
    .ZN(_076_));
 OAI22_X1 _276_ (.A1(_053_),
    .A2(_074_),
    .B1(_076_),
    .B2(_054_),
    .ZN(_012_));
 MUX2_X1 _277_ (.A(net28),
    .B(net14),
    .S(_049_),
    .Z(_077_));
 INV_X1 _278_ (.A(_077_),
    .ZN(_078_));
 MUX2_X1 _279_ (.A(net5),
    .B(net22),
    .S(_048_),
    .Z(_079_));
 INV_X1 _280_ (.A(_079_),
    .ZN(_080_));
 OAI22_X1 _281_ (.A1(_053_),
    .A2(_078_),
    .B1(_080_),
    .B2(_054_),
    .ZN(_013_));
 MUX2_X1 _282_ (.A(net29),
    .B(net15),
    .S(_049_),
    .Z(_081_));
 INV_X1 _283_ (.A(_081_),
    .ZN(_082_));
 MUX2_X1 _284_ (.A(net6),
    .B(net24),
    .S(_048_),
    .Z(_083_));
 INV_X1 _285_ (.A(_083_),
    .ZN(_084_));
 OAI22_X1 _286_ (.A1(_053_),
    .A2(_082_),
    .B1(_084_),
    .B2(_054_),
    .ZN(_014_));
 MUX2_X1 _287_ (.A(net30),
    .B(net16),
    .S(_049_),
    .Z(_085_));
 INV_X1 _288_ (.A(_085_),
    .ZN(_086_));
 MUX2_X1 _289_ (.A(net7),
    .B(net25),
    .S(_048_),
    .Z(_087_));
 INV_X1 _290_ (.A(_087_),
    .ZN(_088_));
 OAI22_X1 _291_ (.A1(_053_),
    .A2(_086_),
    .B1(_088_),
    .B2(_054_),
    .ZN(_015_));
 BUF_X8 _292_ (.A(select[7]),
    .Z(_089_));
 BUF_X8 _293_ (.A(_089_),
    .Z(_090_));
 MUX2_X1 _294_ (.A(net1),
    .B(net8),
    .S(_090_),
    .Z(_091_));
 INV_X1 _295_ (.A(_091_),
    .ZN(_092_));
 INV_X1 _296_ (.A(net36),
    .ZN(_093_));
 NAND2_X4 _297_ (.A1(_093_),
    .A2(_163_),
    .ZN(_094_));
 NAND2_X4 _298_ (.A1(net36),
    .A2(_163_),
    .ZN(_095_));
 MUX2_X1 _299_ (.A(net31),
    .B(net17),
    .S(_089_),
    .Z(_096_));
 INV_X1 _300_ (.A(_096_),
    .ZN(_097_));
 OAI22_X1 _301_ (.A1(_092_),
    .A2(_094_),
    .B1(_095_),
    .B2(_097_),
    .ZN(_016_));
 MUX2_X1 _302_ (.A(net12),
    .B(net9),
    .S(_090_),
    .Z(_098_));
 INV_X1 _303_ (.A(_098_),
    .ZN(_099_));
 MUX2_X1 _304_ (.A(net32),
    .B(net18),
    .S(_090_),
    .Z(_100_));
 INV_X1 _305_ (.A(_100_),
    .ZN(_101_));
 OAI22_X1 _306_ (.A1(_094_),
    .A2(_099_),
    .B1(_101_),
    .B2(_095_),
    .ZN(_017_));
 MUX2_X1 _307_ (.A(net23),
    .B(net10),
    .S(_090_),
    .Z(_102_));
 INV_X1 _308_ (.A(_102_),
    .ZN(_103_));
 MUX2_X1 _309_ (.A(net2),
    .B(net19),
    .S(_090_),
    .Z(_104_));
 INV_X1 _310_ (.A(_104_),
    .ZN(_105_));
 OAI22_X1 _311_ (.A1(_094_),
    .A2(_103_),
    .B1(_105_),
    .B2(_095_),
    .ZN(_018_));
 MUX2_X1 _312_ (.A(net26),
    .B(net11),
    .S(_090_),
    .Z(_106_));
 INV_X1 _313_ (.A(_106_),
    .ZN(_107_));
 MUX2_X1 _314_ (.A(net3),
    .B(net20),
    .S(_089_),
    .Z(_108_));
 INV_X1 _315_ (.A(_108_),
    .ZN(_109_));
 OAI22_X1 _316_ (.A1(_094_),
    .A2(_107_),
    .B1(_109_),
    .B2(_095_),
    .ZN(_019_));
 MUX2_X1 _317_ (.A(net27),
    .B(net13),
    .S(_090_),
    .Z(_110_));
 INV_X1 _318_ (.A(_110_),
    .ZN(_111_));
 MUX2_X1 _319_ (.A(net4),
    .B(net21),
    .S(_089_),
    .Z(_112_));
 INV_X1 _320_ (.A(_112_),
    .ZN(_113_));
 OAI22_X1 _321_ (.A1(_094_),
    .A2(_111_),
    .B1(_113_),
    .B2(_095_),
    .ZN(_020_));
 MUX2_X1 _322_ (.A(net28),
    .B(net14),
    .S(_090_),
    .Z(_114_));
 INV_X1 _323_ (.A(_114_),
    .ZN(_115_));
 MUX2_X1 _324_ (.A(net5),
    .B(net22),
    .S(_089_),
    .Z(_116_));
 INV_X1 _325_ (.A(_116_),
    .ZN(_117_));
 OAI22_X1 _326_ (.A1(_094_),
    .A2(_115_),
    .B1(_117_),
    .B2(_095_),
    .ZN(_021_));
 MUX2_X1 _327_ (.A(net23),
    .B(net10),
    .S(_159_),
    .Z(_118_));
 INV_X1 _328_ (.A(_118_),
    .ZN(_119_));
 MUX2_X1 _329_ (.A(net2),
    .B(net19),
    .S(_159_),
    .Z(_120_));
 INV_X1 _330_ (.A(_120_),
    .ZN(_121_));
 OAI22_X1 _331_ (.A1(_164_),
    .A2(_119_),
    .B1(_121_),
    .B2(_165_),
    .ZN(_022_));
 MUX2_X1 _332_ (.A(net29),
    .B(net15),
    .S(_090_),
    .Z(_122_));
 INV_X1 _333_ (.A(_122_),
    .ZN(_123_));
 MUX2_X1 _334_ (.A(net6),
    .B(net24),
    .S(_089_),
    .Z(_124_));
 INV_X1 _335_ (.A(_124_),
    .ZN(_125_));
 OAI22_X1 _336_ (.A1(_094_),
    .A2(_123_),
    .B1(_125_),
    .B2(_095_),
    .ZN(_023_));
 MUX2_X1 _337_ (.A(net30),
    .B(net16),
    .S(_090_),
    .Z(_126_));
 INV_X1 _338_ (.A(_126_),
    .ZN(_127_));
 MUX2_X1 _339_ (.A(net7),
    .B(net25),
    .S(_089_),
    .Z(_128_));
 INV_X1 _340_ (.A(_128_),
    .ZN(_129_));
 OAI22_X1 _341_ (.A1(_094_),
    .A2(_127_),
    .B1(_129_),
    .B2(_095_),
    .ZN(_024_));
 MUX2_X1 _342_ (.A(net26),
    .B(net11),
    .S(_159_),
    .Z(_130_));
 INV_X1 _343_ (.A(_130_),
    .ZN(_131_));
 MUX2_X1 _344_ (.A(net3),
    .B(net20),
    .S(_158_),
    .Z(_132_));
 INV_X1 _345_ (.A(_132_),
    .ZN(_133_));
 OAI22_X1 _346_ (.A1(_164_),
    .A2(_131_),
    .B1(_133_),
    .B2(_165_),
    .ZN(_025_));
 MUX2_X1 _347_ (.A(net27),
    .B(net13),
    .S(_159_),
    .Z(_134_));
 INV_X1 _348_ (.A(_134_),
    .ZN(_135_));
 MUX2_X1 _349_ (.A(net4),
    .B(net21),
    .S(_158_),
    .Z(_136_));
 INV_X1 _350_ (.A(_136_),
    .ZN(_137_));
 OAI22_X1 _351_ (.A1(_164_),
    .A2(_135_),
    .B1(_137_),
    .B2(_165_),
    .ZN(_026_));
 MUX2_X1 _352_ (.A(net28),
    .B(net14),
    .S(_159_),
    .Z(_138_));
 INV_X1 _353_ (.A(_138_),
    .ZN(_139_));
 MUX2_X1 _354_ (.A(net5),
    .B(net22),
    .S(_158_),
    .Z(_140_));
 INV_X1 _355_ (.A(_140_),
    .ZN(_141_));
 OAI22_X1 _356_ (.A1(_164_),
    .A2(_139_),
    .B1(_141_),
    .B2(_165_),
    .ZN(_027_));
 MUX2_X1 _357_ (.A(net29),
    .B(net15),
    .S(_159_),
    .Z(_142_));
 INV_X1 _358_ (.A(_142_),
    .ZN(_143_));
 MUX2_X1 _359_ (.A(net6),
    .B(net24),
    .S(_158_),
    .Z(_144_));
 INV_X1 _360_ (.A(_144_),
    .ZN(_145_));
 OAI22_X1 _361_ (.A1(_164_),
    .A2(_143_),
    .B1(_145_),
    .B2(_165_),
    .ZN(_028_));
 MUX2_X1 _362_ (.A(net30),
    .B(net16),
    .S(_159_),
    .Z(_146_));
 INV_X1 _363_ (.A(_146_),
    .ZN(_147_));
 MUX2_X1 _364_ (.A(net7),
    .B(net25),
    .S(_158_),
    .Z(_148_));
 INV_X1 _365_ (.A(_148_),
    .ZN(_149_));
 OAI22_X1 _366_ (.A1(_164_),
    .A2(_147_),
    .B1(_149_),
    .B2(_165_),
    .ZN(_029_));
 MUX2_X1 _367_ (.A(net1),
    .B(net8),
    .S(_169_),
    .Z(_150_));
 INV_X1 _368_ (.A(_150_),
    .ZN(_151_));
 MUX2_X1 _369_ (.A(net31),
    .B(net17),
    .S(_168_),
    .Z(_152_));
 INV_X1 _370_ (.A(_152_),
    .ZN(_153_));
 OAI22_X1 _371_ (.A1(_173_),
    .A2(_151_),
    .B1(_153_),
    .B2(_174_),
    .ZN(_030_));
 MUX2_X1 _372_ (.A(net12),
    .B(net9),
    .S(_169_),
    .Z(_154_));
 INV_X1 _373_ (.A(_154_),
    .ZN(_155_));
 MUX2_X1 _374_ (.A(net32),
    .B(net18),
    .S(_168_),
    .Z(_156_));
 INV_X1 _375_ (.A(_156_),
    .ZN(_157_));
 OAI22_X1 _376_ (.A1(_173_),
    .A2(_155_),
    .B1(_157_),
    .B2(_174_),
    .ZN(_031_));
 BUF_X8 _377_ (.A(select[1]),
    .Z(_158_));
 BUF_X8 _378_ (.A(_158_),
    .Z(_159_));
 MUX2_X1 _379_ (.A(net1),
    .B(net8),
    .S(_159_),
    .Z(_160_));
 INV_X1 _380_ (.A(_160_),
    .ZN(_161_));
 INV_X1 _381_ (.A(net33),
    .ZN(_162_));
 BUF_X8 _382_ (.A(rst_n),
    .Z(_163_));
 NAND2_X4 _383_ (.A1(_162_),
    .A2(_163_),
    .ZN(_164_));
 NAND2_X4 _384_ (.A1(net33),
    .A2(_163_),
    .ZN(_165_));
 MUX2_X1 _385_ (.A(net31),
    .B(net17),
    .S(_158_),
    .Z(_166_));
 INV_X1 _386_ (.A(_166_),
    .ZN(_167_));
 OAI22_X1 _387_ (.A1(_161_),
    .A2(_164_),
    .B1(_165_),
    .B2(_167_),
    .ZN(_000_));
 BUF_X8 _388_ (.A(select[3]),
    .Z(_168_));
 BUF_X8 _389_ (.A(_168_),
    .Z(_169_));
 MUX2_X1 _390_ (.A(net23),
    .B(net10),
    .S(_169_),
    .Z(_170_));
 INV_X1 _391_ (.A(_170_),
    .ZN(_171_));
 INV_X1 _392_ (.A(net34),
    .ZN(_172_));
 NAND2_X4 _393_ (.A1(_172_),
    .A2(_163_),
    .ZN(_173_));
 DFF_X1 \data_out[0]$_SDFF_PN0_  (.D(_000_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net37),
    .QN(_212_));
 DFF_X1 \data_out[10]$_SDFF_PN0_  (.D(_001_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net38),
    .QN(_211_));
 DFF_X1 \data_out[11]$_SDFF_PN0_  (.D(_002_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net39),
    .QN(_210_));
 DFF_X1 \data_out[12]$_SDFF_PN0_  (.D(_003_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net40),
    .QN(_209_));
 DFF_X1 \data_out[13]$_SDFF_PN0_  (.D(_004_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net41),
    .QN(_208_));
 DFF_X1 \data_out[14]$_SDFF_PN0_  (.D(_005_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net42),
    .QN(_207_));
 DFF_X1 \data_out[15]$_SDFF_PN0_  (.D(_006_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net43),
    .QN(_206_));
 DFF_X1 \data_out[16]$_SDFF_PN0_  (.D(_007_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net44),
    .QN(_205_));
 DFF_X1 \data_out[17]$_SDFF_PN0_  (.D(_008_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net45),
    .QN(_204_));
 DFF_X1 \data_out[18]$_SDFF_PN0_  (.D(_009_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net46),
    .QN(_203_));
 DFF_X1 \data_out[19]$_SDFF_PN0_  (.D(_010_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net47),
    .QN(_202_));
 DFF_X1 \data_out[1]$_SDFF_PN0_  (.D(_011_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net48),
    .QN(_201_));
 DFF_X1 \data_out[20]$_SDFF_PN0_  (.D(_012_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net49),
    .QN(_200_));
 DFF_X1 \data_out[21]$_SDFF_PN0_  (.D(_013_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net50),
    .QN(_199_));
 DFF_X1 \data_out[22]$_SDFF_PN0_  (.D(_014_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net51),
    .QN(_198_));
 DFF_X1 \data_out[23]$_SDFF_PN0_  (.D(_015_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net52),
    .QN(_197_));
 DFF_X1 \data_out[24]$_SDFF_PN0_  (.D(_016_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net53),
    .QN(_196_));
 DFF_X1 \data_out[25]$_SDFF_PN0_  (.D(_017_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net54),
    .QN(_195_));
 DFF_X1 \data_out[26]$_SDFF_PN0_  (.D(_018_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net55),
    .QN(_194_));
 DFF_X1 \data_out[27]$_SDFF_PN0_  (.D(_019_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net56),
    .QN(_193_));
 DFF_X1 \data_out[28]$_SDFF_PN0_  (.D(_020_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net57),
    .QN(_192_));
 DFF_X1 \data_out[29]$_SDFF_PN0_  (.D(_021_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net58),
    .QN(_191_));
 DFF_X1 \data_out[2]$_SDFF_PN0_  (.D(_022_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net59),
    .QN(_190_));
 DFF_X1 \data_out[30]$_SDFF_PN0_  (.D(_023_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net60),
    .QN(_189_));
 DFF_X1 \data_out[31]$_SDFF_PN0_  (.D(_024_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net61),
    .QN(_188_));
 DFF_X1 \data_out[3]$_SDFF_PN0_  (.D(_025_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net62),
    .QN(_187_));
 DFF_X1 \data_out[4]$_SDFF_PN0_  (.D(_026_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net63),
    .QN(_186_));
 DFF_X1 \data_out[5]$_SDFF_PN0_  (.D(_027_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net64),
    .QN(_185_));
 DFF_X1 \data_out[6]$_SDFF_PN0_  (.D(_028_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net65),
    .QN(_184_));
 DFF_X1 \data_out[7]$_SDFF_PN0_  (.D(_029_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net66),
    .QN(_183_));
 DFF_X1 \data_out[8]$_SDFF_PN0_  (.D(_030_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net67),
    .QN(_182_));
 DFF_X1 \data_out[9]$_SDFF_PN0_  (.D(_031_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net68),
    .QN(_181_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_61 ();
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[10]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[11]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[12]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[13]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[14]),
    .Z(net6));
 BUF_X1 input7 (.A(data_in[15]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[16]),
    .Z(net8));
 BUF_X1 input9 (.A(data_in[17]),
    .Z(net9));
 BUF_X1 input10 (.A(data_in[18]),
    .Z(net10));
 BUF_X1 input11 (.A(data_in[19]),
    .Z(net11));
 BUF_X1 input12 (.A(data_in[1]),
    .Z(net12));
 BUF_X1 input13 (.A(data_in[20]),
    .Z(net13));
 BUF_X1 input14 (.A(data_in[21]),
    .Z(net14));
 BUF_X1 input15 (.A(data_in[22]),
    .Z(net15));
 BUF_X1 input16 (.A(data_in[23]),
    .Z(net16));
 BUF_X1 input17 (.A(data_in[24]),
    .Z(net17));
 BUF_X1 input18 (.A(data_in[25]),
    .Z(net18));
 BUF_X1 input19 (.A(data_in[26]),
    .Z(net19));
 BUF_X1 input20 (.A(data_in[27]),
    .Z(net20));
 BUF_X1 input21 (.A(data_in[28]),
    .Z(net21));
 BUF_X1 input22 (.A(data_in[29]),
    .Z(net22));
 BUF_X1 input23 (.A(data_in[2]),
    .Z(net23));
 BUF_X1 input24 (.A(data_in[30]),
    .Z(net24));
 BUF_X1 input25 (.A(data_in[31]),
    .Z(net25));
 BUF_X1 input26 (.A(data_in[3]),
    .Z(net26));
 BUF_X1 input27 (.A(data_in[4]),
    .Z(net27));
 BUF_X1 input28 (.A(data_in[5]),
    .Z(net28));
 BUF_X1 input29 (.A(data_in[6]),
    .Z(net29));
 BUF_X1 input30 (.A(data_in[7]),
    .Z(net30));
 BUF_X1 input31 (.A(data_in[8]),
    .Z(net31));
 BUF_X1 input32 (.A(data_in[9]),
    .Z(net32));
 BUF_X1 input33 (.A(select[0]),
    .Z(net33));
 BUF_X1 input34 (.A(select[2]),
    .Z(net34));
 BUF_X1 input35 (.A(select[4]),
    .Z(net35));
 BUF_X1 input36 (.A(select[6]),
    .Z(net36));
 BUF_X1 output37 (.A(net37),
    .Z(data_out[0]));
 BUF_X1 output38 (.A(net38),
    .Z(data_out[10]));
 BUF_X1 output39 (.A(net39),
    .Z(data_out[11]));
 BUF_X1 output40 (.A(net40),
    .Z(data_out[12]));
 BUF_X1 output41 (.A(net41),
    .Z(data_out[13]));
 BUF_X1 output42 (.A(net42),
    .Z(data_out[14]));
 BUF_X1 output43 (.A(net43),
    .Z(data_out[15]));
 BUF_X1 output44 (.A(net44),
    .Z(data_out[16]));
 BUF_X1 output45 (.A(net45),
    .Z(data_out[17]));
 BUF_X1 output46 (.A(net46),
    .Z(data_out[18]));
 BUF_X1 output47 (.A(net47),
    .Z(data_out[19]));
 BUF_X1 output48 (.A(net48),
    .Z(data_out[1]));
 BUF_X1 output49 (.A(net49),
    .Z(data_out[20]));
 BUF_X1 output50 (.A(net50),
    .Z(data_out[21]));
 BUF_X1 output51 (.A(net51),
    .Z(data_out[22]));
 BUF_X1 output52 (.A(net52),
    .Z(data_out[23]));
 BUF_X1 output53 (.A(net53),
    .Z(data_out[24]));
 BUF_X1 output54 (.A(net54),
    .Z(data_out[25]));
 BUF_X1 output55 (.A(net55),
    .Z(data_out[26]));
 BUF_X1 output56 (.A(net56),
    .Z(data_out[27]));
 BUF_X1 output57 (.A(net57),
    .Z(data_out[28]));
 BUF_X1 output58 (.A(net58),
    .Z(data_out[29]));
 BUF_X1 output59 (.A(net59),
    .Z(data_out[2]));
 BUF_X1 output60 (.A(net60),
    .Z(data_out[30]));
 BUF_X1 output61 (.A(net61),
    .Z(data_out[31]));
 BUF_X1 output62 (.A(net62),
    .Z(data_out[3]));
 BUF_X1 output63 (.A(net63),
    .Z(data_out[4]));
 BUF_X1 output64 (.A(net64),
    .Z(data_out[5]));
 BUF_X1 output65 (.A(net65),
    .Z(data_out[6]));
 BUF_X1 output66 (.A(net66),
    .Z(data_out[7]));
 BUF_X1 output67 (.A(net67),
    .Z(data_out[8]));
 BUF_X1 output68 (.A(net68),
    .Z(data_out[9]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X1 clkload0 (.A(clknet_2_0__leaf_clk));
 CLKBUF_X1 clkload1 (.A(clknet_2_2__leaf_clk));
 CLKBUF_X1 clkload2 (.A(clknet_2_3__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X16 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_49 ();
 FILLCELL_X4 FILLER_0_57 ();
 FILLCELL_X1 FILLER_0_61 ();
 FILLCELL_X16 FILLER_0_68 ();
 FILLCELL_X4 FILLER_0_84 ();
 FILLCELL_X1 FILLER_0_88 ();
 FILLCELL_X2 FILLER_0_95 ();
 FILLCELL_X1 FILLER_0_97 ();
 FILLCELL_X8 FILLER_0_101 ();
 FILLCELL_X2 FILLER_0_118 ();
 FILLCELL_X1 FILLER_0_120 ();
 FILLCELL_X8 FILLER_0_130 ();
 FILLCELL_X4 FILLER_0_138 ();
 FILLCELL_X2 FILLER_0_145 ();
 FILLCELL_X1 FILLER_0_150 ();
 FILLCELL_X8 FILLER_0_154 ();
 FILLCELL_X4 FILLER_0_162 ();
 FILLCELL_X2 FILLER_0_166 ();
 FILLCELL_X16 FILLER_0_171 ();
 FILLCELL_X2 FILLER_0_187 ();
 FILLCELL_X32 FILLER_0_192 ();
 FILLCELL_X4 FILLER_0_224 ();
 FILLCELL_X2 FILLER_0_228 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X8 FILLER_1_65 ();
 FILLCELL_X4 FILLER_1_73 ();
 FILLCELL_X2 FILLER_1_77 ();
 FILLCELL_X8 FILLER_1_82 ();
 FILLCELL_X2 FILLER_1_90 ();
 FILLCELL_X1 FILLER_1_92 ();
 FILLCELL_X16 FILLER_1_110 ();
 FILLCELL_X1 FILLER_1_126 ();
 FILLCELL_X8 FILLER_1_144 ();
 FILLCELL_X4 FILLER_1_152 ();
 FILLCELL_X2 FILLER_1_173 ();
 FILLCELL_X1 FILLER_1_175 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X4 FILLER_1_225 ();
 FILLCELL_X1 FILLER_1_229 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X2 FILLER_2_65 ();
 FILLCELL_X8 FILLER_2_101 ();
 FILLCELL_X4 FILLER_2_109 ();
 FILLCELL_X32 FILLER_2_130 ();
 FILLCELL_X32 FILLER_2_162 ();
 FILLCELL_X32 FILLER_2_194 ();
 FILLCELL_X4 FILLER_2_226 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X16 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_49 ();
 FILLCELL_X4 FILLER_3_57 ();
 FILLCELL_X1 FILLER_3_61 ();
 FILLCELL_X8 FILLER_3_71 ();
 FILLCELL_X2 FILLER_3_79 ();
 FILLCELL_X1 FILLER_3_81 ();
 FILLCELL_X32 FILLER_3_91 ();
 FILLCELL_X32 FILLER_3_123 ();
 FILLCELL_X1 FILLER_3_155 ();
 FILLCELL_X8 FILLER_3_163 ();
 FILLCELL_X1 FILLER_3_171 ();
 FILLCELL_X32 FILLER_3_174 ();
 FILLCELL_X16 FILLER_3_206 ();
 FILLCELL_X8 FILLER_3_222 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X4 FILLER_4_65 ();
 FILLCELL_X4 FILLER_4_74 ();
 FILLCELL_X1 FILLER_4_78 ();
 FILLCELL_X2 FILLER_4_88 ();
 FILLCELL_X1 FILLER_4_95 ();
 FILLCELL_X8 FILLER_4_98 ();
 FILLCELL_X4 FILLER_4_106 ();
 FILLCELL_X2 FILLER_4_110 ();
 FILLCELL_X1 FILLER_4_112 ();
 FILLCELL_X4 FILLER_4_122 ();
 FILLCELL_X16 FILLER_4_133 ();
 FILLCELL_X1 FILLER_4_156 ();
 FILLCELL_X8 FILLER_4_164 ();
 FILLCELL_X2 FILLER_4_172 ();
 FILLCELL_X1 FILLER_4_179 ();
 FILLCELL_X32 FILLER_4_182 ();
 FILLCELL_X16 FILLER_4_214 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X16 FILLER_5_65 ();
 FILLCELL_X8 FILLER_5_81 ();
 FILLCELL_X1 FILLER_5_89 ();
 FILLCELL_X16 FILLER_5_97 ();
 FILLCELL_X8 FILLER_5_113 ();
 FILLCELL_X2 FILLER_5_121 ();
 FILLCELL_X1 FILLER_5_123 ();
 FILLCELL_X32 FILLER_5_131 ();
 FILLCELL_X4 FILLER_5_163 ();
 FILLCELL_X2 FILLER_5_167 ();
 FILLCELL_X1 FILLER_5_171 ();
 FILLCELL_X32 FILLER_5_186 ();
 FILLCELL_X8 FILLER_5_218 ();
 FILLCELL_X4 FILLER_5_226 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X4 FILLER_6_65 ();
 FILLCELL_X1 FILLER_6_76 ();
 FILLCELL_X32 FILLER_6_86 ();
 FILLCELL_X16 FILLER_6_132 ();
 FILLCELL_X1 FILLER_6_148 ();
 FILLCELL_X4 FILLER_6_163 ();
 FILLCELL_X1 FILLER_6_167 ();
 FILLCELL_X32 FILLER_6_170 ();
 FILLCELL_X4 FILLER_6_202 ();
 FILLCELL_X2 FILLER_6_206 ();
 FILLCELL_X16 FILLER_6_211 ();
 FILLCELL_X2 FILLER_6_227 ();
 FILLCELL_X1 FILLER_6_229 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_65 ();
 FILLCELL_X2 FILLER_7_73 ();
 FILLCELL_X4 FILLER_7_77 ();
 FILLCELL_X1 FILLER_7_81 ();
 FILLCELL_X8 FILLER_7_105 ();
 FILLCELL_X4 FILLER_7_113 ();
 FILLCELL_X2 FILLER_7_117 ();
 FILLCELL_X8 FILLER_7_121 ();
 FILLCELL_X32 FILLER_7_134 ();
 FILLCELL_X4 FILLER_7_166 ();
 FILLCELL_X2 FILLER_7_170 ();
 FILLCELL_X2 FILLER_7_195 ();
 FILLCELL_X4 FILLER_7_200 ();
 FILLCELL_X2 FILLER_7_221 ();
 FILLCELL_X1 FILLER_7_223 ();
 FILLCELL_X2 FILLER_7_227 ();
 FILLCELL_X1 FILLER_7_229 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X8 FILLER_8_65 ();
 FILLCELL_X4 FILLER_8_73 ();
 FILLCELL_X16 FILLER_8_82 ();
 FILLCELL_X8 FILLER_8_98 ();
 FILLCELL_X4 FILLER_8_106 ();
 FILLCELL_X2 FILLER_8_110 ();
 FILLCELL_X1 FILLER_8_112 ();
 FILLCELL_X2 FILLER_8_120 ();
 FILLCELL_X1 FILLER_8_122 ();
 FILLCELL_X32 FILLER_8_139 ();
 FILLCELL_X16 FILLER_8_171 ();
 FILLCELL_X2 FILLER_8_187 ();
 FILLCELL_X4 FILLER_8_213 ();
 FILLCELL_X1 FILLER_8_217 ();
 FILLCELL_X8 FILLER_8_221 ();
 FILLCELL_X1 FILLER_8_229 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X2 FILLER_9_17 ();
 FILLCELL_X1 FILLER_9_19 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X8 FILLER_9_49 ();
 FILLCELL_X2 FILLER_9_57 ();
 FILLCELL_X32 FILLER_9_76 ();
 FILLCELL_X16 FILLER_9_108 ();
 FILLCELL_X8 FILLER_9_124 ();
 FILLCELL_X4 FILLER_9_132 ();
 FILLCELL_X2 FILLER_9_136 ();
 FILLCELL_X32 FILLER_9_140 ();
 FILLCELL_X4 FILLER_9_172 ();
 FILLCELL_X2 FILLER_9_176 ();
 FILLCELL_X1 FILLER_9_178 ();
 FILLCELL_X32 FILLER_9_184 ();
 FILLCELL_X8 FILLER_9_216 ();
 FILLCELL_X4 FILLER_9_224 ();
 FILLCELL_X2 FILLER_9_228 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X2 FILLER_10_9 ();
 FILLCELL_X32 FILLER_10_14 ();
 FILLCELL_X32 FILLER_10_46 ();
 FILLCELL_X16 FILLER_10_78 ();
 FILLCELL_X1 FILLER_10_127 ();
 FILLCELL_X2 FILLER_10_132 ();
 FILLCELL_X32 FILLER_10_139 ();
 FILLCELL_X2 FILLER_10_171 ();
 FILLCELL_X1 FILLER_10_173 ();
 FILLCELL_X2 FILLER_10_179 ();
 FILLCELL_X1 FILLER_10_181 ();
 FILLCELL_X8 FILLER_10_184 ();
 FILLCELL_X2 FILLER_10_192 ();
 FILLCELL_X4 FILLER_10_211 ();
 FILLCELL_X2 FILLER_10_215 ();
 FILLCELL_X1 FILLER_10_217 ();
 FILLCELL_X8 FILLER_10_221 ();
 FILLCELL_X1 FILLER_10_229 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X16 FILLER_11_97 ();
 FILLCELL_X4 FILLER_11_113 ();
 FILLCELL_X1 FILLER_11_126 ();
 FILLCELL_X16 FILLER_11_132 ();
 FILLCELL_X4 FILLER_11_148 ();
 FILLCELL_X2 FILLER_11_152 ();
 FILLCELL_X1 FILLER_11_154 ();
 FILLCELL_X2 FILLER_11_174 ();
 FILLCELL_X8 FILLER_11_192 ();
 FILLCELL_X4 FILLER_11_203 ();
 FILLCELL_X2 FILLER_11_224 ();
 FILLCELL_X1 FILLER_11_226 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_20 ();
 FILLCELL_X2 FILLER_12_24 ();
 FILLCELL_X1 FILLER_12_26 ();
 FILLCELL_X16 FILLER_12_40 ();
 FILLCELL_X4 FILLER_12_56 ();
 FILLCELL_X32 FILLER_12_71 ();
 FILLCELL_X32 FILLER_12_103 ();
 FILLCELL_X16 FILLER_12_135 ();
 FILLCELL_X8 FILLER_12_151 ();
 FILLCELL_X4 FILLER_12_159 ();
 FILLCELL_X1 FILLER_12_163 ();
 FILLCELL_X2 FILLER_12_178 ();
 FILLCELL_X1 FILLER_12_187 ();
 FILLCELL_X8 FILLER_12_200 ();
 FILLCELL_X16 FILLER_12_211 ();
 FILLCELL_X2 FILLER_12_227 ();
 FILLCELL_X1 FILLER_12_229 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_9 ();
 FILLCELL_X16 FILLER_13_17 ();
 FILLCELL_X2 FILLER_13_33 ();
 FILLCELL_X1 FILLER_13_35 ();
 FILLCELL_X32 FILLER_13_74 ();
 FILLCELL_X16 FILLER_13_106 ();
 FILLCELL_X2 FILLER_13_122 ();
 FILLCELL_X1 FILLER_13_124 ();
 FILLCELL_X16 FILLER_13_142 ();
 FILLCELL_X4 FILLER_13_158 ();
 FILLCELL_X2 FILLER_13_162 ();
 FILLCELL_X1 FILLER_13_164 ();
 FILLCELL_X4 FILLER_13_172 ();
 FILLCELL_X1 FILLER_13_176 ();
 FILLCELL_X4 FILLER_13_186 ();
 FILLCELL_X1 FILLER_13_190 ();
 FILLCELL_X4 FILLER_13_196 ();
 FILLCELL_X2 FILLER_13_217 ();
 FILLCELL_X1 FILLER_13_219 ();
 FILLCELL_X4 FILLER_13_223 ();
 FILLCELL_X2 FILLER_13_227 ();
 FILLCELL_X1 FILLER_13_229 ();
 FILLCELL_X1 FILLER_14_14 ();
 FILLCELL_X16 FILLER_14_18 ();
 FILLCELL_X4 FILLER_14_34 ();
 FILLCELL_X1 FILLER_14_38 ();
 FILLCELL_X8 FILLER_14_59 ();
 FILLCELL_X1 FILLER_14_67 ();
 FILLCELL_X16 FILLER_14_79 ();
 FILLCELL_X2 FILLER_14_95 ();
 FILLCELL_X16 FILLER_14_123 ();
 FILLCELL_X1 FILLER_14_139 ();
 FILLCELL_X16 FILLER_14_145 ();
 FILLCELL_X2 FILLER_14_168 ();
 FILLCELL_X8 FILLER_14_172 ();
 FILLCELL_X2 FILLER_14_190 ();
 FILLCELL_X2 FILLER_14_209 ();
 FILLCELL_X1 FILLER_14_211 ();
 FILLCELL_X8 FILLER_14_215 ();
 FILLCELL_X4 FILLER_14_223 ();
 FILLCELL_X2 FILLER_14_227 ();
 FILLCELL_X1 FILLER_14_229 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X4 FILLER_15_17 ();
 FILLCELL_X1 FILLER_15_21 ();
 FILLCELL_X32 FILLER_15_35 ();
 FILLCELL_X32 FILLER_15_67 ();
 FILLCELL_X32 FILLER_15_99 ();
 FILLCELL_X16 FILLER_15_131 ();
 FILLCELL_X8 FILLER_15_147 ();
 FILLCELL_X1 FILLER_15_155 ();
 FILLCELL_X32 FILLER_15_173 ();
 FILLCELL_X16 FILLER_15_205 ();
 FILLCELL_X2 FILLER_15_221 ();
 FILLCELL_X1 FILLER_15_223 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X16 FILLER_16_161 ();
 FILLCELL_X8 FILLER_16_177 ();
 FILLCELL_X2 FILLER_16_185 ();
 FILLCELL_X1 FILLER_16_187 ();
 FILLCELL_X16 FILLER_16_208 ();
 FILLCELL_X4 FILLER_16_224 ();
 FILLCELL_X2 FILLER_16_228 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_9 ();
 FILLCELL_X16 FILLER_17_16 ();
 FILLCELL_X8 FILLER_17_32 ();
 FILLCELL_X1 FILLER_17_40 ();
 FILLCELL_X2 FILLER_17_48 ();
 FILLCELL_X1 FILLER_17_50 ();
 FILLCELL_X16 FILLER_17_70 ();
 FILLCELL_X8 FILLER_17_86 ();
 FILLCELL_X2 FILLER_17_94 ();
 FILLCELL_X8 FILLER_17_98 ();
 FILLCELL_X4 FILLER_17_106 ();
 FILLCELL_X2 FILLER_17_110 ();
 FILLCELL_X16 FILLER_17_119 ();
 FILLCELL_X8 FILLER_17_135 ();
 FILLCELL_X4 FILLER_17_143 ();
 FILLCELL_X1 FILLER_17_147 ();
 FILLCELL_X16 FILLER_17_157 ();
 FILLCELL_X8 FILLER_17_182 ();
 FILLCELL_X4 FILLER_17_207 ();
 FILLCELL_X1 FILLER_17_211 ();
 FILLCELL_X8 FILLER_17_218 ();
 FILLCELL_X4 FILLER_17_226 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_9 ();
 FILLCELL_X8 FILLER_18_14 ();
 FILLCELL_X4 FILLER_18_22 ();
 FILLCELL_X2 FILLER_18_26 ();
 FILLCELL_X1 FILLER_18_28 ();
 FILLCELL_X4 FILLER_18_39 ();
 FILLCELL_X1 FILLER_18_50 ();
 FILLCELL_X4 FILLER_18_53 ();
 FILLCELL_X2 FILLER_18_57 ();
 FILLCELL_X1 FILLER_18_59 ();
 FILLCELL_X8 FILLER_18_76 ();
 FILLCELL_X4 FILLER_18_84 ();
 FILLCELL_X1 FILLER_18_88 ();
 FILLCELL_X1 FILLER_18_103 ();
 FILLCELL_X2 FILLER_18_106 ();
 FILLCELL_X8 FILLER_18_115 ();
 FILLCELL_X4 FILLER_18_123 ();
 FILLCELL_X2 FILLER_18_127 ();
 FILLCELL_X1 FILLER_18_129 ();
 FILLCELL_X2 FILLER_18_146 ();
 FILLCELL_X4 FILLER_18_162 ();
 FILLCELL_X2 FILLER_18_166 ();
 FILLCELL_X4 FILLER_18_196 ();
 FILLCELL_X2 FILLER_18_200 ();
 FILLCELL_X1 FILLER_18_202 ();
 FILLCELL_X2 FILLER_18_206 ();
 FILLCELL_X1 FILLER_18_208 ();
 FILLCELL_X8 FILLER_18_212 ();
 FILLCELL_X4 FILLER_18_220 ();
 FILLCELL_X1 FILLER_18_224 ();
 FILLCELL_X2 FILLER_18_228 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X16 FILLER_19_33 ();
 FILLCELL_X8 FILLER_19_49 ();
 FILLCELL_X4 FILLER_19_57 ();
 FILLCELL_X2 FILLER_19_61 ();
 FILLCELL_X32 FILLER_19_68 ();
 FILLCELL_X4 FILLER_19_100 ();
 FILLCELL_X2 FILLER_19_104 ();
 FILLCELL_X1 FILLER_19_106 ();
 FILLCELL_X32 FILLER_19_121 ();
 FILLCELL_X1 FILLER_19_153 ();
 FILLCELL_X16 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_177 ();
 FILLCELL_X1 FILLER_19_181 ();
 FILLCELL_X4 FILLER_19_184 ();
 FILLCELL_X1 FILLER_19_193 ();
 FILLCELL_X4 FILLER_19_196 ();
 FILLCELL_X2 FILLER_19_200 ();
 FILLCELL_X16 FILLER_19_205 ();
 FILLCELL_X8 FILLER_19_221 ();
 FILLCELL_X1 FILLER_19_229 ();
 FILLCELL_X16 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_17 ();
 FILLCELL_X2 FILLER_20_21 ();
 FILLCELL_X1 FILLER_20_23 ();
 FILLCELL_X4 FILLER_20_37 ();
 FILLCELL_X2 FILLER_20_41 ();
 FILLCELL_X2 FILLER_20_50 ();
 FILLCELL_X8 FILLER_20_59 ();
 FILLCELL_X1 FILLER_20_67 ();
 FILLCELL_X8 FILLER_20_75 ();
 FILLCELL_X2 FILLER_20_83 ();
 FILLCELL_X32 FILLER_20_92 ();
 FILLCELL_X8 FILLER_20_124 ();
 FILLCELL_X2 FILLER_20_132 ();
 FILLCELL_X4 FILLER_20_148 ();
 FILLCELL_X1 FILLER_20_152 ();
 FILLCELL_X2 FILLER_20_160 ();
 FILLCELL_X1 FILLER_20_162 ();
 FILLCELL_X16 FILLER_20_178 ();
 FILLCELL_X8 FILLER_20_194 ();
 FILLCELL_X4 FILLER_20_202 ();
 FILLCELL_X2 FILLER_20_209 ();
 FILLCELL_X2 FILLER_20_228 ();
 FILLCELL_X1 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_5 ();
 FILLCELL_X4 FILLER_21_13 ();
 FILLCELL_X1 FILLER_21_17 ();
 FILLCELL_X16 FILLER_21_21 ();
 FILLCELL_X4 FILLER_21_37 ();
 FILLCELL_X2 FILLER_21_41 ();
 FILLCELL_X1 FILLER_21_50 ();
 FILLCELL_X16 FILLER_21_57 ();
 FILLCELL_X1 FILLER_21_73 ();
 FILLCELL_X16 FILLER_21_76 ();
 FILLCELL_X2 FILLER_21_92 ();
 FILLCELL_X2 FILLER_21_103 ();
 FILLCELL_X4 FILLER_21_114 ();
 FILLCELL_X2 FILLER_21_118 ();
 FILLCELL_X2 FILLER_21_128 ();
 FILLCELL_X2 FILLER_21_137 ();
 FILLCELL_X1 FILLER_21_139 ();
 FILLCELL_X8 FILLER_21_142 ();
 FILLCELL_X8 FILLER_21_152 ();
 FILLCELL_X4 FILLER_21_160 ();
 FILLCELL_X2 FILLER_21_164 ();
 FILLCELL_X1 FILLER_21_175 ();
 FILLCELL_X16 FILLER_21_196 ();
 FILLCELL_X8 FILLER_21_212 ();
 FILLCELL_X4 FILLER_21_220 ();
 FILLCELL_X2 FILLER_21_224 ();
 FILLCELL_X1 FILLER_21_226 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X16 FILLER_22_33 ();
 FILLCELL_X4 FILLER_22_49 ();
 FILLCELL_X8 FILLER_22_58 ();
 FILLCELL_X2 FILLER_22_66 ();
 FILLCELL_X16 FILLER_22_73 ();
 FILLCELL_X4 FILLER_22_89 ();
 FILLCELL_X2 FILLER_22_93 ();
 FILLCELL_X4 FILLER_22_100 ();
 FILLCELL_X2 FILLER_22_104 ();
 FILLCELL_X1 FILLER_22_115 ();
 FILLCELL_X16 FILLER_22_118 ();
 FILLCELL_X2 FILLER_22_136 ();
 FILLCELL_X1 FILLER_22_138 ();
 FILLCELL_X4 FILLER_22_141 ();
 FILLCELL_X2 FILLER_22_145 ();
 FILLCELL_X16 FILLER_22_152 ();
 FILLCELL_X4 FILLER_22_168 ();
 FILLCELL_X2 FILLER_22_172 ();
 FILLCELL_X1 FILLER_22_174 ();
 FILLCELL_X4 FILLER_22_185 ();
 FILLCELL_X2 FILLER_22_189 ();
 FILLCELL_X16 FILLER_22_208 ();
 FILLCELL_X2 FILLER_22_224 ();
 FILLCELL_X1 FILLER_22_229 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X8 FILLER_23_97 ();
 FILLCELL_X2 FILLER_23_105 ();
 FILLCELL_X1 FILLER_23_107 ();
 FILLCELL_X16 FILLER_23_113 ();
 FILLCELL_X4 FILLER_23_129 ();
 FILLCELL_X2 FILLER_23_133 ();
 FILLCELL_X32 FILLER_23_140 ();
 FILLCELL_X8 FILLER_23_172 ();
 FILLCELL_X4 FILLER_23_180 ();
 FILLCELL_X2 FILLER_23_184 ();
 FILLCELL_X16 FILLER_23_203 ();
 FILLCELL_X8 FILLER_23_219 ();
 FILLCELL_X2 FILLER_23_227 ();
 FILLCELL_X1 FILLER_23_229 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X16 FILLER_24_33 ();
 FILLCELL_X2 FILLER_24_49 ();
 FILLCELL_X32 FILLER_24_85 ();
 FILLCELL_X32 FILLER_24_117 ();
 FILLCELL_X1 FILLER_24_149 ();
 FILLCELL_X32 FILLER_24_167 ();
 FILLCELL_X4 FILLER_24_199 ();
 FILLCELL_X1 FILLER_24_203 ();
 FILLCELL_X16 FILLER_24_207 ();
 FILLCELL_X4 FILLER_24_223 ();
 FILLCELL_X2 FILLER_24_227 ();
 FILLCELL_X1 FILLER_24_229 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X16 FILLER_25_65 ();
 FILLCELL_X8 FILLER_25_81 ();
 FILLCELL_X1 FILLER_25_89 ();
 FILLCELL_X32 FILLER_25_124 ();
 FILLCELL_X32 FILLER_25_156 ();
 FILLCELL_X32 FILLER_25_188 ();
 FILLCELL_X8 FILLER_25_220 ();
 FILLCELL_X2 FILLER_25_228 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X16 FILLER_26_33 ();
 FILLCELL_X8 FILLER_26_49 ();
 FILLCELL_X2 FILLER_26_57 ();
 FILLCELL_X1 FILLER_26_59 ();
 FILLCELL_X32 FILLER_26_77 ();
 FILLCELL_X4 FILLER_26_126 ();
 FILLCELL_X2 FILLER_26_130 ();
 FILLCELL_X1 FILLER_26_132 ();
 FILLCELL_X32 FILLER_26_167 ();
 FILLCELL_X16 FILLER_26_199 ();
 FILLCELL_X8 FILLER_26_215 ();
 FILLCELL_X4 FILLER_26_223 ();
 FILLCELL_X2 FILLER_26_227 ();
 FILLCELL_X1 FILLER_26_229 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X4 FILLER_27_225 ();
 FILLCELL_X1 FILLER_27_229 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X4 FILLER_28_225 ();
 FILLCELL_X1 FILLER_28_229 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X16 FILLER_29_65 ();
 FILLCELL_X2 FILLER_29_81 ();
 FILLCELL_X1 FILLER_29_83 ();
 FILLCELL_X16 FILLER_29_87 ();
 FILLCELL_X2 FILLER_29_103 ();
 FILLCELL_X32 FILLER_29_114 ();
 FILLCELL_X32 FILLER_29_146 ();
 FILLCELL_X32 FILLER_29_178 ();
 FILLCELL_X16 FILLER_29_210 ();
 FILLCELL_X4 FILLER_29_226 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X1 FILLER_30_65 ();
 FILLCELL_X4 FILLER_30_69 ();
 FILLCELL_X2 FILLER_30_73 ();
 FILLCELL_X4 FILLER_30_78 ();
 FILLCELL_X1 FILLER_30_82 ();
 FILLCELL_X2 FILLER_30_86 ();
 FILLCELL_X16 FILLER_30_91 ();
 FILLCELL_X8 FILLER_30_107 ();
 FILLCELL_X4 FILLER_30_115 ();
 FILLCELL_X2 FILLER_30_122 ();
 FILLCELL_X4 FILLER_30_127 ();
 FILLCELL_X1 FILLER_30_131 ();
 FILLCELL_X2 FILLER_30_138 ();
 FILLCELL_X4 FILLER_30_143 ();
 FILLCELL_X2 FILLER_30_147 ();
 FILLCELL_X1 FILLER_30_149 ();
 FILLCELL_X8 FILLER_30_153 ();
 FILLCELL_X4 FILLER_30_161 ();
 FILLCELL_X2 FILLER_30_168 ();
 FILLCELL_X32 FILLER_30_173 ();
 FILLCELL_X16 FILLER_30_205 ();
 FILLCELL_X8 FILLER_30_221 ();
 FILLCELL_X1 FILLER_30_229 ();
endmodule
