module network_interface_cdc (dst_clk,
    dst_rst_n,
    mem_read,
    mem_ready,
    mem_write,
    router_in_ready,
    router_in_valid,
    router_out_ready,
    router_out_valid,
    src_clk,
    src_rst_n,
    dest_id,
    mem_addr,
    mem_rdata,
    mem_wdata,
    msg_type,
    router_in_data,
    router_out_data);
 input dst_clk;
 input dst_rst_n;
 input mem_read;
 output mem_ready;
 input mem_write;
 input router_in_ready;
 output router_in_valid;
 output router_out_ready;
 input router_out_valid;
 input src_clk;
 input src_rst_n;
 input [7:0] dest_id;
 input [31:0] mem_addr;
 output [31:0] mem_rdata;
 input [31:0] mem_wdata;
 input [2:0] msg_type;
 output [31:0] router_in_data;
 input [31:0] router_out_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire dst_ack;
 wire dst_ack_prev;
 wire dst_ack_sync;
 wire \dst_ack_sync_reg[0] ;
 wire dst_data_valid;
 wire dst_data_valid_sync;
 wire \dst_data_valid_sync_reg[0] ;
 wire dst_is_write_op;
 wire \dst_state[0] ;
 wire \dst_state[1] ;
 wire \dst_state[2] ;
 wire \dst_state[3] ;
 wire \dst_to_src_data[0] ;
 wire \dst_to_src_data[10] ;
 wire \dst_to_src_data[11] ;
 wire \dst_to_src_data[12] ;
 wire \dst_to_src_data[13] ;
 wire \dst_to_src_data[14] ;
 wire \dst_to_src_data[15] ;
 wire \dst_to_src_data[16] ;
 wire \dst_to_src_data[17] ;
 wire \dst_to_src_data[18] ;
 wire \dst_to_src_data[19] ;
 wire \dst_to_src_data[1] ;
 wire \dst_to_src_data[20] ;
 wire \dst_to_src_data[21] ;
 wire \dst_to_src_data[22] ;
 wire \dst_to_src_data[23] ;
 wire \dst_to_src_data[24] ;
 wire \dst_to_src_data[25] ;
 wire \dst_to_src_data[26] ;
 wire \dst_to_src_data[27] ;
 wire \dst_to_src_data[28] ;
 wire \dst_to_src_data[29] ;
 wire \dst_to_src_data[2] ;
 wire \dst_to_src_data[30] ;
 wire \dst_to_src_data[31] ;
 wire \dst_to_src_data[3] ;
 wire \dst_to_src_data[4] ;
 wire \dst_to_src_data[5] ;
 wire \dst_to_src_data[6] ;
 wire \dst_to_src_data[7] ;
 wire \dst_to_src_data[8] ;
 wire \dst_to_src_data[9] ;
 wire src_data_valid;
 wire src_data_valid_sync;
 wire \src_data_valid_sync_reg[0] ;
 wire src_is_write_op_flag;
 wire src_is_write_op_sync;
 wire \src_is_write_op_sync_reg[0] ;
 wire src_req;
 wire src_req_prev;
 wire src_req_sync;
 wire \src_req_sync_reg[0] ;
 wire \src_state[0] ;
 wire \src_state[1] ;
 wire \src_state[2] ;
 wire \src_state[3] ;
 wire \src_to_dst_data[0] ;
 wire \src_to_dst_data[10] ;
 wire \src_to_dst_data[11] ;
 wire \src_to_dst_data[12] ;
 wire \src_to_dst_data[13] ;
 wire \src_to_dst_data[14] ;
 wire \src_to_dst_data[15] ;
 wire \src_to_dst_data[16] ;
 wire \src_to_dst_data[17] ;
 wire \src_to_dst_data[18] ;
 wire \src_to_dst_data[19] ;
 wire \src_to_dst_data[1] ;
 wire \src_to_dst_data[20] ;
 wire \src_to_dst_data[21] ;
 wire \src_to_dst_data[22] ;
 wire \src_to_dst_data[23] ;
 wire \src_to_dst_data[24] ;
 wire \src_to_dst_data[25] ;
 wire \src_to_dst_data[26] ;
 wire \src_to_dst_data[27] ;
 wire \src_to_dst_data[28] ;
 wire \src_to_dst_data[29] ;
 wire \src_to_dst_data[2] ;
 wire \src_to_dst_data[30] ;
 wire \src_to_dst_data[31] ;
 wire \src_to_dst_data[3] ;
 wire \src_to_dst_data[4] ;
 wire \src_to_dst_data[5] ;
 wire \src_to_dst_data[6] ;
 wire \src_to_dst_data[7] ;
 wire \src_to_dst_data[8] ;
 wire \src_to_dst_data[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;

 XOR2_X1 _471_ (.A(src_req_prev),
    .B(src_req_sync),
    .Z(_146_));
 AND2_X1 _472_ (.A1(src_data_valid_sync),
    .A2(_146_),
    .ZN(_147_));
 NAND2_X1 _473_ (.A1(\dst_state[0] ),
    .A2(_147_),
    .ZN(_148_));
 NAND2_X1 _474_ (.A1(net169),
    .A2(net69),
    .ZN(_149_));
 NAND2_X1 _475_ (.A1(\dst_state[2] ),
    .A2(_149_),
    .ZN(_150_));
 NAND2_X1 _476_ (.A1(_148_),
    .A2(_150_),
    .ZN(_004_));
 BUF_X2 _477_ (.A(\src_state[0] ),
    .Z(_151_));
 NOR2_X2 _478_ (.A1(net65),
    .A2(net32),
    .ZN(_152_));
 BUF_X2 _479_ (.A(_009_),
    .Z(_153_));
 XNOR2_X2 _480_ (.A(dst_ack_prev),
    .B(dst_ack_sync),
    .ZN(_154_));
 NOR2_X1 _481_ (.A1(_153_),
    .A2(_154_),
    .ZN(_155_));
 BUF_X2 _482_ (.A(\src_state[1] ),
    .Z(_156_));
 AOI221_X2 _483_ (.A(\src_state[3] ),
    .B1(_151_),
    .B2(_152_),
    .C1(_155_),
    .C2(_156_),
    .ZN(_157_));
 INV_X1 _484_ (.A(_157_),
    .ZN(_006_));
 BUF_X8 _485_ (.A(\src_state[2] ),
    .Z(_158_));
 XOR2_X2 _486_ (.A(dst_ack_prev),
    .B(dst_ack_sync),
    .Z(_159_));
 BUF_X1 _487_ (.A(dst_data_valid_sync),
    .Z(_160_));
 OAI22_X1 _488_ (.A1(_160_),
    .A2(src_is_write_op_flag),
    .B1(_159_),
    .B2(_153_),
    .ZN(_161_));
 AOI22_X1 _489_ (.A1(_158_),
    .A2(_159_),
    .B1(_161_),
    .B2(_156_),
    .ZN(_162_));
 INV_X1 _490_ (.A(_162_),
    .ZN(_007_));
 INV_X1 _491_ (.A(\dst_state[0] ),
    .ZN(_163_));
 BUF_X2 _492_ (.A(dst_is_write_op),
    .Z(_164_));
 MUX2_X1 _493_ (.A(src_data_valid_sync),
    .B(_149_),
    .S(_164_),
    .Z(_165_));
 INV_X1 _494_ (.A(\dst_state[3] ),
    .ZN(_166_));
 OAI22_X1 _495_ (.A1(_163_),
    .A2(_147_),
    .B1(_165_),
    .B2(_166_),
    .ZN(_002_));
 BUF_X2 _496_ (.A(\dst_state[1] ),
    .Z(_167_));
 BUF_X1 _497_ (.A(router_out_valid),
    .Z(_168_));
 NOR2_X1 _498_ (.A1(_164_),
    .A2(_168_),
    .ZN(_169_));
 AOI21_X1 _499_ (.A(_011_),
    .B1(_146_),
    .B2(src_data_valid_sync),
    .ZN(_170_));
 OAI21_X1 _500_ (.A(_167_),
    .B1(_169_),
    .B2(_170_),
    .ZN(_171_));
 INV_X1 _501_ (.A(\dst_state[2] ),
    .ZN(_172_));
 OAI21_X1 _502_ (.A(_171_),
    .B1(_149_),
    .B2(_172_),
    .ZN(_003_));
 NAND3_X1 _503_ (.A1(_167_),
    .A2(_164_),
    .A3(_147_),
    .ZN(_173_));
 INV_X1 _504_ (.A(_164_),
    .ZN(_174_));
 NAND2_X1 _505_ (.A1(_167_),
    .A2(_174_),
    .ZN(_175_));
 INV_X1 _506_ (.A(_168_),
    .ZN(_176_));
 INV_X1 _507_ (.A(_011_),
    .ZN(_177_));
 AOI22_X1 _508_ (.A1(src_data_valid_sync),
    .A2(_174_),
    .B1(_177_),
    .B2(_149_),
    .ZN(_178_));
 OAI221_X1 _509_ (.A(_173_),
    .B1(_175_),
    .B2(_176_),
    .C1(_178_),
    .C2(_166_),
    .ZN(_005_));
 NAND2_X2 _510_ (.A1(_158_),
    .A2(_154_),
    .ZN(_179_));
 INV_X1 _511_ (.A(_151_),
    .ZN(_180_));
 OAI21_X1 _512_ (.A(_179_),
    .B1(_152_),
    .B2(_180_),
    .ZN(_008_));
 OR2_X1 _513_ (.A1(\dst_state[3] ),
    .A2(_167_),
    .ZN(net170));
 AOI21_X1 _514_ (.A(\dst_state[3] ),
    .B1(_167_),
    .B2(_168_),
    .ZN(_181_));
 NOR2_X1 _515_ (.A1(_164_),
    .A2(_181_),
    .ZN(_469_));
 NAND2_X1 _516_ (.A1(\dst_state[3] ),
    .A2(_164_),
    .ZN(_182_));
 NAND4_X1 _517_ (.A1(_148_),
    .A2(_150_),
    .A3(_173_),
    .A4(_182_),
    .ZN(_470_));
 AOI21_X1 _518_ (.A(_158_),
    .B1(_154_),
    .B2(_156_),
    .ZN(_183_));
 OAI221_X1 _519_ (.A(_179_),
    .B1(_183_),
    .B2(_153_),
    .C1(_010_),
    .C2(_152_),
    .ZN(_468_));
 INV_X1 _520_ (.A(_156_),
    .ZN(_184_));
 INV_X1 _521_ (.A(_160_),
    .ZN(_185_));
 NOR3_X1 _522_ (.A1(_184_),
    .A2(_185_),
    .A3(src_is_write_op_flag),
    .ZN(_001_));
 MUX2_X1 _523_ (.A(\dst_state[0] ),
    .B(_164_),
    .S(_167_),
    .Z(_186_));
 NAND2_X4 _524_ (.A1(_147_),
    .A2(_186_),
    .ZN(_187_));
 BUF_X4 _525_ (.A(_187_),
    .Z(_188_));
 MUX2_X1 _526_ (.A(_012_),
    .B(dst_ack),
    .S(_188_),
    .Z(_013_));
 MUX2_X1 _527_ (.A(\src_to_dst_data[0] ),
    .B(net137),
    .S(_188_),
    .Z(_014_));
 MUX2_X1 _528_ (.A(\src_to_dst_data[10] ),
    .B(net138),
    .S(_188_),
    .Z(_015_));
 MUX2_X1 _529_ (.A(\src_to_dst_data[11] ),
    .B(net139),
    .S(_188_),
    .Z(_016_));
 MUX2_X1 _530_ (.A(\src_to_dst_data[12] ),
    .B(net140),
    .S(_188_),
    .Z(_017_));
 MUX2_X1 _531_ (.A(\src_to_dst_data[13] ),
    .B(net141),
    .S(_188_),
    .Z(_018_));
 MUX2_X1 _532_ (.A(\src_to_dst_data[14] ),
    .B(net142),
    .S(_188_),
    .Z(_019_));
 MUX2_X1 _533_ (.A(\src_to_dst_data[15] ),
    .B(net143),
    .S(_188_),
    .Z(_020_));
 MUX2_X1 _534_ (.A(\src_to_dst_data[16] ),
    .B(net144),
    .S(_188_),
    .Z(_021_));
 MUX2_X1 _535_ (.A(\src_to_dst_data[17] ),
    .B(net145),
    .S(_188_),
    .Z(_022_));
 BUF_X4 _536_ (.A(_187_),
    .Z(_189_));
 MUX2_X1 _537_ (.A(\src_to_dst_data[18] ),
    .B(net146),
    .S(_189_),
    .Z(_023_));
 MUX2_X1 _538_ (.A(\src_to_dst_data[19] ),
    .B(net147),
    .S(_189_),
    .Z(_024_));
 MUX2_X1 _539_ (.A(\src_to_dst_data[1] ),
    .B(net148),
    .S(_189_),
    .Z(_025_));
 MUX2_X1 _540_ (.A(\src_to_dst_data[20] ),
    .B(net149),
    .S(_189_),
    .Z(_026_));
 MUX2_X1 _541_ (.A(\src_to_dst_data[21] ),
    .B(net150),
    .S(_189_),
    .Z(_027_));
 MUX2_X1 _542_ (.A(\src_to_dst_data[22] ),
    .B(net151),
    .S(_189_),
    .Z(_028_));
 MUX2_X1 _543_ (.A(\src_to_dst_data[23] ),
    .B(net152),
    .S(_189_),
    .Z(_029_));
 MUX2_X1 _544_ (.A(\src_to_dst_data[24] ),
    .B(net153),
    .S(_189_),
    .Z(_030_));
 MUX2_X1 _545_ (.A(\src_to_dst_data[25] ),
    .B(net154),
    .S(_189_),
    .Z(_031_));
 MUX2_X1 _546_ (.A(\src_to_dst_data[26] ),
    .B(net155),
    .S(_189_),
    .Z(_032_));
 BUF_X4 _547_ (.A(_187_),
    .Z(_190_));
 MUX2_X1 _548_ (.A(\src_to_dst_data[27] ),
    .B(net156),
    .S(_190_),
    .Z(_033_));
 MUX2_X1 _549_ (.A(\src_to_dst_data[28] ),
    .B(net157),
    .S(_190_),
    .Z(_034_));
 MUX2_X1 _550_ (.A(\src_to_dst_data[29] ),
    .B(net158),
    .S(_190_),
    .Z(_035_));
 MUX2_X1 _551_ (.A(\src_to_dst_data[2] ),
    .B(net159),
    .S(_190_),
    .Z(_036_));
 MUX2_X1 _552_ (.A(\src_to_dst_data[30] ),
    .B(net160),
    .S(_190_),
    .Z(_037_));
 MUX2_X1 _553_ (.A(\src_to_dst_data[31] ),
    .B(net161),
    .S(_190_),
    .Z(_038_));
 MUX2_X1 _554_ (.A(\src_to_dst_data[3] ),
    .B(net162),
    .S(_190_),
    .Z(_039_));
 MUX2_X1 _555_ (.A(\src_to_dst_data[4] ),
    .B(net163),
    .S(_190_),
    .Z(_040_));
 MUX2_X1 _556_ (.A(\src_to_dst_data[5] ),
    .B(net164),
    .S(_190_),
    .Z(_041_));
 MUX2_X1 _557_ (.A(\src_to_dst_data[6] ),
    .B(net165),
    .S(_190_),
    .Z(_042_));
 MUX2_X1 _558_ (.A(\src_to_dst_data[7] ),
    .B(net166),
    .S(_187_),
    .Z(_043_));
 MUX2_X1 _559_ (.A(\src_to_dst_data[8] ),
    .B(net167),
    .S(_187_),
    .Z(_044_));
 MUX2_X1 _560_ (.A(\src_to_dst_data[9] ),
    .B(net168),
    .S(_187_),
    .Z(_045_));
 MUX2_X1 _561_ (.A(src_is_write_op_sync),
    .B(_164_),
    .S(_148_),
    .Z(_046_));
 NAND3_X2 _562_ (.A1(_167_),
    .A2(_011_),
    .A3(_168_),
    .ZN(_191_));
 CLKBUF_X3 _563_ (.A(_191_),
    .Z(_192_));
 MUX2_X1 _564_ (.A(net70),
    .B(\dst_to_src_data[0] ),
    .S(_192_),
    .Z(_047_));
 MUX2_X1 _565_ (.A(net71),
    .B(\dst_to_src_data[10] ),
    .S(_192_),
    .Z(_048_));
 MUX2_X1 _566_ (.A(net72),
    .B(\dst_to_src_data[11] ),
    .S(_192_),
    .Z(_049_));
 MUX2_X1 _567_ (.A(net73),
    .B(\dst_to_src_data[12] ),
    .S(_192_),
    .Z(_050_));
 MUX2_X1 _568_ (.A(net74),
    .B(\dst_to_src_data[13] ),
    .S(_192_),
    .Z(_051_));
 MUX2_X1 _569_ (.A(net75),
    .B(\dst_to_src_data[14] ),
    .S(_192_),
    .Z(_052_));
 MUX2_X1 _570_ (.A(net76),
    .B(\dst_to_src_data[15] ),
    .S(_192_),
    .Z(_053_));
 MUX2_X1 _571_ (.A(net77),
    .B(\dst_to_src_data[16] ),
    .S(_192_),
    .Z(_054_));
 MUX2_X1 _572_ (.A(net78),
    .B(\dst_to_src_data[17] ),
    .S(_192_),
    .Z(_055_));
 MUX2_X1 _573_ (.A(net79),
    .B(\dst_to_src_data[18] ),
    .S(_192_),
    .Z(_056_));
 CLKBUF_X3 _574_ (.A(_191_),
    .Z(_193_));
 MUX2_X1 _575_ (.A(net80),
    .B(\dst_to_src_data[19] ),
    .S(_193_),
    .Z(_057_));
 MUX2_X1 _576_ (.A(net81),
    .B(\dst_to_src_data[1] ),
    .S(_193_),
    .Z(_058_));
 MUX2_X1 _577_ (.A(net82),
    .B(\dst_to_src_data[20] ),
    .S(_193_),
    .Z(_059_));
 MUX2_X1 _578_ (.A(net83),
    .B(\dst_to_src_data[21] ),
    .S(_193_),
    .Z(_060_));
 MUX2_X1 _579_ (.A(net84),
    .B(\dst_to_src_data[22] ),
    .S(_193_),
    .Z(_061_));
 MUX2_X1 _580_ (.A(net85),
    .B(\dst_to_src_data[23] ),
    .S(_193_),
    .Z(_062_));
 MUX2_X1 _581_ (.A(net86),
    .B(\dst_to_src_data[24] ),
    .S(_193_),
    .Z(_063_));
 MUX2_X1 _582_ (.A(net87),
    .B(\dst_to_src_data[25] ),
    .S(_193_),
    .Z(_064_));
 MUX2_X1 _583_ (.A(net88),
    .B(\dst_to_src_data[26] ),
    .S(_193_),
    .Z(_065_));
 MUX2_X1 _584_ (.A(net89),
    .B(\dst_to_src_data[27] ),
    .S(_193_),
    .Z(_066_));
 CLKBUF_X3 _585_ (.A(_191_),
    .Z(_194_));
 MUX2_X1 _586_ (.A(net90),
    .B(\dst_to_src_data[28] ),
    .S(_194_),
    .Z(_067_));
 MUX2_X1 _587_ (.A(net91),
    .B(\dst_to_src_data[29] ),
    .S(_194_),
    .Z(_068_));
 MUX2_X1 _588_ (.A(net92),
    .B(\dst_to_src_data[2] ),
    .S(_194_),
    .Z(_069_));
 MUX2_X1 _589_ (.A(net93),
    .B(\dst_to_src_data[30] ),
    .S(_194_),
    .Z(_070_));
 MUX2_X1 _590_ (.A(net94),
    .B(\dst_to_src_data[31] ),
    .S(_194_),
    .Z(_071_));
 MUX2_X1 _591_ (.A(net95),
    .B(\dst_to_src_data[3] ),
    .S(_194_),
    .Z(_072_));
 MUX2_X1 _592_ (.A(net96),
    .B(\dst_to_src_data[4] ),
    .S(_194_),
    .Z(_073_));
 MUX2_X1 _593_ (.A(net97),
    .B(\dst_to_src_data[5] ),
    .S(_194_),
    .Z(_074_));
 MUX2_X1 _594_ (.A(net98),
    .B(\dst_to_src_data[6] ),
    .S(_194_),
    .Z(_075_));
 MUX2_X1 _595_ (.A(net99),
    .B(\dst_to_src_data[7] ),
    .S(_194_),
    .Z(_076_));
 MUX2_X1 _596_ (.A(net100),
    .B(\dst_to_src_data[8] ),
    .S(_191_),
    .Z(_077_));
 MUX2_X1 _597_ (.A(net101),
    .B(\dst_to_src_data[9] ),
    .S(_191_),
    .Z(_078_));
 NAND3_X2 _598_ (.A1(_156_),
    .A2(_160_),
    .A3(_153_),
    .ZN(_195_));
 CLKBUF_X3 _599_ (.A(_195_),
    .Z(_196_));
 MUX2_X1 _600_ (.A(\dst_to_src_data[0] ),
    .B(net104),
    .S(_196_),
    .Z(_079_));
 MUX2_X1 _601_ (.A(\dst_to_src_data[10] ),
    .B(net105),
    .S(_196_),
    .Z(_080_));
 MUX2_X1 _602_ (.A(\dst_to_src_data[11] ),
    .B(net106),
    .S(_196_),
    .Z(_081_));
 MUX2_X1 _603_ (.A(\dst_to_src_data[12] ),
    .B(net107),
    .S(_196_),
    .Z(_082_));
 MUX2_X1 _604_ (.A(\dst_to_src_data[13] ),
    .B(net108),
    .S(_196_),
    .Z(_083_));
 MUX2_X1 _605_ (.A(\dst_to_src_data[14] ),
    .B(net109),
    .S(_196_),
    .Z(_084_));
 MUX2_X1 _606_ (.A(\dst_to_src_data[15] ),
    .B(net110),
    .S(_196_),
    .Z(_085_));
 MUX2_X1 _607_ (.A(\dst_to_src_data[16] ),
    .B(net111),
    .S(_196_),
    .Z(_086_));
 MUX2_X1 _608_ (.A(\dst_to_src_data[17] ),
    .B(net112),
    .S(_196_),
    .Z(_087_));
 MUX2_X1 _609_ (.A(\dst_to_src_data[18] ),
    .B(net113),
    .S(_196_),
    .Z(_088_));
 CLKBUF_X3 _610_ (.A(_195_),
    .Z(_197_));
 MUX2_X1 _611_ (.A(\dst_to_src_data[19] ),
    .B(net114),
    .S(_197_),
    .Z(_089_));
 MUX2_X1 _612_ (.A(\dst_to_src_data[1] ),
    .B(net115),
    .S(_197_),
    .Z(_090_));
 MUX2_X1 _613_ (.A(\dst_to_src_data[20] ),
    .B(net116),
    .S(_197_),
    .Z(_091_));
 MUX2_X1 _614_ (.A(\dst_to_src_data[21] ),
    .B(net117),
    .S(_197_),
    .Z(_092_));
 MUX2_X1 _615_ (.A(\dst_to_src_data[22] ),
    .B(net118),
    .S(_197_),
    .Z(_093_));
 MUX2_X1 _616_ (.A(\dst_to_src_data[23] ),
    .B(net119),
    .S(_197_),
    .Z(_094_));
 MUX2_X1 _617_ (.A(\dst_to_src_data[24] ),
    .B(net120),
    .S(_197_),
    .Z(_095_));
 MUX2_X1 _618_ (.A(\dst_to_src_data[25] ),
    .B(net121),
    .S(_197_),
    .Z(_096_));
 MUX2_X1 _619_ (.A(\dst_to_src_data[26] ),
    .B(net122),
    .S(_197_),
    .Z(_097_));
 MUX2_X1 _620_ (.A(\dst_to_src_data[27] ),
    .B(net123),
    .S(_197_),
    .Z(_098_));
 CLKBUF_X3 _621_ (.A(_195_),
    .Z(_198_));
 MUX2_X1 _622_ (.A(\dst_to_src_data[28] ),
    .B(net124),
    .S(_198_),
    .Z(_099_));
 MUX2_X1 _623_ (.A(\dst_to_src_data[29] ),
    .B(net125),
    .S(_198_),
    .Z(_100_));
 MUX2_X1 _624_ (.A(\dst_to_src_data[2] ),
    .B(net126),
    .S(_198_),
    .Z(_101_));
 MUX2_X1 _625_ (.A(\dst_to_src_data[30] ),
    .B(net127),
    .S(_198_),
    .Z(_102_));
 MUX2_X1 _626_ (.A(\dst_to_src_data[31] ),
    .B(net128),
    .S(_198_),
    .Z(_103_));
 MUX2_X1 _627_ (.A(\dst_to_src_data[3] ),
    .B(net129),
    .S(_198_),
    .Z(_104_));
 MUX2_X1 _628_ (.A(\dst_to_src_data[4] ),
    .B(net130),
    .S(_198_),
    .Z(_105_));
 MUX2_X1 _629_ (.A(\dst_to_src_data[5] ),
    .B(net131),
    .S(_198_),
    .Z(_106_));
 MUX2_X1 _630_ (.A(\dst_to_src_data[6] ),
    .B(net132),
    .S(_198_),
    .Z(_107_));
 MUX2_X1 _631_ (.A(\dst_to_src_data[7] ),
    .B(net133),
    .S(_198_),
    .Z(_108_));
 MUX2_X1 _632_ (.A(\dst_to_src_data[8] ),
    .B(net134),
    .S(_195_),
    .Z(_109_));
 MUX2_X1 _633_ (.A(\dst_to_src_data[9] ),
    .B(net135),
    .S(_195_),
    .Z(_110_));
 INV_X1 _634_ (.A(net136),
    .ZN(_199_));
 OR2_X1 _635_ (.A1(\src_state[3] ),
    .A2(_151_),
    .ZN(_200_));
 MUX2_X1 _636_ (.A(_160_),
    .B(_159_),
    .S(src_is_write_op_flag),
    .Z(_201_));
 MUX2_X1 _637_ (.A(_199_),
    .B(_200_),
    .S(_201_),
    .Z(_202_));
 OAI22_X1 _638_ (.A1(_199_),
    .A2(_200_),
    .B1(_202_),
    .B2(_184_),
    .ZN(_111_));
 INV_X1 _639_ (.A(net32),
    .ZN(_203_));
 OAI21_X1 _640_ (.A(src_is_write_op_flag),
    .B1(_203_),
    .B2(_010_),
    .ZN(_204_));
 INV_X1 _641_ (.A(net65),
    .ZN(_205_));
 OAI21_X1 _642_ (.A(_204_),
    .B1(_010_),
    .B2(_205_),
    .ZN(_112_));
 NAND2_X1 _643_ (.A1(_151_),
    .A2(_152_),
    .ZN(_206_));
 NOR2_X1 _644_ (.A1(_151_),
    .A2(_158_),
    .ZN(_207_));
 AOI21_X2 _645_ (.A(_207_),
    .B1(_158_),
    .B2(_153_),
    .ZN(_208_));
 NAND3_X4 _646_ (.A1(_206_),
    .A2(_179_),
    .A3(_208_),
    .ZN(_209_));
 BUF_X8 _647_ (.A(_209_),
    .Z(_210_));
 MUX2_X1 _648_ (.A(_000_),
    .B(src_req),
    .S(_210_),
    .Z(_113_));
 OR3_X2 _649_ (.A1(_180_),
    .A2(_158_),
    .A3(_152_),
    .ZN(_211_));
 CLKBUF_X3 _650_ (.A(_211_),
    .Z(_212_));
 NOR2_X1 _651_ (.A1(net11),
    .A2(_212_),
    .ZN(_213_));
 AND3_X2 _652_ (.A1(_158_),
    .A2(_155_),
    .A3(_206_),
    .ZN(_214_));
 INV_X1 _653_ (.A(net33),
    .ZN(_215_));
 INV_X1 _654_ (.A(\src_to_dst_data[0] ),
    .ZN(_216_));
 AOI221_X1 _655_ (.A(_213_),
    .B1(_214_),
    .B2(_215_),
    .C1(_216_),
    .C2(_210_),
    .ZN(_114_));
 NOR2_X1 _656_ (.A1(net12),
    .A2(_212_),
    .ZN(_217_));
 INV_X1 _657_ (.A(\src_to_dst_data[10] ),
    .ZN(_218_));
 INV_X1 _658_ (.A(net34),
    .ZN(_219_));
 BUF_X4 _659_ (.A(_214_),
    .Z(_220_));
 AOI221_X1 _660_ (.A(_217_),
    .B1(_210_),
    .B2(_218_),
    .C1(_219_),
    .C2(_220_),
    .ZN(_115_));
 NOR2_X1 _661_ (.A1(net13),
    .A2(_212_),
    .ZN(_221_));
 INV_X1 _662_ (.A(\src_to_dst_data[11] ),
    .ZN(_222_));
 INV_X1 _663_ (.A(net35),
    .ZN(_223_));
 AOI221_X1 _664_ (.A(_221_),
    .B1(_210_),
    .B2(_222_),
    .C1(_223_),
    .C2(_220_),
    .ZN(_116_));
 NOR2_X1 _665_ (.A1(net14),
    .A2(_212_),
    .ZN(_224_));
 INV_X1 _666_ (.A(\src_to_dst_data[12] ),
    .ZN(_225_));
 INV_X1 _667_ (.A(net36),
    .ZN(_226_));
 AOI221_X1 _668_ (.A(_224_),
    .B1(_210_),
    .B2(_225_),
    .C1(_226_),
    .C2(_220_),
    .ZN(_117_));
 NOR2_X1 _669_ (.A1(net15),
    .A2(_212_),
    .ZN(_227_));
 INV_X1 _670_ (.A(\src_to_dst_data[13] ),
    .ZN(_228_));
 INV_X1 _671_ (.A(net37),
    .ZN(_229_));
 AOI221_X1 _672_ (.A(_227_),
    .B1(_210_),
    .B2(_228_),
    .C1(_229_),
    .C2(_220_),
    .ZN(_118_));
 NOR2_X1 _673_ (.A1(net16),
    .A2(_212_),
    .ZN(_230_));
 INV_X1 _674_ (.A(\src_to_dst_data[14] ),
    .ZN(_231_));
 INV_X1 _675_ (.A(net38),
    .ZN(_232_));
 AOI221_X1 _676_ (.A(_230_),
    .B1(_210_),
    .B2(_231_),
    .C1(_232_),
    .C2(_220_),
    .ZN(_119_));
 NOR2_X1 _677_ (.A1(net17),
    .A2(_212_),
    .ZN(_233_));
 INV_X1 _678_ (.A(\src_to_dst_data[15] ),
    .ZN(_234_));
 INV_X1 _679_ (.A(net39),
    .ZN(_235_));
 AOI221_X1 _680_ (.A(_233_),
    .B1(_210_),
    .B2(_234_),
    .C1(_235_),
    .C2(_220_),
    .ZN(_120_));
 NOR2_X1 _681_ (.A1(net18),
    .A2(_212_),
    .ZN(_236_));
 INV_X1 _682_ (.A(\src_to_dst_data[16] ),
    .ZN(_237_));
 INV_X1 _683_ (.A(net40),
    .ZN(_238_));
 AOI221_X1 _684_ (.A(_236_),
    .B1(_210_),
    .B2(_237_),
    .C1(_238_),
    .C2(_220_),
    .ZN(_121_));
 NOR2_X1 _685_ (.A1(net19),
    .A2(_212_),
    .ZN(_239_));
 BUF_X8 _686_ (.A(_209_),
    .Z(_240_));
 INV_X1 _687_ (.A(\src_to_dst_data[17] ),
    .ZN(_241_));
 INV_X1 _688_ (.A(net41),
    .ZN(_242_));
 AOI221_X1 _689_ (.A(_239_),
    .B1(_240_),
    .B2(_241_),
    .C1(_242_),
    .C2(_220_),
    .ZN(_122_));
 NOR2_X1 _690_ (.A1(net20),
    .A2(_212_),
    .ZN(_243_));
 INV_X1 _691_ (.A(\src_to_dst_data[18] ),
    .ZN(_244_));
 INV_X1 _692_ (.A(net42),
    .ZN(_245_));
 AOI221_X1 _693_ (.A(_243_),
    .B1(_240_),
    .B2(_244_),
    .C1(_245_),
    .C2(_220_),
    .ZN(_123_));
 CLKBUF_X3 _694_ (.A(_211_),
    .Z(_246_));
 NOR2_X1 _695_ (.A1(net21),
    .A2(_246_),
    .ZN(_247_));
 INV_X1 _696_ (.A(\src_to_dst_data[19] ),
    .ZN(_248_));
 INV_X1 _697_ (.A(net43),
    .ZN(_249_));
 AOI221_X1 _698_ (.A(_247_),
    .B1(_240_),
    .B2(_248_),
    .C1(_249_),
    .C2(_220_),
    .ZN(_124_));
 NOR2_X1 _699_ (.A1(net22),
    .A2(_246_),
    .ZN(_250_));
 INV_X1 _700_ (.A(\src_to_dst_data[1] ),
    .ZN(_251_));
 INV_X1 _701_ (.A(net44),
    .ZN(_252_));
 BUF_X4 _702_ (.A(_214_),
    .Z(_253_));
 AOI221_X1 _703_ (.A(_250_),
    .B1(_240_),
    .B2(_251_),
    .C1(_252_),
    .C2(_253_),
    .ZN(_125_));
 NOR3_X1 _704_ (.A1(net65),
    .A2(_158_),
    .A3(net23),
    .ZN(_254_));
 INV_X1 _705_ (.A(net45),
    .ZN(_255_));
 AOI21_X1 _706_ (.A(_254_),
    .B1(_255_),
    .B2(_158_),
    .ZN(_256_));
 MUX2_X1 _707_ (.A(_256_),
    .B(\src_to_dst_data[20] ),
    .S(_210_),
    .Z(_126_));
 NOR2_X1 _708_ (.A1(net66),
    .A2(_246_),
    .ZN(_257_));
 INV_X1 _709_ (.A(\src_to_dst_data[21] ),
    .ZN(_258_));
 INV_X1 _710_ (.A(net46),
    .ZN(_259_));
 AOI221_X1 _711_ (.A(_257_),
    .B1(_240_),
    .B2(_258_),
    .C1(_259_),
    .C2(_253_),
    .ZN(_127_));
 NOR2_X1 _712_ (.A1(net67),
    .A2(_246_),
    .ZN(_260_));
 INV_X1 _713_ (.A(\src_to_dst_data[22] ),
    .ZN(_261_));
 INV_X1 _714_ (.A(net47),
    .ZN(_262_));
 AOI221_X1 _715_ (.A(_260_),
    .B1(_240_),
    .B2(_261_),
    .C1(_262_),
    .C2(_253_),
    .ZN(_128_));
 NOR2_X1 _716_ (.A1(net68),
    .A2(_246_),
    .ZN(_263_));
 INV_X1 _717_ (.A(\src_to_dst_data[23] ),
    .ZN(_264_));
 INV_X1 _718_ (.A(net48),
    .ZN(_265_));
 AOI221_X1 _719_ (.A(_263_),
    .B1(_240_),
    .B2(_264_),
    .C1(_265_),
    .C2(_253_),
    .ZN(_129_));
 NOR2_X1 _720_ (.A1(net1),
    .A2(_246_),
    .ZN(_266_));
 INV_X1 _721_ (.A(\src_to_dst_data[24] ),
    .ZN(_267_));
 INV_X1 _722_ (.A(net49),
    .ZN(_268_));
 AOI221_X1 _723_ (.A(_266_),
    .B1(_240_),
    .B2(_267_),
    .C1(_268_),
    .C2(_253_),
    .ZN(_130_));
 NOR2_X1 _724_ (.A1(net2),
    .A2(_246_),
    .ZN(_269_));
 INV_X1 _725_ (.A(\src_to_dst_data[25] ),
    .ZN(_270_));
 INV_X1 _726_ (.A(net50),
    .ZN(_271_));
 AOI221_X1 _727_ (.A(_269_),
    .B1(_240_),
    .B2(_270_),
    .C1(_271_),
    .C2(_253_),
    .ZN(_131_));
 NOR2_X1 _728_ (.A1(net3),
    .A2(_246_),
    .ZN(_272_));
 INV_X1 _729_ (.A(\src_to_dst_data[26] ),
    .ZN(_273_));
 INV_X1 _730_ (.A(net51),
    .ZN(_274_));
 AOI221_X1 _731_ (.A(_272_),
    .B1(_240_),
    .B2(_273_),
    .C1(_274_),
    .C2(_253_),
    .ZN(_132_));
 NOR2_X1 _732_ (.A1(net4),
    .A2(_246_),
    .ZN(_275_));
 BUF_X8 _733_ (.A(_209_),
    .Z(_276_));
 INV_X1 _734_ (.A(\src_to_dst_data[27] ),
    .ZN(_277_));
 INV_X1 _735_ (.A(net52),
    .ZN(_278_));
 AOI221_X1 _736_ (.A(_275_),
    .B1(_276_),
    .B2(_277_),
    .C1(_278_),
    .C2(_253_),
    .ZN(_133_));
 NOR2_X1 _737_ (.A1(net5),
    .A2(_246_),
    .ZN(_279_));
 INV_X1 _738_ (.A(\src_to_dst_data[28] ),
    .ZN(_280_));
 INV_X1 _739_ (.A(net53),
    .ZN(_281_));
 AOI221_X1 _740_ (.A(_279_),
    .B1(_276_),
    .B2(_280_),
    .C1(_281_),
    .C2(_253_),
    .ZN(_134_));
 CLKBUF_X3 _741_ (.A(_211_),
    .Z(_282_));
 NOR2_X1 _742_ (.A1(net6),
    .A2(_282_),
    .ZN(_283_));
 INV_X1 _743_ (.A(\src_to_dst_data[29] ),
    .ZN(_284_));
 INV_X1 _744_ (.A(net54),
    .ZN(_285_));
 AOI221_X1 _745_ (.A(_283_),
    .B1(_276_),
    .B2(_284_),
    .C1(_285_),
    .C2(_253_),
    .ZN(_135_));
 NOR2_X1 _746_ (.A1(net24),
    .A2(_282_),
    .ZN(_286_));
 INV_X1 _747_ (.A(\src_to_dst_data[2] ),
    .ZN(_287_));
 INV_X1 _748_ (.A(net55),
    .ZN(_288_));
 BUF_X4 _749_ (.A(_214_),
    .Z(_289_));
 AOI221_X1 _750_ (.A(_286_),
    .B1(_276_),
    .B2(_287_),
    .C1(_288_),
    .C2(_289_),
    .ZN(_136_));
 NOR2_X1 _751_ (.A1(net7),
    .A2(_282_),
    .ZN(_290_));
 INV_X1 _752_ (.A(\src_to_dst_data[30] ),
    .ZN(_291_));
 INV_X1 _753_ (.A(net56),
    .ZN(_292_));
 AOI221_X1 _754_ (.A(_290_),
    .B1(_276_),
    .B2(_291_),
    .C1(_292_),
    .C2(_289_),
    .ZN(_137_));
 NOR2_X1 _755_ (.A1(net8),
    .A2(_282_),
    .ZN(_293_));
 INV_X1 _756_ (.A(\src_to_dst_data[31] ),
    .ZN(_294_));
 INV_X1 _757_ (.A(net57),
    .ZN(_295_));
 AOI221_X1 _758_ (.A(_293_),
    .B1(_276_),
    .B2(_294_),
    .C1(_295_),
    .C2(_289_),
    .ZN(_138_));
 NOR2_X1 _759_ (.A1(net25),
    .A2(_282_),
    .ZN(_296_));
 INV_X1 _760_ (.A(\src_to_dst_data[3] ),
    .ZN(_297_));
 INV_X1 _761_ (.A(net58),
    .ZN(_298_));
 AOI221_X1 _762_ (.A(_296_),
    .B1(_276_),
    .B2(_297_),
    .C1(_298_),
    .C2(_289_),
    .ZN(_139_));
 NOR2_X1 _763_ (.A1(net26),
    .A2(_282_),
    .ZN(_299_));
 INV_X1 _764_ (.A(\src_to_dst_data[4] ),
    .ZN(_300_));
 INV_X1 _765_ (.A(net59),
    .ZN(_301_));
 AOI221_X1 _766_ (.A(_299_),
    .B1(_276_),
    .B2(_300_),
    .C1(_301_),
    .C2(_289_),
    .ZN(_140_));
 NOR2_X1 _767_ (.A1(net27),
    .A2(_282_),
    .ZN(_302_));
 INV_X1 _768_ (.A(\src_to_dst_data[5] ),
    .ZN(_303_));
 INV_X1 _769_ (.A(net60),
    .ZN(_304_));
 AOI221_X1 _770_ (.A(_302_),
    .B1(_276_),
    .B2(_303_),
    .C1(_304_),
    .C2(_289_),
    .ZN(_141_));
 NOR2_X1 _771_ (.A1(net28),
    .A2(_282_),
    .ZN(_305_));
 INV_X1 _772_ (.A(\src_to_dst_data[6] ),
    .ZN(_306_));
 INV_X1 _773_ (.A(net61),
    .ZN(_307_));
 AOI221_X1 _774_ (.A(_305_),
    .B1(_276_),
    .B2(_306_),
    .C1(_307_),
    .C2(_289_),
    .ZN(_142_));
 NOR2_X1 _775_ (.A1(net29),
    .A2(_282_),
    .ZN(_308_));
 INV_X1 _776_ (.A(\src_to_dst_data[7] ),
    .ZN(_309_));
 INV_X1 _777_ (.A(net62),
    .ZN(_310_));
 AOI221_X1 _778_ (.A(_308_),
    .B1(_209_),
    .B2(_309_),
    .C1(_310_),
    .C2(_289_),
    .ZN(_143_));
 NOR2_X1 _779_ (.A1(net30),
    .A2(_282_),
    .ZN(_311_));
 INV_X1 _780_ (.A(\src_to_dst_data[8] ),
    .ZN(_312_));
 INV_X1 _781_ (.A(net63),
    .ZN(_313_));
 AOI221_X1 _782_ (.A(_311_),
    .B1(_209_),
    .B2(_312_),
    .C1(_313_),
    .C2(_289_),
    .ZN(_144_));
 NOR2_X1 _783_ (.A1(net31),
    .A2(_211_),
    .ZN(_314_));
 INV_X1 _784_ (.A(\src_to_dst_data[9] ),
    .ZN(_315_));
 INV_X1 _785_ (.A(net64),
    .ZN(_316_));
 AOI221_X1 _786_ (.A(_314_),
    .B1(_209_),
    .B2(_315_),
    .C1(_316_),
    .C2(_289_),
    .ZN(_145_));
 DFFR_X1 \dst_ack$_DFFE_PN0P_  (.D(_013_),
    .RN(net10),
    .CK(net9),
    .Q(dst_ack),
    .QN(_012_));
 DFFR_X1 \dst_ack_prev$_DFF_PN0_  (.D(dst_ack_sync),
    .RN(net103),
    .CK(net102),
    .Q(dst_ack_prev),
    .QN(_450_));
 DFFR_X1 \dst_ack_sync_reg[0]$_DFF_PN0_  (.D(dst_ack),
    .RN(net103),
    .CK(net102),
    .Q(\dst_ack_sync_reg[0] ),
    .QN(_451_));
 DFFR_X2 \dst_ack_sync_reg[1]$_DFF_PN0_  (.D(\dst_ack_sync_reg[0] ),
    .RN(net103),
    .CK(net102),
    .Q(dst_ack_sync),
    .QN(_449_));
 DFFR_X1 \dst_data_reg[0]$_DFFE_PN0P_  (.D(_014_),
    .RN(net10),
    .CK(net9),
    .Q(net137),
    .QN(_448_));
 DFFR_X1 \dst_data_reg[10]$_DFFE_PN0P_  (.D(_015_),
    .RN(net10),
    .CK(net9),
    .Q(net138),
    .QN(_447_));
 DFFR_X1 \dst_data_reg[11]$_DFFE_PN0P_  (.D(_016_),
    .RN(net10),
    .CK(net9),
    .Q(net139),
    .QN(_446_));
 DFFR_X1 \dst_data_reg[12]$_DFFE_PN0P_  (.D(_017_),
    .RN(net10),
    .CK(net9),
    .Q(net140),
    .QN(_445_));
 DFFR_X1 \dst_data_reg[13]$_DFFE_PN0P_  (.D(_018_),
    .RN(net10),
    .CK(net9),
    .Q(net141),
    .QN(_444_));
 DFFR_X1 \dst_data_reg[14]$_DFFE_PN0P_  (.D(_019_),
    .RN(net10),
    .CK(net9),
    .Q(net142),
    .QN(_443_));
 DFFR_X1 \dst_data_reg[15]$_DFFE_PN0P_  (.D(_020_),
    .RN(net10),
    .CK(net9),
    .Q(net143),
    .QN(_442_));
 DFFR_X1 \dst_data_reg[16]$_DFFE_PN0P_  (.D(_021_),
    .RN(net10),
    .CK(net9),
    .Q(net144),
    .QN(_441_));
 DFFR_X1 \dst_data_reg[17]$_DFFE_PN0P_  (.D(_022_),
    .RN(net10),
    .CK(net9),
    .Q(net145),
    .QN(_440_));
 DFFR_X1 \dst_data_reg[18]$_DFFE_PN0P_  (.D(_023_),
    .RN(net10),
    .CK(net9),
    .Q(net146),
    .QN(_439_));
 DFFR_X1 \dst_data_reg[19]$_DFFE_PN0P_  (.D(_024_),
    .RN(net10),
    .CK(net9),
    .Q(net147),
    .QN(_438_));
 DFFR_X1 \dst_data_reg[1]$_DFFE_PN0P_  (.D(_025_),
    .RN(net10),
    .CK(net9),
    .Q(net148),
    .QN(_437_));
 DFFR_X1 \dst_data_reg[20]$_DFFE_PN0P_  (.D(_026_),
    .RN(net10),
    .CK(net9),
    .Q(net149),
    .QN(_436_));
 DFFR_X1 \dst_data_reg[21]$_DFFE_PN0P_  (.D(_027_),
    .RN(net10),
    .CK(net9),
    .Q(net150),
    .QN(_435_));
 DFFR_X1 \dst_data_reg[22]$_DFFE_PN0P_  (.D(_028_),
    .RN(net10),
    .CK(net9),
    .Q(net151),
    .QN(_434_));
 DFFR_X1 \dst_data_reg[23]$_DFFE_PN0P_  (.D(_029_),
    .RN(net10),
    .CK(net9),
    .Q(net152),
    .QN(_433_));
 DFFR_X1 \dst_data_reg[24]$_DFFE_PN0P_  (.D(_030_),
    .RN(net10),
    .CK(net9),
    .Q(net153),
    .QN(_432_));
 DFFR_X1 \dst_data_reg[25]$_DFFE_PN0P_  (.D(_031_),
    .RN(net10),
    .CK(net9),
    .Q(net154),
    .QN(_431_));
 DFFR_X1 \dst_data_reg[26]$_DFFE_PN0P_  (.D(_032_),
    .RN(net10),
    .CK(net9),
    .Q(net155),
    .QN(_430_));
 DFFR_X1 \dst_data_reg[27]$_DFFE_PN0P_  (.D(_033_),
    .RN(net10),
    .CK(net9),
    .Q(net156),
    .QN(_429_));
 DFFR_X1 \dst_data_reg[28]$_DFFE_PN0P_  (.D(_034_),
    .RN(net10),
    .CK(net9),
    .Q(net157),
    .QN(_428_));
 DFFR_X1 \dst_data_reg[29]$_DFFE_PN0P_  (.D(_035_),
    .RN(net10),
    .CK(net9),
    .Q(net158),
    .QN(_427_));
 DFFR_X1 \dst_data_reg[2]$_DFFE_PN0P_  (.D(_036_),
    .RN(net10),
    .CK(net9),
    .Q(net159),
    .QN(_426_));
 DFFR_X1 \dst_data_reg[30]$_DFFE_PN0P_  (.D(_037_),
    .RN(net10),
    .CK(net9),
    .Q(net160),
    .QN(_425_));
 DFFR_X1 \dst_data_reg[31]$_DFFE_PN0P_  (.D(_038_),
    .RN(net10),
    .CK(net9),
    .Q(net161),
    .QN(_424_));
 DFFR_X1 \dst_data_reg[3]$_DFFE_PN0P_  (.D(_039_),
    .RN(net10),
    .CK(net9),
    .Q(net162),
    .QN(_423_));
 DFFR_X1 \dst_data_reg[4]$_DFFE_PN0P_  (.D(_040_),
    .RN(net10),
    .CK(net9),
    .Q(net163),
    .QN(_422_));
 DFFR_X1 \dst_data_reg[5]$_DFFE_PN0P_  (.D(_041_),
    .RN(net10),
    .CK(net9),
    .Q(net164),
    .QN(_421_));
 DFFR_X1 \dst_data_reg[6]$_DFFE_PN0P_  (.D(_042_),
    .RN(net10),
    .CK(net9),
    .Q(net165),
    .QN(_420_));
 DFFR_X1 \dst_data_reg[7]$_DFFE_PN0P_  (.D(_043_),
    .RN(net10),
    .CK(net9),
    .Q(net166),
    .QN(_419_));
 DFFR_X1 \dst_data_reg[8]$_DFFE_PN0P_  (.D(_044_),
    .RN(net10),
    .CK(net9),
    .Q(net167),
    .QN(_418_));
 DFFR_X1 \dst_data_reg[9]$_DFFE_PN0P_  (.D(_045_),
    .RN(net10),
    .CK(net9),
    .Q(net168),
    .QN(_452_));
 DFFR_X1 \dst_data_valid$_DFF_PN0_  (.D(_469_),
    .RN(net10),
    .CK(net9),
    .Q(dst_data_valid),
    .QN(_453_));
 DFFR_X1 \dst_data_valid_sync_reg[0]$_DFF_PN0_  (.D(dst_data_valid),
    .RN(net103),
    .CK(net102),
    .Q(\dst_data_valid_sync_reg[0] ),
    .QN(_454_));
 DFFR_X1 \dst_data_valid_sync_reg[1]$_DFF_PN0_  (.D(\dst_data_valid_sync_reg[0] ),
    .RN(net103),
    .CK(net102),
    .Q(dst_data_valid_sync),
    .QN(_417_));
 DFFR_X1 \dst_is_write_op$_DFFE_PN0P_  (.D(_046_),
    .RN(net10),
    .CK(net9),
    .Q(dst_is_write_op),
    .QN(_011_));
 DFFS_X1 \dst_state[0]$_DFF_PN1_  (.D(_002_),
    .SN(net10),
    .CK(net9),
    .Q(\dst_state[0] ),
    .QN(_455_));
 DFFR_X1 \dst_state[1]$_DFF_PN0_  (.D(_003_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_state[1] ),
    .QN(_456_));
 DFFR_X1 \dst_state[2]$_DFF_PN0_  (.D(_004_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_state[2] ),
    .QN(_457_));
 DFFR_X1 \dst_state[3]$_DFF_PN0_  (.D(_005_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_state[3] ),
    .QN(_416_));
 DFFR_X1 \dst_to_src_data[0]$_DFFE_PN0P_  (.D(_047_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[0] ),
    .QN(_415_));
 DFFR_X1 \dst_to_src_data[10]$_DFFE_PN0P_  (.D(_048_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[10] ),
    .QN(_414_));
 DFFR_X1 \dst_to_src_data[11]$_DFFE_PN0P_  (.D(_049_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[11] ),
    .QN(_413_));
 DFFR_X1 \dst_to_src_data[12]$_DFFE_PN0P_  (.D(_050_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[12] ),
    .QN(_412_));
 DFFR_X1 \dst_to_src_data[13]$_DFFE_PN0P_  (.D(_051_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[13] ),
    .QN(_411_));
 DFFR_X1 \dst_to_src_data[14]$_DFFE_PN0P_  (.D(_052_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[14] ),
    .QN(_410_));
 DFFR_X1 \dst_to_src_data[15]$_DFFE_PN0P_  (.D(_053_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[15] ),
    .QN(_409_));
 DFFR_X1 \dst_to_src_data[16]$_DFFE_PN0P_  (.D(_054_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[16] ),
    .QN(_408_));
 DFFR_X1 \dst_to_src_data[17]$_DFFE_PN0P_  (.D(_055_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[17] ),
    .QN(_407_));
 DFFR_X1 \dst_to_src_data[18]$_DFFE_PN0P_  (.D(_056_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[18] ),
    .QN(_406_));
 DFFR_X1 \dst_to_src_data[19]$_DFFE_PN0P_  (.D(_057_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[19] ),
    .QN(_405_));
 DFFR_X1 \dst_to_src_data[1]$_DFFE_PN0P_  (.D(_058_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[1] ),
    .QN(_404_));
 DFFR_X1 \dst_to_src_data[20]$_DFFE_PN0P_  (.D(_059_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[20] ),
    .QN(_403_));
 DFFR_X1 \dst_to_src_data[21]$_DFFE_PN0P_  (.D(_060_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[21] ),
    .QN(_402_));
 DFFR_X1 \dst_to_src_data[22]$_DFFE_PN0P_  (.D(_061_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[22] ),
    .QN(_401_));
 DFFR_X1 \dst_to_src_data[23]$_DFFE_PN0P_  (.D(_062_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[23] ),
    .QN(_400_));
 DFFR_X1 \dst_to_src_data[24]$_DFFE_PN0P_  (.D(_063_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[24] ),
    .QN(_399_));
 DFFR_X1 \dst_to_src_data[25]$_DFFE_PN0P_  (.D(_064_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[25] ),
    .QN(_398_));
 DFFR_X1 \dst_to_src_data[26]$_DFFE_PN0P_  (.D(_065_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[26] ),
    .QN(_397_));
 DFFR_X1 \dst_to_src_data[27]$_DFFE_PN0P_  (.D(_066_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[27] ),
    .QN(_396_));
 DFFR_X1 \dst_to_src_data[28]$_DFFE_PN0P_  (.D(_067_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[28] ),
    .QN(_395_));
 DFFR_X1 \dst_to_src_data[29]$_DFFE_PN0P_  (.D(_068_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[29] ),
    .QN(_394_));
 DFFR_X1 \dst_to_src_data[2]$_DFFE_PN0P_  (.D(_069_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[2] ),
    .QN(_393_));
 DFFR_X1 \dst_to_src_data[30]$_DFFE_PN0P_  (.D(_070_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[30] ),
    .QN(_392_));
 DFFR_X1 \dst_to_src_data[31]$_DFFE_PN0P_  (.D(_071_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[31] ),
    .QN(_391_));
 DFFR_X1 \dst_to_src_data[3]$_DFFE_PN0P_  (.D(_072_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[3] ),
    .QN(_390_));
 DFFR_X1 \dst_to_src_data[4]$_DFFE_PN0P_  (.D(_073_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[4] ),
    .QN(_389_));
 DFFR_X1 \dst_to_src_data[5]$_DFFE_PN0P_  (.D(_074_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[5] ),
    .QN(_388_));
 DFFR_X1 \dst_to_src_data[6]$_DFFE_PN0P_  (.D(_075_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[6] ),
    .QN(_387_));
 DFFR_X1 \dst_to_src_data[7]$_DFFE_PN0P_  (.D(_076_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[7] ),
    .QN(_386_));
 DFFR_X1 \dst_to_src_data[8]$_DFFE_PN0P_  (.D(_077_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[8] ),
    .QN(_385_));
 DFFR_X1 \dst_to_src_data[9]$_DFFE_PN0P_  (.D(_078_),
    .RN(net10),
    .CK(net9),
    .Q(\dst_to_src_data[9] ),
    .QN(_458_));
 DFFR_X1 \dst_valid$_DFF_PN0_  (.D(_470_),
    .RN(net10),
    .CK(net9),
    .Q(net169),
    .QN(_384_));
 DFFR_X1 \mem_rdata[0]$_DFFE_PN0P_  (.D(_079_),
    .RN(net103),
    .CK(net102),
    .Q(net104),
    .QN(_383_));
 DFFR_X1 \mem_rdata[10]$_DFFE_PN0P_  (.D(_080_),
    .RN(net103),
    .CK(net102),
    .Q(net105),
    .QN(_382_));
 DFFR_X1 \mem_rdata[11]$_DFFE_PN0P_  (.D(_081_),
    .RN(net103),
    .CK(net102),
    .Q(net106),
    .QN(_381_));
 DFFR_X1 \mem_rdata[12]$_DFFE_PN0P_  (.D(_082_),
    .RN(net103),
    .CK(net102),
    .Q(net107),
    .QN(_380_));
 DFFR_X1 \mem_rdata[13]$_DFFE_PN0P_  (.D(_083_),
    .RN(net103),
    .CK(net102),
    .Q(net108),
    .QN(_379_));
 DFFR_X1 \mem_rdata[14]$_DFFE_PN0P_  (.D(_084_),
    .RN(net103),
    .CK(net102),
    .Q(net109),
    .QN(_378_));
 DFFR_X1 \mem_rdata[15]$_DFFE_PN0P_  (.D(_085_),
    .RN(net103),
    .CK(net102),
    .Q(net110),
    .QN(_377_));
 DFFR_X1 \mem_rdata[16]$_DFFE_PN0P_  (.D(_086_),
    .RN(net103),
    .CK(net102),
    .Q(net111),
    .QN(_376_));
 DFFR_X1 \mem_rdata[17]$_DFFE_PN0P_  (.D(_087_),
    .RN(net103),
    .CK(net102),
    .Q(net112),
    .QN(_375_));
 DFFR_X1 \mem_rdata[18]$_DFFE_PN0P_  (.D(_088_),
    .RN(net103),
    .CK(net102),
    .Q(net113),
    .QN(_374_));
 DFFR_X1 \mem_rdata[19]$_DFFE_PN0P_  (.D(_089_),
    .RN(net103),
    .CK(net102),
    .Q(net114),
    .QN(_373_));
 DFFR_X1 \mem_rdata[1]$_DFFE_PN0P_  (.D(_090_),
    .RN(net103),
    .CK(net102),
    .Q(net115),
    .QN(_372_));
 DFFR_X1 \mem_rdata[20]$_DFFE_PN0P_  (.D(_091_),
    .RN(net103),
    .CK(net102),
    .Q(net116),
    .QN(_371_));
 DFFR_X1 \mem_rdata[21]$_DFFE_PN0P_  (.D(_092_),
    .RN(net103),
    .CK(net102),
    .Q(net117),
    .QN(_370_));
 DFFR_X1 \mem_rdata[22]$_DFFE_PN0P_  (.D(_093_),
    .RN(net103),
    .CK(net102),
    .Q(net118),
    .QN(_369_));
 DFFR_X1 \mem_rdata[23]$_DFFE_PN0P_  (.D(_094_),
    .RN(net103),
    .CK(net102),
    .Q(net119),
    .QN(_368_));
 DFFR_X1 \mem_rdata[24]$_DFFE_PN0P_  (.D(_095_),
    .RN(net103),
    .CK(net102),
    .Q(net120),
    .QN(_367_));
 DFFR_X1 \mem_rdata[25]$_DFFE_PN0P_  (.D(_096_),
    .RN(net103),
    .CK(net102),
    .Q(net121),
    .QN(_366_));
 DFFR_X1 \mem_rdata[26]$_DFFE_PN0P_  (.D(_097_),
    .RN(net103),
    .CK(net102),
    .Q(net122),
    .QN(_365_));
 DFFR_X1 \mem_rdata[27]$_DFFE_PN0P_  (.D(_098_),
    .RN(net103),
    .CK(net102),
    .Q(net123),
    .QN(_364_));
 DFFR_X1 \mem_rdata[28]$_DFFE_PN0P_  (.D(_099_),
    .RN(net103),
    .CK(net102),
    .Q(net124),
    .QN(_363_));
 DFFR_X1 \mem_rdata[29]$_DFFE_PN0P_  (.D(_100_),
    .RN(net103),
    .CK(net102),
    .Q(net125),
    .QN(_362_));
 DFFR_X1 \mem_rdata[2]$_DFFE_PN0P_  (.D(_101_),
    .RN(net103),
    .CK(net102),
    .Q(net126),
    .QN(_361_));
 DFFR_X1 \mem_rdata[30]$_DFFE_PN0P_  (.D(_102_),
    .RN(net103),
    .CK(net102),
    .Q(net127),
    .QN(_360_));
 DFFR_X1 \mem_rdata[31]$_DFFE_PN0P_  (.D(_103_),
    .RN(net103),
    .CK(net102),
    .Q(net128),
    .QN(_359_));
 DFFR_X1 \mem_rdata[3]$_DFFE_PN0P_  (.D(_104_),
    .RN(net103),
    .CK(net102),
    .Q(net129),
    .QN(_358_));
 DFFR_X1 \mem_rdata[4]$_DFFE_PN0P_  (.D(_105_),
    .RN(net103),
    .CK(net102),
    .Q(net130),
    .QN(_357_));
 DFFR_X1 \mem_rdata[5]$_DFFE_PN0P_  (.D(_106_),
    .RN(net103),
    .CK(net102),
    .Q(net131),
    .QN(_356_));
 DFFR_X1 \mem_rdata[6]$_DFFE_PN0P_  (.D(_107_),
    .RN(net103),
    .CK(net102),
    .Q(net132),
    .QN(_355_));
 DFFR_X1 \mem_rdata[7]$_DFFE_PN0P_  (.D(_108_),
    .RN(net103),
    .CK(net102),
    .Q(net133),
    .QN(_354_));
 DFFR_X1 \mem_rdata[8]$_DFFE_PN0P_  (.D(_109_),
    .RN(net103),
    .CK(net102),
    .Q(net134),
    .QN(_353_));
 DFFR_X1 \mem_rdata[9]$_DFFE_PN0P_  (.D(_110_),
    .RN(net103),
    .CK(net102),
    .Q(net135),
    .QN(_352_));
 DFFR_X1 \mem_ready$_DFFE_PN0P_  (.D(_111_),
    .RN(net103),
    .CK(net102),
    .Q(net136),
    .QN(_459_));
 DFFR_X1 \src_data_valid$_DFF_PN0_  (.D(_468_),
    .RN(net103),
    .CK(net102),
    .Q(src_data_valid),
    .QN(_460_));
 DFFR_X1 \src_data_valid_sync_reg[0]$_DFF_PN0_  (.D(src_data_valid),
    .RN(net10),
    .CK(net9),
    .Q(\src_data_valid_sync_reg[0] ),
    .QN(_461_));
 DFFR_X1 \src_data_valid_sync_reg[1]$_DFF_PN0_  (.D(\src_data_valid_sync_reg[0] ),
    .RN(net10),
    .CK(net9),
    .Q(src_data_valid_sync),
    .QN(_351_));
 DFFR_X2 \src_is_write_op$_DFFE_PN0P_  (.D(_112_),
    .RN(net103),
    .CK(net102),
    .Q(src_is_write_op_flag),
    .QN(_009_));
 DFFR_X1 \src_is_write_op_sync_reg[0]$_DFF_PN0_  (.D(src_is_write_op_flag),
    .RN(net10),
    .CK(net9),
    .Q(\src_is_write_op_sync_reg[0] ),
    .QN(_462_));
 DFFR_X1 \src_is_write_op_sync_reg[1]$_DFF_PN0_  (.D(\src_is_write_op_sync_reg[0] ),
    .RN(net10),
    .CK(net9),
    .Q(src_is_write_op_sync),
    .QN(_350_));
 DFFR_X1 \src_req$_DFFE_PN0P_  (.D(_113_),
    .RN(net103),
    .CK(net102),
    .Q(src_req),
    .QN(_000_));
 DFFR_X1 \src_req_prev$_DFF_PN0_  (.D(src_req_sync),
    .RN(net10),
    .CK(net9),
    .Q(src_req_prev),
    .QN(_463_));
 DFFR_X1 \src_req_sync_reg[0]$_DFF_PN0_  (.D(src_req),
    .RN(net10),
    .CK(net9),
    .Q(\src_req_sync_reg[0] ),
    .QN(_464_));
 DFFR_X1 \src_req_sync_reg[1]$_DFF_PN0_  (.D(\src_req_sync_reg[0] ),
    .RN(net10),
    .CK(net9),
    .Q(src_req_sync),
    .QN(_465_));
 DFFS_X1 \src_state[0]$_DFF_PN1_  (.D(_006_),
    .SN(net103),
    .CK(net102),
    .Q(\src_state[0] ),
    .QN(_010_));
 DFFR_X1 \src_state[1]$_DFF_PN0_  (.D(_007_),
    .RN(net103),
    .CK(net102),
    .Q(\src_state[1] ),
    .QN(_466_));
 DFFR_X1 \src_state[2]$_DFF_PN0_  (.D(_008_),
    .RN(net103),
    .CK(net102),
    .Q(\src_state[2] ),
    .QN(_467_));
 DFFR_X1 \src_state[3]$_DFF_PN0_  (.D(_001_),
    .RN(net103),
    .CK(net102),
    .Q(\src_state[3] ),
    .QN(_349_));
 DFFR_X1 \src_to_dst_data[0]$_DFFE_PN0P_  (.D(_114_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[0] ),
    .QN(_348_));
 DFFR_X1 \src_to_dst_data[10]$_DFFE_PN0P_  (.D(_115_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[10] ),
    .QN(_347_));
 DFFR_X1 \src_to_dst_data[11]$_DFFE_PN0P_  (.D(_116_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[11] ),
    .QN(_346_));
 DFFR_X1 \src_to_dst_data[12]$_DFFE_PN0P_  (.D(_117_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[12] ),
    .QN(_345_));
 DFFR_X1 \src_to_dst_data[13]$_DFFE_PN0P_  (.D(_118_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[13] ),
    .QN(_344_));
 DFFR_X1 \src_to_dst_data[14]$_DFFE_PN0P_  (.D(_119_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[14] ),
    .QN(_343_));
 DFFR_X1 \src_to_dst_data[15]$_DFFE_PN0P_  (.D(_120_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[15] ),
    .QN(_342_));
 DFFR_X1 \src_to_dst_data[16]$_DFFE_PN0P_  (.D(_121_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[16] ),
    .QN(_341_));
 DFFR_X1 \src_to_dst_data[17]$_DFFE_PN0P_  (.D(_122_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[17] ),
    .QN(_340_));
 DFFR_X1 \src_to_dst_data[18]$_DFFE_PN0P_  (.D(_123_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[18] ),
    .QN(_339_));
 DFFR_X1 \src_to_dst_data[19]$_DFFE_PN0P_  (.D(_124_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[19] ),
    .QN(_338_));
 DFFR_X1 \src_to_dst_data[1]$_DFFE_PN0P_  (.D(_125_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[1] ),
    .QN(_337_));
 DFFR_X1 \src_to_dst_data[20]$_DFFE_PN0P_  (.D(_126_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[20] ),
    .QN(_336_));
 DFFR_X1 \src_to_dst_data[21]$_DFFE_PN0P_  (.D(_127_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[21] ),
    .QN(_335_));
 DFFR_X1 \src_to_dst_data[22]$_DFFE_PN0P_  (.D(_128_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[22] ),
    .QN(_334_));
 DFFR_X1 \src_to_dst_data[23]$_DFFE_PN0P_  (.D(_129_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[23] ),
    .QN(_333_));
 DFFR_X1 \src_to_dst_data[24]$_DFFE_PN0P_  (.D(_130_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[24] ),
    .QN(_332_));
 DFFR_X1 \src_to_dst_data[25]$_DFFE_PN0P_  (.D(_131_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[25] ),
    .QN(_331_));
 DFFR_X1 \src_to_dst_data[26]$_DFFE_PN0P_  (.D(_132_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[26] ),
    .QN(_330_));
 DFFR_X1 \src_to_dst_data[27]$_DFFE_PN0P_  (.D(_133_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[27] ),
    .QN(_329_));
 DFFR_X1 \src_to_dst_data[28]$_DFFE_PN0P_  (.D(_134_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[28] ),
    .QN(_328_));
 DFFR_X1 \src_to_dst_data[29]$_DFFE_PN0P_  (.D(_135_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[29] ),
    .QN(_327_));
 DFFR_X1 \src_to_dst_data[2]$_DFFE_PN0P_  (.D(_136_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[2] ),
    .QN(_326_));
 DFFR_X1 \src_to_dst_data[30]$_DFFE_PN0P_  (.D(_137_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[30] ),
    .QN(_325_));
 DFFR_X1 \src_to_dst_data[31]$_DFFE_PN0P_  (.D(_138_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[31] ),
    .QN(_324_));
 DFFR_X1 \src_to_dst_data[3]$_DFFE_PN0P_  (.D(_139_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[3] ),
    .QN(_323_));
 DFFR_X1 \src_to_dst_data[4]$_DFFE_PN0P_  (.D(_140_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[4] ),
    .QN(_322_));
 DFFR_X1 \src_to_dst_data[5]$_DFFE_PN0P_  (.D(_141_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[5] ),
    .QN(_321_));
 DFFR_X1 \src_to_dst_data[6]$_DFFE_PN0P_  (.D(_142_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[6] ),
    .QN(_320_));
 DFFR_X1 \src_to_dst_data[7]$_DFFE_PN0P_  (.D(_143_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[7] ),
    .QN(_319_));
 DFFR_X1 \src_to_dst_data[8]$_DFFE_PN0P_  (.D(_144_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[8] ),
    .QN(_318_));
 DFFR_X1 \src_to_dst_data[9]$_DFFE_PN0P_  (.D(_145_),
    .RN(net103),
    .CK(net102),
    .Q(\src_to_dst_data[9] ),
    .QN(_317_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_69 ();
 BUF_X1 input1 (.A(dest_id[0]),
    .Z(net1));
 BUF_X1 input2 (.A(dest_id[1]),
    .Z(net2));
 BUF_X1 input3 (.A(dest_id[2]),
    .Z(net3));
 BUF_X1 input4 (.A(dest_id[3]),
    .Z(net4));
 BUF_X1 input5 (.A(dest_id[4]),
    .Z(net5));
 BUF_X1 input6 (.A(dest_id[5]),
    .Z(net6));
 BUF_X1 input7 (.A(dest_id[6]),
    .Z(net7));
 BUF_X1 input8 (.A(dest_id[7]),
    .Z(net8));
 BUF_X16 input9 (.A(dst_clk),
    .Z(net9));
 BUF_X16 input10 (.A(dst_rst_n),
    .Z(net10));
 BUF_X1 input11 (.A(mem_addr[0]),
    .Z(net11));
 BUF_X1 input12 (.A(mem_addr[10]),
    .Z(net12));
 BUF_X1 input13 (.A(mem_addr[11]),
    .Z(net13));
 BUF_X1 input14 (.A(mem_addr[12]),
    .Z(net14));
 BUF_X1 input15 (.A(mem_addr[13]),
    .Z(net15));
 BUF_X1 input16 (.A(mem_addr[14]),
    .Z(net16));
 BUF_X1 input17 (.A(mem_addr[15]),
    .Z(net17));
 BUF_X1 input18 (.A(mem_addr[16]),
    .Z(net18));
 BUF_X1 input19 (.A(mem_addr[17]),
    .Z(net19));
 BUF_X1 input20 (.A(mem_addr[18]),
    .Z(net20));
 BUF_X1 input21 (.A(mem_addr[19]),
    .Z(net21));
 BUF_X1 input22 (.A(mem_addr[1]),
    .Z(net22));
 BUF_X1 input23 (.A(mem_addr[20]),
    .Z(net23));
 BUF_X1 input24 (.A(mem_addr[2]),
    .Z(net24));
 BUF_X1 input25 (.A(mem_addr[3]),
    .Z(net25));
 BUF_X1 input26 (.A(mem_addr[4]),
    .Z(net26));
 BUF_X1 input27 (.A(mem_addr[5]),
    .Z(net27));
 BUF_X1 input28 (.A(mem_addr[6]),
    .Z(net28));
 BUF_X1 input29 (.A(mem_addr[7]),
    .Z(net29));
 BUF_X1 input30 (.A(mem_addr[8]),
    .Z(net30));
 BUF_X1 input31 (.A(mem_addr[9]),
    .Z(net31));
 BUF_X1 input32 (.A(mem_read),
    .Z(net32));
 BUF_X1 input33 (.A(mem_wdata[0]),
    .Z(net33));
 BUF_X1 input34 (.A(mem_wdata[10]),
    .Z(net34));
 BUF_X1 input35 (.A(mem_wdata[11]),
    .Z(net35));
 BUF_X1 input36 (.A(mem_wdata[12]),
    .Z(net36));
 BUF_X1 input37 (.A(mem_wdata[13]),
    .Z(net37));
 BUF_X1 input38 (.A(mem_wdata[14]),
    .Z(net38));
 BUF_X1 input39 (.A(mem_wdata[15]),
    .Z(net39));
 BUF_X1 input40 (.A(mem_wdata[16]),
    .Z(net40));
 BUF_X1 input41 (.A(mem_wdata[17]),
    .Z(net41));
 BUF_X1 input42 (.A(mem_wdata[18]),
    .Z(net42));
 BUF_X1 input43 (.A(mem_wdata[19]),
    .Z(net43));
 BUF_X1 input44 (.A(mem_wdata[1]),
    .Z(net44));
 BUF_X1 input45 (.A(mem_wdata[20]),
    .Z(net45));
 BUF_X1 input46 (.A(mem_wdata[21]),
    .Z(net46));
 BUF_X1 input47 (.A(mem_wdata[22]),
    .Z(net47));
 BUF_X1 input48 (.A(mem_wdata[23]),
    .Z(net48));
 BUF_X1 input49 (.A(mem_wdata[24]),
    .Z(net49));
 BUF_X1 input50 (.A(mem_wdata[25]),
    .Z(net50));
 BUF_X1 input51 (.A(mem_wdata[26]),
    .Z(net51));
 BUF_X1 input52 (.A(mem_wdata[27]),
    .Z(net52));
 BUF_X1 input53 (.A(mem_wdata[28]),
    .Z(net53));
 BUF_X1 input54 (.A(mem_wdata[29]),
    .Z(net54));
 BUF_X1 input55 (.A(mem_wdata[2]),
    .Z(net55));
 BUF_X1 input56 (.A(mem_wdata[30]),
    .Z(net56));
 BUF_X1 input57 (.A(mem_wdata[31]),
    .Z(net57));
 BUF_X1 input58 (.A(mem_wdata[3]),
    .Z(net58));
 BUF_X1 input59 (.A(mem_wdata[4]),
    .Z(net59));
 BUF_X1 input60 (.A(mem_wdata[5]),
    .Z(net60));
 BUF_X1 input61 (.A(mem_wdata[6]),
    .Z(net61));
 BUF_X1 input62 (.A(mem_wdata[7]),
    .Z(net62));
 BUF_X1 input63 (.A(mem_wdata[8]),
    .Z(net63));
 BUF_X1 input64 (.A(mem_wdata[9]),
    .Z(net64));
 BUF_X1 input65 (.A(mem_write),
    .Z(net65));
 BUF_X1 input66 (.A(msg_type[0]),
    .Z(net66));
 BUF_X1 input67 (.A(msg_type[1]),
    .Z(net67));
 BUF_X1 input68 (.A(msg_type[2]),
    .Z(net68));
 BUF_X1 input69 (.A(router_in_ready),
    .Z(net69));
 BUF_X1 input70 (.A(router_out_data[0]),
    .Z(net70));
 BUF_X1 input71 (.A(router_out_data[10]),
    .Z(net71));
 BUF_X1 input72 (.A(router_out_data[11]),
    .Z(net72));
 BUF_X1 input73 (.A(router_out_data[12]),
    .Z(net73));
 BUF_X1 input74 (.A(router_out_data[13]),
    .Z(net74));
 BUF_X1 input75 (.A(router_out_data[14]),
    .Z(net75));
 BUF_X1 input76 (.A(router_out_data[15]),
    .Z(net76));
 BUF_X1 input77 (.A(router_out_data[16]),
    .Z(net77));
 BUF_X1 input78 (.A(router_out_data[17]),
    .Z(net78));
 BUF_X1 input79 (.A(router_out_data[18]),
    .Z(net79));
 BUF_X1 input80 (.A(router_out_data[19]),
    .Z(net80));
 BUF_X1 input81 (.A(router_out_data[1]),
    .Z(net81));
 BUF_X1 input82 (.A(router_out_data[20]),
    .Z(net82));
 BUF_X1 input83 (.A(router_out_data[21]),
    .Z(net83));
 BUF_X1 input84 (.A(router_out_data[22]),
    .Z(net84));
 BUF_X1 input85 (.A(router_out_data[23]),
    .Z(net85));
 BUF_X1 input86 (.A(router_out_data[24]),
    .Z(net86));
 BUF_X1 input87 (.A(router_out_data[25]),
    .Z(net87));
 BUF_X1 input88 (.A(router_out_data[26]),
    .Z(net88));
 BUF_X1 input89 (.A(router_out_data[27]),
    .Z(net89));
 BUF_X1 input90 (.A(router_out_data[28]),
    .Z(net90));
 BUF_X1 input91 (.A(router_out_data[29]),
    .Z(net91));
 BUF_X1 input92 (.A(router_out_data[2]),
    .Z(net92));
 BUF_X1 input93 (.A(router_out_data[30]),
    .Z(net93));
 BUF_X1 input94 (.A(router_out_data[31]),
    .Z(net94));
 BUF_X1 input95 (.A(router_out_data[3]),
    .Z(net95));
 BUF_X1 input96 (.A(router_out_data[4]),
    .Z(net96));
 BUF_X1 input97 (.A(router_out_data[5]),
    .Z(net97));
 BUF_X1 input98 (.A(router_out_data[6]),
    .Z(net98));
 BUF_X1 input99 (.A(router_out_data[7]),
    .Z(net99));
 BUF_X1 input100 (.A(router_out_data[8]),
    .Z(net100));
 BUF_X1 input101 (.A(router_out_data[9]),
    .Z(net101));
 BUF_X16 input102 (.A(src_clk),
    .Z(net102));
 BUF_X16 input103 (.A(src_rst_n),
    .Z(net103));
 BUF_X1 output104 (.A(net104),
    .Z(mem_rdata[0]));
 BUF_X1 output105 (.A(net105),
    .Z(mem_rdata[10]));
 BUF_X1 output106 (.A(net106),
    .Z(mem_rdata[11]));
 BUF_X1 output107 (.A(net107),
    .Z(mem_rdata[12]));
 BUF_X1 output108 (.A(net108),
    .Z(mem_rdata[13]));
 BUF_X1 output109 (.A(net109),
    .Z(mem_rdata[14]));
 BUF_X1 output110 (.A(net110),
    .Z(mem_rdata[15]));
 BUF_X1 output111 (.A(net111),
    .Z(mem_rdata[16]));
 BUF_X1 output112 (.A(net112),
    .Z(mem_rdata[17]));
 BUF_X1 output113 (.A(net113),
    .Z(mem_rdata[18]));
 BUF_X1 output114 (.A(net114),
    .Z(mem_rdata[19]));
 BUF_X1 output115 (.A(net115),
    .Z(mem_rdata[1]));
 BUF_X1 output116 (.A(net116),
    .Z(mem_rdata[20]));
 BUF_X1 output117 (.A(net117),
    .Z(mem_rdata[21]));
 BUF_X1 output118 (.A(net118),
    .Z(mem_rdata[22]));
 BUF_X1 output119 (.A(net119),
    .Z(mem_rdata[23]));
 BUF_X1 output120 (.A(net120),
    .Z(mem_rdata[24]));
 BUF_X1 output121 (.A(net121),
    .Z(mem_rdata[25]));
 BUF_X1 output122 (.A(net122),
    .Z(mem_rdata[26]));
 BUF_X1 output123 (.A(net123),
    .Z(mem_rdata[27]));
 BUF_X1 output124 (.A(net124),
    .Z(mem_rdata[28]));
 BUF_X1 output125 (.A(net125),
    .Z(mem_rdata[29]));
 BUF_X1 output126 (.A(net126),
    .Z(mem_rdata[2]));
 BUF_X1 output127 (.A(net127),
    .Z(mem_rdata[30]));
 BUF_X1 output128 (.A(net128),
    .Z(mem_rdata[31]));
 BUF_X1 output129 (.A(net129),
    .Z(mem_rdata[3]));
 BUF_X1 output130 (.A(net130),
    .Z(mem_rdata[4]));
 BUF_X1 output131 (.A(net131),
    .Z(mem_rdata[5]));
 BUF_X1 output132 (.A(net132),
    .Z(mem_rdata[6]));
 BUF_X1 output133 (.A(net133),
    .Z(mem_rdata[7]));
 BUF_X1 output134 (.A(net134),
    .Z(mem_rdata[8]));
 BUF_X1 output135 (.A(net135),
    .Z(mem_rdata[9]));
 BUF_X1 output136 (.A(net136),
    .Z(mem_ready));
 BUF_X1 output137 (.A(net137),
    .Z(router_in_data[0]));
 BUF_X1 output138 (.A(net138),
    .Z(router_in_data[10]));
 BUF_X1 output139 (.A(net139),
    .Z(router_in_data[11]));
 BUF_X1 output140 (.A(net140),
    .Z(router_in_data[12]));
 BUF_X1 output141 (.A(net141),
    .Z(router_in_data[13]));
 BUF_X1 output142 (.A(net142),
    .Z(router_in_data[14]));
 BUF_X1 output143 (.A(net143),
    .Z(router_in_data[15]));
 BUF_X1 output144 (.A(net144),
    .Z(router_in_data[16]));
 BUF_X1 output145 (.A(net145),
    .Z(router_in_data[17]));
 BUF_X1 output146 (.A(net146),
    .Z(router_in_data[18]));
 BUF_X1 output147 (.A(net147),
    .Z(router_in_data[19]));
 BUF_X1 output148 (.A(net148),
    .Z(router_in_data[1]));
 BUF_X1 output149 (.A(net149),
    .Z(router_in_data[20]));
 BUF_X1 output150 (.A(net150),
    .Z(router_in_data[21]));
 BUF_X1 output151 (.A(net151),
    .Z(router_in_data[22]));
 BUF_X1 output152 (.A(net152),
    .Z(router_in_data[23]));
 BUF_X1 output153 (.A(net153),
    .Z(router_in_data[24]));
 BUF_X1 output154 (.A(net154),
    .Z(router_in_data[25]));
 BUF_X1 output155 (.A(net155),
    .Z(router_in_data[26]));
 BUF_X1 output156 (.A(net156),
    .Z(router_in_data[27]));
 BUF_X1 output157 (.A(net157),
    .Z(router_in_data[28]));
 BUF_X1 output158 (.A(net158),
    .Z(router_in_data[29]));
 BUF_X1 output159 (.A(net159),
    .Z(router_in_data[2]));
 BUF_X1 output160 (.A(net160),
    .Z(router_in_data[30]));
 BUF_X1 output161 (.A(net161),
    .Z(router_in_data[31]));
 BUF_X1 output162 (.A(net162),
    .Z(router_in_data[3]));
 BUF_X1 output163 (.A(net163),
    .Z(router_in_data[4]));
 BUF_X1 output164 (.A(net164),
    .Z(router_in_data[5]));
 BUF_X1 output165 (.A(net165),
    .Z(router_in_data[6]));
 BUF_X1 output166 (.A(net166),
    .Z(router_in_data[7]));
 BUF_X1 output167 (.A(net167),
    .Z(router_in_data[8]));
 BUF_X1 output168 (.A(net168),
    .Z(router_in_data[9]));
 BUF_X1 output169 (.A(net169),
    .Z(router_in_valid));
 BUF_X1 output170 (.A(net170),
    .Z(router_out_ready));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X4 FILLER_0_17 ();
 FILLCELL_X32 FILLER_0_80 ();
 FILLCELL_X16 FILLER_0_112 ();
 FILLCELL_X8 FILLER_0_128 ();
 FILLCELL_X1 FILLER_0_136 ();
 FILLCELL_X8 FILLER_0_166 ();
 FILLCELL_X2 FILLER_0_174 ();
 FILLCELL_X1 FILLER_0_176 ();
 FILLCELL_X1 FILLER_0_180 ();
 FILLCELL_X2 FILLER_0_191 ();
 FILLCELL_X2 FILLER_0_196 ();
 FILLCELL_X2 FILLER_0_211 ();
 FILLCELL_X2 FILLER_0_219 ();
 FILLCELL_X4 FILLER_0_238 ();
 FILLCELL_X1 FILLER_0_242 ();
 FILLCELL_X1 FILLER_0_263 ();
 FILLCELL_X4 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_5 ();
 FILLCELL_X2 FILLER_1_9 ();
 FILLCELL_X2 FILLER_1_43 ();
 FILLCELL_X1 FILLER_1_68 ();
 FILLCELL_X32 FILLER_1_89 ();
 FILLCELL_X8 FILLER_1_121 ();
 FILLCELL_X2 FILLER_1_129 ();
 FILLCELL_X1 FILLER_1_131 ();
 FILLCELL_X8 FILLER_1_158 ();
 FILLCELL_X4 FILLER_1_166 ();
 FILLCELL_X2 FILLER_1_190 ();
 FILLCELL_X1 FILLER_1_192 ();
 FILLCELL_X4 FILLER_1_200 ();
 FILLCELL_X1 FILLER_1_204 ();
 FILLCELL_X4 FILLER_1_245 ();
 FILLCELL_X8 FILLER_1_256 ();
 FILLCELL_X2 FILLER_2_1 ();
 FILLCELL_X4 FILLER_2_56 ();
 FILLCELL_X2 FILLER_2_60 ();
 FILLCELL_X2 FILLER_2_68 ();
 FILLCELL_X32 FILLER_2_72 ();
 FILLCELL_X32 FILLER_2_104 ();
 FILLCELL_X4 FILLER_2_136 ();
 FILLCELL_X2 FILLER_2_140 ();
 FILLCELL_X1 FILLER_2_142 ();
 FILLCELL_X8 FILLER_2_166 ();
 FILLCELL_X2 FILLER_2_241 ();
 FILLCELL_X1 FILLER_2_263 ();
 FILLCELL_X2 FILLER_3_1 ();
 FILLCELL_X1 FILLER_3_3 ();
 FILLCELL_X8 FILLER_3_27 ();
 FILLCELL_X4 FILLER_3_35 ();
 FILLCELL_X8 FILLER_3_50 ();
 FILLCELL_X32 FILLER_3_78 ();
 FILLCELL_X32 FILLER_3_110 ();
 FILLCELL_X4 FILLER_3_142 ();
 FILLCELL_X2 FILLER_3_149 ();
 FILLCELL_X4 FILLER_3_157 ();
 FILLCELL_X8 FILLER_3_165 ();
 FILLCELL_X4 FILLER_3_173 ();
 FILLCELL_X2 FILLER_3_177 ();
 FILLCELL_X4 FILLER_3_206 ();
 FILLCELL_X1 FILLER_3_210 ();
 FILLCELL_X8 FILLER_3_218 ();
 FILLCELL_X4 FILLER_3_226 ();
 FILLCELL_X2 FILLER_3_230 ();
 FILLCELL_X32 FILLER_4_27 ();
 FILLCELL_X32 FILLER_4_79 ();
 FILLCELL_X16 FILLER_4_111 ();
 FILLCELL_X8 FILLER_4_127 ();
 FILLCELL_X4 FILLER_4_135 ();
 FILLCELL_X2 FILLER_4_139 ();
 FILLCELL_X1 FILLER_4_141 ();
 FILLCELL_X16 FILLER_4_166 ();
 FILLCELL_X4 FILLER_4_182 ();
 FILLCELL_X16 FILLER_4_206 ();
 FILLCELL_X8 FILLER_4_222 ();
 FILLCELL_X4 FILLER_4_237 ();
 FILLCELL_X8 FILLER_4_248 ();
 FILLCELL_X2 FILLER_4_256 ();
 FILLCELL_X1 FILLER_5_4 ();
 FILLCELL_X1 FILLER_5_7 ();
 FILLCELL_X1 FILLER_5_17 ();
 FILLCELL_X1 FILLER_5_20 ();
 FILLCELL_X8 FILLER_5_48 ();
 FILLCELL_X4 FILLER_5_56 ();
 FILLCELL_X2 FILLER_5_60 ();
 FILLCELL_X8 FILLER_5_135 ();
 FILLCELL_X32 FILLER_5_178 ();
 FILLCELL_X8 FILLER_5_210 ();
 FILLCELL_X4 FILLER_5_238 ();
 FILLCELL_X1 FILLER_5_242 ();
 FILLCELL_X1 FILLER_5_263 ();
 FILLCELL_X2 FILLER_6_1 ();
 FILLCELL_X1 FILLER_6_3 ();
 FILLCELL_X8 FILLER_6_13 ();
 FILLCELL_X4 FILLER_6_21 ();
 FILLCELL_X2 FILLER_6_25 ();
 FILLCELL_X1 FILLER_6_27 ();
 FILLCELL_X32 FILLER_6_35 ();
 FILLCELL_X32 FILLER_6_67 ();
 FILLCELL_X16 FILLER_6_99 ();
 FILLCELL_X4 FILLER_6_115 ();
 FILLCELL_X1 FILLER_6_119 ();
 FILLCELL_X1 FILLER_6_151 ();
 FILLCELL_X1 FILLER_6_175 ();
 FILLCELL_X32 FILLER_6_178 ();
 FILLCELL_X4 FILLER_6_210 ();
 FILLCELL_X4 FILLER_6_234 ();
 FILLCELL_X1 FILLER_6_238 ();
 FILLCELL_X2 FILLER_6_262 ();
 FILLCELL_X2 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_51 ();
 FILLCELL_X16 FILLER_7_83 ();
 FILLCELL_X8 FILLER_7_99 ();
 FILLCELL_X2 FILLER_7_107 ();
 FILLCELL_X8 FILLER_7_129 ();
 FILLCELL_X4 FILLER_7_137 ();
 FILLCELL_X1 FILLER_7_141 ();
 FILLCELL_X32 FILLER_7_183 ();
 FILLCELL_X8 FILLER_7_215 ();
 FILLCELL_X4 FILLER_7_223 ();
 FILLCELL_X4 FILLER_7_234 ();
 FILLCELL_X2 FILLER_7_238 ();
 FILLCELL_X4 FILLER_7_247 ();
 FILLCELL_X1 FILLER_7_251 ();
 FILLCELL_X2 FILLER_7_255 ();
 FILLCELL_X1 FILLER_7_257 ();
 FILLCELL_X1 FILLER_8_7 ();
 FILLCELL_X8 FILLER_8_10 ();
 FILLCELL_X1 FILLER_8_18 ();
 FILLCELL_X8 FILLER_8_22 ();
 FILLCELL_X1 FILLER_8_30 ();
 FILLCELL_X8 FILLER_8_78 ();
 FILLCELL_X4 FILLER_8_86 ();
 FILLCELL_X8 FILLER_8_110 ();
 FILLCELL_X2 FILLER_8_118 ();
 FILLCELL_X1 FILLER_8_120 ();
 FILLCELL_X16 FILLER_8_172 ();
 FILLCELL_X4 FILLER_8_188 ();
 FILLCELL_X1 FILLER_8_192 ();
 FILLCELL_X32 FILLER_8_198 ();
 FILLCELL_X2 FILLER_8_230 ();
 FILLCELL_X2 FILLER_8_239 ();
 FILLCELL_X4 FILLER_8_248 ();
 FILLCELL_X1 FILLER_8_252 ();
 FILLCELL_X2 FILLER_8_256 ();
 FILLCELL_X1 FILLER_9_6 ();
 FILLCELL_X1 FILLER_9_13 ();
 FILLCELL_X1 FILLER_9_34 ();
 FILLCELL_X16 FILLER_9_62 ();
 FILLCELL_X2 FILLER_9_78 ();
 FILLCELL_X16 FILLER_9_122 ();
 FILLCELL_X8 FILLER_9_138 ();
 FILLCELL_X4 FILLER_9_146 ();
 FILLCELL_X2 FILLER_9_150 ();
 FILLCELL_X2 FILLER_9_155 ();
 FILLCELL_X1 FILLER_9_157 ();
 FILLCELL_X16 FILLER_9_162 ();
 FILLCELL_X8 FILLER_9_178 ();
 FILLCELL_X4 FILLER_9_186 ();
 FILLCELL_X2 FILLER_9_190 ();
 FILLCELL_X1 FILLER_9_192 ();
 FILLCELL_X8 FILLER_9_213 ();
 FILLCELL_X2 FILLER_9_241 ();
 FILLCELL_X1 FILLER_9_263 ();
 FILLCELL_X2 FILLER_10_4 ();
 FILLCELL_X1 FILLER_10_6 ();
 FILLCELL_X4 FILLER_10_20 ();
 FILLCELL_X1 FILLER_10_24 ();
 FILLCELL_X16 FILLER_10_32 ();
 FILLCELL_X8 FILLER_10_48 ();
 FILLCELL_X4 FILLER_10_56 ();
 FILLCELL_X2 FILLER_10_60 ();
 FILLCELL_X1 FILLER_10_62 ();
 FILLCELL_X16 FILLER_10_70 ();
 FILLCELL_X4 FILLER_10_86 ();
 FILLCELL_X16 FILLER_10_119 ();
 FILLCELL_X16 FILLER_10_175 ();
 FILLCELL_X8 FILLER_10_191 ();
 FILLCELL_X4 FILLER_10_199 ();
 FILLCELL_X1 FILLER_10_203 ();
 FILLCELL_X4 FILLER_10_218 ();
 FILLCELL_X1 FILLER_10_222 ();
 FILLCELL_X1 FILLER_10_263 ();
 FILLCELL_X1 FILLER_11_1 ();
 FILLCELL_X1 FILLER_11_27 ();
 FILLCELL_X32 FILLER_11_48 ();
 FILLCELL_X16 FILLER_11_80 ();
 FILLCELL_X1 FILLER_11_96 ();
 FILLCELL_X4 FILLER_11_107 ();
 FILLCELL_X1 FILLER_11_111 ();
 FILLCELL_X32 FILLER_11_134 ();
 FILLCELL_X1 FILLER_11_166 ();
 FILLCELL_X8 FILLER_11_187 ();
 FILLCELL_X4 FILLER_11_195 ();
 FILLCELL_X2 FILLER_11_199 ();
 FILLCELL_X1 FILLER_11_201 ();
 FILLCELL_X4 FILLER_11_227 ();
 FILLCELL_X1 FILLER_11_231 ();
 FILLCELL_X2 FILLER_11_239 ();
 FILLCELL_X4 FILLER_11_248 ();
 FILLCELL_X2 FILLER_11_258 ();
 FILLCELL_X1 FILLER_11_260 ();
 FILLCELL_X2 FILLER_12_1 ();
 FILLCELL_X2 FILLER_12_6 ();
 FILLCELL_X1 FILLER_12_8 ();
 FILLCELL_X4 FILLER_12_15 ();
 FILLCELL_X2 FILLER_12_19 ();
 FILLCELL_X1 FILLER_12_21 ();
 FILLCELL_X4 FILLER_12_25 ();
 FILLCELL_X2 FILLER_12_29 ();
 FILLCELL_X16 FILLER_12_34 ();
 FILLCELL_X2 FILLER_12_50 ();
 FILLCELL_X2 FILLER_12_79 ();
 FILLCELL_X8 FILLER_12_107 ();
 FILLCELL_X2 FILLER_12_115 ();
 FILLCELL_X32 FILLER_12_139 ();
 FILLCELL_X4 FILLER_12_171 ();
 FILLCELL_X2 FILLER_12_175 ();
 FILLCELL_X4 FILLER_12_197 ();
 FILLCELL_X2 FILLER_12_201 ();
 FILLCELL_X2 FILLER_12_230 ();
 FILLCELL_X1 FILLER_12_232 ();
 FILLCELL_X4 FILLER_12_236 ();
 FILLCELL_X1 FILLER_12_240 ();
 FILLCELL_X1 FILLER_12_248 ();
 FILLCELL_X2 FILLER_12_252 ();
 FILLCELL_X1 FILLER_12_254 ();
 FILLCELL_X4 FILLER_13_13 ();
 FILLCELL_X1 FILLER_13_17 ();
 FILLCELL_X2 FILLER_13_45 ();
 FILLCELL_X2 FILLER_13_74 ();
 FILLCELL_X4 FILLER_13_86 ();
 FILLCELL_X1 FILLER_13_100 ();
 FILLCELL_X32 FILLER_13_141 ();
 FILLCELL_X16 FILLER_13_173 ();
 FILLCELL_X2 FILLER_13_189 ();
 FILLCELL_X1 FILLER_13_191 ();
 FILLCELL_X2 FILLER_13_199 ();
 FILLCELL_X2 FILLER_14_26 ();
 FILLCELL_X8 FILLER_14_33 ();
 FILLCELL_X1 FILLER_14_41 ();
 FILLCELL_X8 FILLER_14_53 ();
 FILLCELL_X4 FILLER_14_85 ();
 FILLCELL_X1 FILLER_14_89 ();
 FILLCELL_X2 FILLER_14_92 ();
 FILLCELL_X1 FILLER_14_109 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X16 FILLER_14_193 ();
 FILLCELL_X1 FILLER_14_209 ();
 FILLCELL_X4 FILLER_14_217 ();
 FILLCELL_X2 FILLER_14_221 ();
 FILLCELL_X1 FILLER_14_263 ();
 FILLCELL_X1 FILLER_15_12 ();
 FILLCELL_X4 FILLER_15_18 ();
 FILLCELL_X2 FILLER_15_22 ();
 FILLCELL_X1 FILLER_15_24 ();
 FILLCELL_X1 FILLER_15_31 ();
 FILLCELL_X4 FILLER_15_36 ();
 FILLCELL_X2 FILLER_15_40 ();
 FILLCELL_X16 FILLER_15_62 ();
 FILLCELL_X8 FILLER_15_78 ();
 FILLCELL_X1 FILLER_15_86 ();
 FILLCELL_X8 FILLER_15_89 ();
 FILLCELL_X1 FILLER_15_97 ();
 FILLCELL_X4 FILLER_15_111 ();
 FILLCELL_X32 FILLER_15_135 ();
 FILLCELL_X16 FILLER_15_167 ();
 FILLCELL_X4 FILLER_15_190 ();
 FILLCELL_X1 FILLER_15_194 ();
 FILLCELL_X2 FILLER_15_222 ();
 FILLCELL_X1 FILLER_15_224 ();
 FILLCELL_X2 FILLER_15_228 ();
 FILLCELL_X1 FILLER_15_230 ();
 FILLCELL_X2 FILLER_15_255 ();
 FILLCELL_X1 FILLER_15_257 ();
 FILLCELL_X1 FILLER_16_15 ();
 FILLCELL_X8 FILLER_16_36 ();
 FILLCELL_X2 FILLER_16_44 ();
 FILLCELL_X4 FILLER_16_66 ();
 FILLCELL_X8 FILLER_16_75 ();
 FILLCELL_X4 FILLER_16_93 ();
 FILLCELL_X32 FILLER_16_116 ();
 FILLCELL_X16 FILLER_16_148 ();
 FILLCELL_X2 FILLER_16_164 ();
 FILLCELL_X2 FILLER_16_193 ();
 FILLCELL_X1 FILLER_16_195 ();
 FILLCELL_X16 FILLER_16_216 ();
 FILLCELL_X4 FILLER_16_232 ();
 FILLCELL_X1 FILLER_16_236 ();
 FILLCELL_X1 FILLER_16_260 ();
 FILLCELL_X2 FILLER_17_10 ();
 FILLCELL_X4 FILLER_17_15 ();
 FILLCELL_X2 FILLER_17_22 ();
 FILLCELL_X1 FILLER_17_24 ();
 FILLCELL_X2 FILLER_17_86 ();
 FILLCELL_X32 FILLER_17_121 ();
 FILLCELL_X32 FILLER_17_153 ();
 FILLCELL_X4 FILLER_17_185 ();
 FILLCELL_X1 FILLER_17_189 ();
 FILLCELL_X4 FILLER_17_210 ();
 FILLCELL_X2 FILLER_17_241 ();
 FILLCELL_X1 FILLER_17_263 ();
 FILLCELL_X4 FILLER_18_12 ();
 FILLCELL_X2 FILLER_18_16 ();
 FILLCELL_X4 FILLER_18_20 ();
 FILLCELL_X2 FILLER_18_24 ();
 FILLCELL_X1 FILLER_18_26 ();
 FILLCELL_X4 FILLER_18_34 ();
 FILLCELL_X2 FILLER_18_38 ();
 FILLCELL_X32 FILLER_18_53 ();
 FILLCELL_X32 FILLER_18_85 ();
 FILLCELL_X32 FILLER_18_117 ();
 FILLCELL_X32 FILLER_18_149 ();
 FILLCELL_X16 FILLER_18_181 ();
 FILLCELL_X4 FILLER_18_197 ();
 FILLCELL_X2 FILLER_18_201 ();
 FILLCELL_X8 FILLER_18_217 ();
 FILLCELL_X2 FILLER_18_259 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_5 ();
 FILLCELL_X1 FILLER_19_30 ();
 FILLCELL_X32 FILLER_19_51 ();
 FILLCELL_X32 FILLER_19_83 ();
 FILLCELL_X32 FILLER_19_115 ();
 FILLCELL_X32 FILLER_19_147 ();
 FILLCELL_X16 FILLER_19_179 ();
 FILLCELL_X8 FILLER_19_195 ();
 FILLCELL_X4 FILLER_19_203 ();
 FILLCELL_X2 FILLER_19_227 ();
 FILLCELL_X1 FILLER_19_229 ();
 FILLCELL_X8 FILLER_19_233 ();
 FILLCELL_X1 FILLER_19_241 ();
 FILLCELL_X2 FILLER_19_252 ();
 FILLCELL_X1 FILLER_19_254 ();
 FILLCELL_X2 FILLER_19_258 ();
 FILLCELL_X1 FILLER_19_260 ();
 FILLCELL_X8 FILLER_20_4 ();
 FILLCELL_X4 FILLER_20_12 ();
 FILLCELL_X2 FILLER_20_16 ();
 FILLCELL_X1 FILLER_20_18 ();
 FILLCELL_X8 FILLER_20_22 ();
 FILLCELL_X2 FILLER_20_30 ();
 FILLCELL_X1 FILLER_20_35 ();
 FILLCELL_X32 FILLER_20_63 ();
 FILLCELL_X32 FILLER_20_95 ();
 FILLCELL_X16 FILLER_20_127 ();
 FILLCELL_X4 FILLER_20_143 ();
 FILLCELL_X8 FILLER_20_174 ();
 FILLCELL_X2 FILLER_20_182 ();
 FILLCELL_X1 FILLER_20_184 ();
 FILLCELL_X16 FILLER_20_212 ();
 FILLCELL_X4 FILLER_20_228 ();
 FILLCELL_X1 FILLER_20_232 ();
 FILLCELL_X1 FILLER_20_263 ();
 FILLCELL_X32 FILLER_21_37 ();
 FILLCELL_X4 FILLER_21_69 ();
 FILLCELL_X1 FILLER_21_73 ();
 FILLCELL_X32 FILLER_21_91 ();
 FILLCELL_X32 FILLER_21_123 ();
 FILLCELL_X32 FILLER_21_155 ();
 FILLCELL_X8 FILLER_21_187 ();
 FILLCELL_X4 FILLER_21_195 ();
 FILLCELL_X2 FILLER_21_199 ();
 FILLCELL_X2 FILLER_21_259 ();
 FILLCELL_X2 FILLER_22_13 ();
 FILLCELL_X8 FILLER_22_17 ();
 FILLCELL_X2 FILLER_22_25 ();
 FILLCELL_X4 FILLER_22_29 ();
 FILLCELL_X2 FILLER_22_63 ();
 FILLCELL_X1 FILLER_22_65 ();
 FILLCELL_X2 FILLER_22_68 ();
 FILLCELL_X2 FILLER_22_81 ();
 FILLCELL_X1 FILLER_22_83 ();
 FILLCELL_X32 FILLER_22_91 ();
 FILLCELL_X2 FILLER_22_123 ();
 FILLCELL_X8 FILLER_22_147 ();
 FILLCELL_X1 FILLER_22_155 ();
 FILLCELL_X4 FILLER_22_183 ();
 FILLCELL_X2 FILLER_22_187 ();
 FILLCELL_X1 FILLER_22_189 ();
 FILLCELL_X4 FILLER_22_195 ();
 FILLCELL_X1 FILLER_22_199 ();
 FILLCELL_X2 FILLER_22_205 ();
 FILLCELL_X2 FILLER_22_214 ();
 FILLCELL_X4 FILLER_22_253 ();
 FILLCELL_X1 FILLER_22_257 ();
 FILLCELL_X2 FILLER_23_16 ();
 FILLCELL_X16 FILLER_23_38 ();
 FILLCELL_X4 FILLER_23_54 ();
 FILLCELL_X8 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_100 ();
 FILLCELL_X8 FILLER_23_116 ();
 FILLCELL_X2 FILLER_23_124 ();
 FILLCELL_X2 FILLER_23_132 ();
 FILLCELL_X1 FILLER_23_134 ();
 FILLCELL_X8 FILLER_23_157 ();
 FILLCELL_X2 FILLER_23_165 ();
 FILLCELL_X16 FILLER_23_187 ();
 FILLCELL_X8 FILLER_23_203 ();
 FILLCELL_X2 FILLER_23_211 ();
 FILLCELL_X1 FILLER_23_213 ();
 FILLCELL_X2 FILLER_23_241 ();
 FILLCELL_X1 FILLER_23_263 ();
 FILLCELL_X1 FILLER_24_4 ();
 FILLCELL_X2 FILLER_24_33 ();
 FILLCELL_X1 FILLER_24_35 ();
 FILLCELL_X16 FILLER_24_63 ();
 FILLCELL_X4 FILLER_24_79 ();
 FILLCELL_X2 FILLER_24_83 ();
 FILLCELL_X8 FILLER_24_105 ();
 FILLCELL_X4 FILLER_24_113 ();
 FILLCELL_X1 FILLER_24_117 ();
 FILLCELL_X1 FILLER_24_133 ();
 FILLCELL_X16 FILLER_24_142 ();
 FILLCELL_X8 FILLER_24_158 ();
 FILLCELL_X2 FILLER_24_166 ();
 FILLCELL_X1 FILLER_24_168 ();
 FILLCELL_X4 FILLER_24_176 ();
 FILLCELL_X16 FILLER_24_212 ();
 FILLCELL_X8 FILLER_24_228 ();
 FILLCELL_X1 FILLER_24_263 ();
 FILLCELL_X2 FILLER_25_37 ();
 FILLCELL_X1 FILLER_25_39 ();
 FILLCELL_X16 FILLER_25_67 ();
 FILLCELL_X4 FILLER_25_83 ();
 FILLCELL_X2 FILLER_25_87 ();
 FILLCELL_X1 FILLER_25_89 ();
 FILLCELL_X16 FILLER_25_97 ();
 FILLCELL_X8 FILLER_25_113 ();
 FILLCELL_X2 FILLER_25_121 ();
 FILLCELL_X1 FILLER_25_123 ();
 FILLCELL_X32 FILLER_25_130 ();
 FILLCELL_X32 FILLER_25_162 ();
 FILLCELL_X32 FILLER_25_194 ();
 FILLCELL_X4 FILLER_25_246 ();
 FILLCELL_X1 FILLER_25_250 ();
 FILLCELL_X1 FILLER_25_257 ();
 FILLCELL_X4 FILLER_26_1 ();
 FILLCELL_X1 FILLER_26_5 ();
 FILLCELL_X1 FILLER_26_12 ();
 FILLCELL_X32 FILLER_26_21 ();
 FILLCELL_X8 FILLER_26_53 ();
 FILLCELL_X4 FILLER_26_61 ();
 FILLCELL_X4 FILLER_26_85 ();
 FILLCELL_X1 FILLER_26_89 ();
 FILLCELL_X4 FILLER_26_138 ();
 FILLCELL_X16 FILLER_26_169 ();
 FILLCELL_X8 FILLER_26_185 ();
 FILLCELL_X1 FILLER_26_193 ();
 FILLCELL_X16 FILLER_26_214 ();
 FILLCELL_X4 FILLER_26_230 ();
 FILLCELL_X2 FILLER_26_234 ();
 FILLCELL_X1 FILLER_26_257 ();
 FILLCELL_X16 FILLER_27_9 ();
 FILLCELL_X1 FILLER_27_28 ();
 FILLCELL_X16 FILLER_27_56 ();
 FILLCELL_X2 FILLER_27_72 ();
 FILLCELL_X4 FILLER_27_94 ();
 FILLCELL_X2 FILLER_27_98 ();
 FILLCELL_X1 FILLER_27_100 ();
 FILLCELL_X8 FILLER_27_121 ();
 FILLCELL_X2 FILLER_27_129 ();
 FILLCELL_X2 FILLER_27_134 ();
 FILLCELL_X1 FILLER_27_136 ();
 FILLCELL_X32 FILLER_27_139 ();
 FILLCELL_X2 FILLER_27_171 ();
 FILLCELL_X1 FILLER_27_173 ();
 FILLCELL_X16 FILLER_27_201 ();
 FILLCELL_X2 FILLER_27_217 ();
 FILLCELL_X1 FILLER_27_219 ();
 FILLCELL_X1 FILLER_27_243 ();
 FILLCELL_X1 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_30 ();
 FILLCELL_X16 FILLER_28_62 ();
 FILLCELL_X4 FILLER_28_80 ();
 FILLCELL_X2 FILLER_28_84 ();
 FILLCELL_X1 FILLER_28_93 ();
 FILLCELL_X1 FILLER_28_100 ();
 FILLCELL_X1 FILLER_28_103 ();
 FILLCELL_X8 FILLER_28_111 ();
 FILLCELL_X4 FILLER_28_141 ();
 FILLCELL_X4 FILLER_28_172 ();
 FILLCELL_X2 FILLER_28_183 ();
 FILLCELL_X32 FILLER_28_205 ();
 FILLCELL_X8 FILLER_29_70 ();
 FILLCELL_X2 FILLER_29_78 ();
 FILLCELL_X8 FILLER_29_86 ();
 FILLCELL_X1 FILLER_29_94 ();
 FILLCELL_X2 FILLER_29_98 ();
 FILLCELL_X16 FILLER_29_102 ();
 FILLCELL_X2 FILLER_29_118 ();
 FILLCELL_X32 FILLER_29_126 ();
 FILLCELL_X16 FILLER_29_158 ();
 FILLCELL_X8 FILLER_29_174 ();
 FILLCELL_X4 FILLER_29_182 ();
 FILLCELL_X2 FILLER_29_186 ();
 FILLCELL_X4 FILLER_29_195 ();
 FILLCELL_X4 FILLER_29_206 ();
 FILLCELL_X4 FILLER_29_230 ();
 FILLCELL_X2 FILLER_29_234 ();
 FILLCELL_X1 FILLER_29_236 ();
 FILLCELL_X2 FILLER_29_240 ();
 FILLCELL_X1 FILLER_29_242 ();
 FILLCELL_X1 FILLER_29_263 ();
 FILLCELL_X1 FILLER_30_18 ();
 FILLCELL_X32 FILLER_30_21 ();
 FILLCELL_X8 FILLER_30_53 ();
 FILLCELL_X4 FILLER_30_81 ();
 FILLCELL_X1 FILLER_30_87 ();
 FILLCELL_X16 FILLER_30_91 ();
 FILLCELL_X4 FILLER_30_107 ();
 FILLCELL_X1 FILLER_30_118 ();
 FILLCELL_X4 FILLER_30_122 ();
 FILLCELL_X4 FILLER_30_128 ();
 FILLCELL_X2 FILLER_30_132 ();
 FILLCELL_X2 FILLER_30_156 ();
 FILLCELL_X1 FILLER_30_158 ();
 FILLCELL_X1 FILLER_30_166 ();
 FILLCELL_X32 FILLER_30_187 ();
 FILLCELL_X16 FILLER_30_219 ();
 FILLCELL_X8 FILLER_30_242 ();
 FILLCELL_X4 FILLER_30_257 ();
 FILLCELL_X2 FILLER_31_4 ();
 FILLCELL_X8 FILLER_31_53 ();
 FILLCELL_X2 FILLER_31_61 ();
 FILLCELL_X1 FILLER_31_111 ();
 FILLCELL_X4 FILLER_31_132 ();
 FILLCELL_X2 FILLER_31_136 ();
 FILLCELL_X1 FILLER_31_146 ();
 FILLCELL_X16 FILLER_31_150 ();
 FILLCELL_X8 FILLER_31_166 ();
 FILLCELL_X2 FILLER_31_174 ();
 FILLCELL_X16 FILLER_31_216 ();
 FILLCELL_X1 FILLER_31_232 ();
 FILLCELL_X8 FILLER_31_253 ();
 FILLCELL_X2 FILLER_31_261 ();
 FILLCELL_X1 FILLER_31_263 ();
 FILLCELL_X16 FILLER_32_26 ();
 FILLCELL_X4 FILLER_32_42 ();
 FILLCELL_X2 FILLER_32_70 ();
 FILLCELL_X1 FILLER_32_72 ();
 FILLCELL_X4 FILLER_32_99 ();
 FILLCELL_X1 FILLER_32_103 ();
 FILLCELL_X2 FILLER_32_110 ();
 FILLCELL_X1 FILLER_32_114 ();
 FILLCELL_X2 FILLER_32_117 ();
 FILLCELL_X4 FILLER_32_161 ();
 FILLCELL_X2 FILLER_32_165 ();
 FILLCELL_X1 FILLER_32_167 ();
 FILLCELL_X8 FILLER_32_235 ();
 FILLCELL_X1 FILLER_32_263 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X16 FILLER_33_33 ();
 FILLCELL_X4 FILLER_33_49 ();
 FILLCELL_X2 FILLER_33_53 ();
 FILLCELL_X4 FILLER_33_85 ();
 FILLCELL_X1 FILLER_33_92 ();
 FILLCELL_X2 FILLER_33_102 ();
 FILLCELL_X1 FILLER_33_134 ();
 FILLCELL_X2 FILLER_33_147 ();
 FILLCELL_X1 FILLER_33_175 ();
 FILLCELL_X1 FILLER_33_183 ();
 FILLCELL_X1 FILLER_33_191 ();
 FILLCELL_X1 FILLER_33_199 ();
 FILLCELL_X1 FILLER_33_214 ();
 FILLCELL_X8 FILLER_33_255 ();
 FILLCELL_X1 FILLER_33_263 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X16 FILLER_34_33 ();
 FILLCELL_X8 FILLER_34_49 ();
 FILLCELL_X4 FILLER_34_57 ();
 FILLCELL_X1 FILLER_34_61 ();
 FILLCELL_X2 FILLER_34_77 ();
 FILLCELL_X2 FILLER_34_91 ();
 FILLCELL_X1 FILLER_34_93 ();
 FILLCELL_X1 FILLER_34_99 ();
 FILLCELL_X4 FILLER_34_133 ();
 FILLCELL_X1 FILLER_34_143 ();
 FILLCELL_X2 FILLER_34_149 ();
 FILLCELL_X2 FILLER_34_154 ();
 FILLCELL_X1 FILLER_34_156 ();
 FILLCELL_X2 FILLER_34_200 ();
 FILLCELL_X8 FILLER_34_211 ();
 FILLCELL_X4 FILLER_34_219 ();
 FILLCELL_X2 FILLER_34_236 ();
 FILLCELL_X1 FILLER_34_238 ();
 FILLCELL_X8 FILLER_34_249 ();
 FILLCELL_X4 FILLER_34_257 ();
 FILLCELL_X2 FILLER_34_261 ();
 FILLCELL_X1 FILLER_34_263 ();
endmodule
