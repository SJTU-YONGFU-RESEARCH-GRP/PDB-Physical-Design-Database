module booth_multiplier (clk,
    done,
    rst,
    start,
    multiplicand,
    multiplier,
    product);
 input clk;
 output done;
 input rst;
 input start;
 input [7:0] multiplicand;
 input [7:0] multiplier;
 output [15:0] product;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire start_r;
 wire state;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net34;

 sky130_fd_sc_hd__inv_1 _400_ (.A(state),
    .Y(_018_));
 sky130_fd_sc_hd__nand2_2 _401_ (.A(_018_),
    .B(_306_),
    .Y(_019_));
 sky130_fd_sc_hd__clkbuf_4 _402_ (.A(_019_),
    .X(_020_));
 sky130_fd_sc_hd__o21ai_0 _403_ (.A1(_018_),
    .A2(net17),
    .B1(_020_),
    .Y(_399_));
 sky130_fd_sc_hd__clkbuf_4 _404_ (.A(net8),
    .X(_021_));
 sky130_fd_sc_hd__and2_0 _405_ (.A(_021_),
    .B(net2),
    .X(_309_));
 sky130_fd_sc_hd__clkbuf_4 _406_ (.A(multiplier[1]),
    .X(_022_));
 sky130_fd_sc_hd__and2_0 _407_ (.A(net1),
    .B(_022_),
    .X(_308_));
 sky130_fd_sc_hd__nand2_1 _408_ (.A(net1),
    .B(net9),
    .Y(_106_));
 sky130_fd_sc_hd__nand2_1 _409_ (.A(_021_),
    .B(net4),
    .Y(_113_));
 sky130_fd_sc_hd__nand2_1 _410_ (.A(_022_),
    .B(net3),
    .Y(_112_));
 sky130_fd_sc_hd__nand2_1 _411_ (.A(net2),
    .B(net9),
    .Y(_111_));
 sky130_fd_sc_hd__nand2_1 _412_ (.A(net1),
    .B(net10),
    .Y(_116_));
 sky130_fd_sc_hd__nand2_1 _413_ (.A(_021_),
    .B(net5),
    .Y(_120_));
 sky130_fd_sc_hd__nand2_1 _414_ (.A(_022_),
    .B(net4),
    .Y(_119_));
 sky130_fd_sc_hd__nand2_1 _415_ (.A(net3),
    .B(net9),
    .Y(_121_));
 sky130_fd_sc_hd__and2_0 _416_ (.A(net2),
    .B(net10),
    .X(_319_));
 sky130_fd_sc_hd__and2_0 _417_ (.A(net1),
    .B(net11),
    .X(_318_));
 sky130_fd_sc_hd__nand2_1 _418_ (.A(_021_),
    .B(net7),
    .Y(_129_));
 sky130_fd_sc_hd__nand2_1 _419_ (.A(_022_),
    .B(net6),
    .Y(_128_));
 sky130_fd_sc_hd__nand2_1 _420_ (.A(net9),
    .B(net5),
    .Y(_127_));
 sky130_fd_sc_hd__and2_0 _421_ (.A(_022_),
    .B(net5),
    .X(_141_));
 sky130_fd_sc_hd__and2_0 _422_ (.A(net9),
    .B(net4),
    .X(_140_));
 sky130_fd_sc_hd__and2_0 _423_ (.A(net4),
    .B(net10),
    .X(_134_));
 sky130_fd_sc_hd__and2_0 _424_ (.A(net3),
    .B(net11),
    .X(_133_));
 sky130_fd_sc_hd__and2_0 _425_ (.A(net2),
    .B(net12),
    .X(_132_));
 sky130_fd_sc_hd__and2_0 _426_ (.A(net1),
    .B(net13),
    .X(_328_));
 sky130_fd_sc_hd__nand2_1 _427_ (.A(_022_),
    .B(net7),
    .Y(_167_));
 sky130_fd_sc_hd__nand2_1 _428_ (.A(net9),
    .B(net6),
    .Y(_173_));
 sky130_fd_sc_hd__nand2_1 _429_ (.A(net10),
    .B(net5),
    .Y(_171_));
 sky130_fd_sc_hd__nand2_1 _430_ (.A(net4),
    .B(net11),
    .Y(_172_));
 sky130_fd_sc_hd__and2_0 _431_ (.A(net3),
    .B(net12),
    .X(_178_));
 sky130_fd_sc_hd__and2_0 _432_ (.A(net2),
    .B(net13),
    .X(_180_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(net14),
    .Y(_166_));
 sky130_fd_sc_hd__nor2_1 _434_ (.A(net1),
    .B(_166_),
    .Y(_179_));
 sky130_fd_sc_hd__inv_1 _435_ (.A(_190_),
    .Y(_187_));
 sky130_fd_sc_hd__and2_0 _436_ (.A(net9),
    .B(net7),
    .X(_344_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(net10),
    .B(net6),
    .Y(_193_));
 sky130_fd_sc_hd__nand2_1 _438_ (.A(net5),
    .B(net11),
    .Y(_192_));
 sky130_fd_sc_hd__nand2_1 _439_ (.A(net4),
    .B(net12),
    .Y(_191_));
 sky130_fd_sc_hd__and2_0 _440_ (.A(net3),
    .B(net13),
    .X(_348_));
 sky130_fd_sc_hd__nor2_1 _441_ (.A(net2),
    .B(_166_),
    .Y(_349_));
 sky130_fd_sc_hd__buf_2 _442_ (.A(multiplicand[7]),
    .X(_023_));
 sky130_fd_sc_hd__and2_0 _443_ (.A(net9),
    .B(_023_),
    .X(_354_));
 sky130_fd_sc_hd__a31oi_2 _444_ (.A1(_021_),
    .A2(_022_),
    .A3(_023_),
    .B1(_346_),
    .Y(_216_));
 sky130_fd_sc_hd__nand2_1 _445_ (.A(net10),
    .B(net7),
    .Y(_211_));
 sky130_fd_sc_hd__nand2_1 _446_ (.A(net11),
    .B(net6),
    .Y(_212_));
 sky130_fd_sc_hd__nand2_1 _447_ (.A(net5),
    .B(net12),
    .Y(_210_));
 sky130_fd_sc_hd__and2_0 _448_ (.A(net4),
    .B(net13),
    .X(_358_));
 sky130_fd_sc_hd__nor2_1 _449_ (.A(net3),
    .B(_166_),
    .Y(_357_));
 sky130_fd_sc_hd__a31oi_4 _450_ (.A1(_021_),
    .A2(_022_),
    .A3(_023_),
    .B1(_355_),
    .Y(_234_));
 sky130_fd_sc_hd__and2_2 _451_ (.A(net10),
    .B(_023_),
    .X(_229_));
 sky130_fd_sc_hd__and2_0 _452_ (.A(net11),
    .B(net7),
    .X(_230_));
 sky130_fd_sc_hd__and2_0 _453_ (.A(net6),
    .B(net12),
    .X(_231_));
 sky130_fd_sc_hd__and2_0 _454_ (.A(net5),
    .B(net13),
    .X(_362_));
 sky130_fd_sc_hd__nor2_1 _455_ (.A(net4),
    .B(_166_),
    .Y(_363_));
 sky130_fd_sc_hd__inv_1 _456_ (.A(_339_),
    .Y(_163_));
 sky130_fd_sc_hd__and2_0 _457_ (.A(net11),
    .B(_023_),
    .X(_250_));
 sky130_fd_sc_hd__and2_0 _458_ (.A(net7),
    .B(net12),
    .X(_249_));
 sky130_fd_sc_hd__and2_0 _459_ (.A(net6),
    .B(net13),
    .X(_369_));
 sky130_fd_sc_hd__nor2_1 _460_ (.A(net5),
    .B(_166_),
    .Y(_368_));
 sky130_fd_sc_hd__and2_0 _461_ (.A(net12),
    .B(_023_),
    .X(_266_));
 sky130_fd_sc_hd__and2_0 _462_ (.A(net7),
    .B(net13),
    .X(_375_));
 sky130_fd_sc_hd__nor2_1 _463_ (.A(net6),
    .B(_166_),
    .Y(_376_));
 sky130_fd_sc_hd__and2_0 _464_ (.A(net13),
    .B(_023_),
    .X(_384_));
 sky130_fd_sc_hd__nor2_1 _465_ (.A(net7),
    .B(_166_),
    .Y(_385_));
 sky130_fd_sc_hd__inv_6 _466_ (.A(net15),
    .Y(_000_));
 sky130_fd_sc_hd__nand2_1 _467_ (.A(net1),
    .B(net12),
    .Y(_145_));
 sky130_fd_sc_hd__inv_1 _468_ (.A(_320_),
    .Y(_158_));
 sky130_fd_sc_hd__nand2_1 _469_ (.A(net2),
    .B(_022_),
    .Y(_107_));
 sky130_fd_sc_hd__nand2_1 _470_ (.A(net2),
    .B(net11),
    .Y(_146_));
 sky130_fd_sc_hd__nand2_1 _471_ (.A(_021_),
    .B(net3),
    .Y(_108_));
 sky130_fd_sc_hd__nand2_1 _472_ (.A(net3),
    .B(net10),
    .Y(_147_));
 sky130_fd_sc_hd__nand2_1 _473_ (.A(_021_),
    .B(_023_),
    .Y(_168_));
 sky130_fd_sc_hd__inv_1 _474_ (.A(_144_),
    .Y(_156_));
 sky130_fd_sc_hd__inv_1 _475_ (.A(_154_),
    .Y(_331_));
 sky130_fd_sc_hd__inv_1 _476_ (.A(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__inv_1 _477_ (.A(_233_),
    .Y(_235_));
 sky130_fd_sc_hd__inv_1 _478_ (.A(_242_),
    .Y(_243_));
 sky130_fd_sc_hd__inv_1 _479_ (.A(_252_),
    .Y(_253_));
 sky130_fd_sc_hd__inv_1 _480_ (.A(_259_),
    .Y(_260_));
 sky130_fd_sc_hd__inv_1 _481_ (.A(_268_),
    .Y(_269_));
 sky130_fd_sc_hd__inv_1 _482_ (.A(_275_),
    .Y(_276_));
 sky130_fd_sc_hd__inv_1 _483_ (.A(_285_),
    .Y(_286_));
 sky130_fd_sc_hd__inv_1 _484_ (.A(_295_),
    .Y(_296_));
 sky130_fd_sc_hd__inv_1 _485_ (.A(_143_),
    .Y(_137_));
 sky130_fd_sc_hd__inv_1 _486_ (.A(_153_),
    .Y(_186_));
 sky130_fd_sc_hd__inv_1 _487_ (.A(_181_),
    .Y(_199_));
 sky130_fd_sc_hd__inv_1 _488_ (.A(_222_),
    .Y(_246_));
 sky130_fd_sc_hd__inv_1 _489_ (.A(_241_),
    .Y(_263_));
 sky130_fd_sc_hd__inv_1 _490_ (.A(_258_),
    .Y(_279_));
 sky130_fd_sc_hd__inv_1 _491_ (.A(_274_),
    .Y(_289_));
 sky130_fd_sc_hd__inv_1 _492_ (.A(_284_),
    .Y(_299_));
 sky130_fd_sc_hd__inv_1 _493_ (.A(net16),
    .Y(_302_));
 sky130_fd_sc_hd__inv_1 _494_ (.A(_117_),
    .Y(_322_));
 sky130_fd_sc_hd__inv_1 _495_ (.A(_122_),
    .Y(_155_));
 sky130_fd_sc_hd__inv_1 _496_ (.A(_159_),
    .Y(_330_));
 sky130_fd_sc_hd__inv_1 _497_ (.A(_189_),
    .Y(_341_));
 sky130_fd_sc_hd__inv_1 _498_ (.A(_204_),
    .Y(_205_));
 sky130_fd_sc_hd__inv_1 _499_ (.A(_188_),
    .Y(_351_));
 sky130_fd_sc_hd__inv_1 _500_ (.A(_194_),
    .Y(_219_));
 sky130_fd_sc_hd__inv_1 _501_ (.A(_248_),
    .Y(_364_));
 sky130_fd_sc_hd__inv_1 _502_ (.A(_265_),
    .Y(_370_));
 sky130_fd_sc_hd__inv_1 _503_ (.A(_271_),
    .Y(_374_));
 sky130_fd_sc_hd__inv_1 _504_ (.A(_281_),
    .Y(_377_));
 sky130_fd_sc_hd__inv_1 _505_ (.A(_280_),
    .Y(_386_));
 sky130_fd_sc_hd__inv_1 _506_ (.A(_301_),
    .Y(_394_));
 sky130_fd_sc_hd__inv_1 _507_ (.A(start_r),
    .Y(_305_));
 sky130_fd_sc_hd__inv_1 _508_ (.A(_110_),
    .Y(_312_));
 sky130_fd_sc_hd__inv_1 _509_ (.A(_118_),
    .Y(_315_));
 sky130_fd_sc_hd__inv_1 _510_ (.A(_126_),
    .Y(_323_));
 sky130_fd_sc_hd__and2_0 _511_ (.A(_021_),
    .B(net6),
    .X(_142_));
 sky130_fd_sc_hd__inv_1 _512_ (.A(_139_),
    .Y(_152_));
 sky130_fd_sc_hd__inv_1 _513_ (.A(_148_),
    .Y(_329_));
 sky130_fd_sc_hd__inv_1 _514_ (.A(_160_),
    .Y(_337_));
 sky130_fd_sc_hd__inv_1 _515_ (.A(_184_),
    .Y(_206_));
 sky130_fd_sc_hd__xor2_1 _516_ (.A(net8),
    .B(_022_),
    .X(_024_));
 sky130_fd_sc_hd__and2_0 _517_ (.A(_023_),
    .B(_024_),
    .X(_345_));
 sky130_fd_sc_hd__inv_1 _518_ (.A(_228_),
    .Y(_359_));
 sky130_fd_sc_hd__inv_1 _519_ (.A(_213_),
    .Y(_240_));
 sky130_fd_sc_hd__inv_1 _520_ (.A(_227_),
    .Y(_365_));
 sky130_fd_sc_hd__inv_1 _521_ (.A(_247_),
    .Y(_371_));
 sky130_fd_sc_hd__inv_1 _522_ (.A(_264_),
    .Y(_378_));
 sky130_fd_sc_hd__inv_1 _523_ (.A(_270_),
    .Y(_381_));
 sky130_fd_sc_hd__inv_1 _524_ (.A(_291_),
    .Y(_387_));
 sky130_fd_sc_hd__nor2_1 _525_ (.A(_023_),
    .B(_166_),
    .Y(_390_));
 sky130_fd_sc_hd__inv_1 _526_ (.A(_290_),
    .Y(_395_));
 sky130_fd_sc_hd__inv_1 _527_ (.A(_333_),
    .Y(_162_));
 sky130_fd_sc_hd__inv_1 _528_ (.A(_340_),
    .Y(_183_));
 sky130_fd_sc_hd__inv_1 _529_ (.A(_347_),
    .Y(_196_));
 sky130_fd_sc_hd__inv_2 _530_ (.A(_356_),
    .Y(_215_));
 sky130_fd_sc_hd__inv_1 _531_ (.A(_321_),
    .Y(_124_));
 sky130_fd_sc_hd__inv_1 _532_ (.A(_350_),
    .Y(_200_));
 sky130_fd_sc_hd__inv_1 _533_ (.A(_334_),
    .Y(_161_));
 sky130_fd_sc_hd__nand3_1 _534_ (.A(_018_),
    .B(net17),
    .C(_304_),
    .Y(_025_));
 sky130_fd_sc_hd__o21ai_0 _535_ (.A1(_018_),
    .A2(_303_),
    .B1(_025_),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_1 _536_ (.A(net18),
    .B(_020_),
    .Y(_026_));
 sky130_fd_sc_hd__nor2b_1 _537_ (.A(state),
    .B_N(_306_),
    .Y(_027_));
 sky130_fd_sc_hd__clkbuf_4 _538_ (.A(_027_),
    .X(_028_));
 sky130_fd_sc_hd__nand3_1 _539_ (.A(_021_),
    .B(net1),
    .C(_028_),
    .Y(_029_));
 sky130_fd_sc_hd__nand2_1 _540_ (.A(_026_),
    .B(_029_),
    .Y(_002_));
 sky130_fd_sc_hd__clkbuf_2 _541_ (.A(_019_),
    .X(_030_));
 sky130_fd_sc_hd__a211oi_1 _542_ (.A1(_336_),
    .A2(_339_),
    .B1(_335_),
    .C1(_342_),
    .Y(_031_));
 sky130_fd_sc_hd__o21ai_0 _543_ (.A1(_343_),
    .A2(_342_),
    .B1(_353_),
    .Y(_032_));
 sky130_fd_sc_hd__o21bai_1 _544_ (.A1(_031_),
    .A2(_032_),
    .B1_N(_352_),
    .Y(_033_));
 sky130_fd_sc_hd__a21oi_1 _545_ (.A1(_361_),
    .A2(_033_),
    .B1(_360_),
    .Y(_034_));
 sky130_fd_sc_hd__xor2_1 _546_ (.A(_367_),
    .B(_034_),
    .X(_035_));
 sky130_fd_sc_hd__nand2_1 _547_ (.A(net19),
    .B(_030_),
    .Y(_036_));
 sky130_fd_sc_hd__o21ai_0 _548_ (.A1(_030_),
    .A2(_035_),
    .B1(_036_),
    .Y(_003_));
 sky130_fd_sc_hd__clkbuf_2 _549_ (.A(_373_),
    .X(_037_));
 sky130_fd_sc_hd__nor2b_1 _550_ (.A(_164_),
    .B_N(_343_),
    .Y(_038_));
 sky130_fd_sc_hd__o21a_1 _551_ (.A1(_353_),
    .A2(_352_),
    .B1(_361_),
    .X(_039_));
 sky130_fd_sc_hd__o31a_1 _552_ (.A1(_342_),
    .A2(_352_),
    .A3(_038_),
    .B1(_039_),
    .X(_040_));
 sky130_fd_sc_hd__o21a_1 _553_ (.A1(_360_),
    .A2(_040_),
    .B1(_367_),
    .X(_041_));
 sky130_fd_sc_hd__nor3_1 _554_ (.A(_037_),
    .B(_366_),
    .C(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__o21a_1 _555_ (.A1(_366_),
    .A2(_041_),
    .B1(_037_),
    .X(_043_));
 sky130_fd_sc_hd__nand2_1 _556_ (.A(net20),
    .B(_020_),
    .Y(_044_));
 sky130_fd_sc_hd__o31ai_1 _557_ (.A1(_019_),
    .A2(_042_),
    .A3(_043_),
    .B1(_044_),
    .Y(_004_));
 sky130_fd_sc_hd__clkbuf_2 _558_ (.A(_380_),
    .X(_045_));
 sky130_fd_sc_hd__and3_1 _559_ (.A(_361_),
    .B(_367_),
    .C(_037_),
    .X(_046_));
 sky130_fd_sc_hd__a21oi_1 _560_ (.A1(_037_),
    .A2(_366_),
    .B1(_372_),
    .Y(_047_));
 sky130_fd_sc_hd__nand3_1 _561_ (.A(_367_),
    .B(_037_),
    .C(_360_),
    .Y(_048_));
 sky130_fd_sc_hd__nand2_1 _562_ (.A(_047_),
    .B(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__a21oi_1 _563_ (.A1(_033_),
    .A2(_046_),
    .B1(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__xor2_1 _564_ (.A(_045_),
    .B(_050_),
    .X(_051_));
 sky130_fd_sc_hd__nand2_1 _565_ (.A(net21),
    .B(_030_),
    .Y(_052_));
 sky130_fd_sc_hd__o21ai_0 _566_ (.A1(_030_),
    .A2(_051_),
    .B1(_052_),
    .Y(_005_));
 sky130_fd_sc_hd__o2111ai_1 _567_ (.A1(_360_),
    .A2(_040_),
    .B1(_367_),
    .C1(_037_),
    .D1(_045_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2b_1 _568_ (.A(_047_),
    .B_N(_045_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _569_ (.A(_379_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__a211o_1 _570_ (.A1(_053_),
    .A2(_055_),
    .B1(_389_),
    .C1(_019_),
    .X(_056_));
 sky130_fd_sc_hd__nand4_1 _571_ (.A(_389_),
    .B(_028_),
    .C(_053_),
    .D(_055_),
    .Y(_057_));
 sky130_fd_sc_hd__nand2_1 _572_ (.A(net22),
    .B(_030_),
    .Y(_058_));
 sky130_fd_sc_hd__nand3_1 _573_ (.A(_056_),
    .B(_057_),
    .C(_058_),
    .Y(_006_));
 sky130_fd_sc_hd__nor2_1 _574_ (.A(net23),
    .B(_028_),
    .Y(_059_));
 sky130_fd_sc_hd__nand4_1 _575_ (.A(_367_),
    .B(_037_),
    .C(_045_),
    .D(_389_),
    .Y(_060_));
 sky130_fd_sc_hd__nand2_1 _576_ (.A(_397_),
    .B(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__nand2_1 _577_ (.A(_045_),
    .B(_389_),
    .Y(_062_));
 sky130_fd_sc_hd__a21oi_1 _578_ (.A1(_389_),
    .A2(_379_),
    .B1(_388_),
    .Y(_063_));
 sky130_fd_sc_hd__o21ai_1 _579_ (.A1(_047_),
    .A2(_062_),
    .B1(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__mux2i_1 _580_ (.A0(_061_),
    .A1(_397_),
    .S(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__nor2_1 _581_ (.A(_019_),
    .B(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__nor2_1 _582_ (.A(_397_),
    .B(_060_),
    .Y(_067_));
 sky130_fd_sc_hd__inv_1 _583_ (.A(_397_),
    .Y(_068_));
 sky130_fd_sc_hd__nor2_1 _584_ (.A(_068_),
    .B(_064_),
    .Y(_069_));
 sky130_fd_sc_hd__mux2i_1 _585_ (.A0(_067_),
    .A1(_069_),
    .S(_034_),
    .Y(_070_));
 sky130_fd_sc_hd__o22ai_1 _586_ (.A1(_059_),
    .A2(_066_),
    .B1(_070_),
    .B2(_020_),
    .Y(_007_));
 sky130_fd_sc_hd__nand4_1 _587_ (.A(_037_),
    .B(_045_),
    .C(_389_),
    .D(_397_),
    .Y(_071_));
 sky130_fd_sc_hd__nor2_1 _588_ (.A(_367_),
    .B(_366_),
    .Y(_072_));
 sky130_fd_sc_hd__nor2_1 _589_ (.A(_071_),
    .B(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__o31ai_1 _590_ (.A1(_360_),
    .A2(_366_),
    .A3(_040_),
    .B1(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__a21o_1 _591_ (.A1(_045_),
    .A2(_372_),
    .B1(_379_),
    .X(_075_));
 sky130_fd_sc_hd__nand3_1 _592_ (.A(_389_),
    .B(_397_),
    .C(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__a21oi_1 _593_ (.A1(_397_),
    .A2(_388_),
    .B1(_396_),
    .Y(_077_));
 sky130_fd_sc_hd__xor2_1 _594_ (.A(_294_),
    .B(_393_),
    .X(_078_));
 sky130_fd_sc_hd__xnor2_1 _595_ (.A(_297_),
    .B(_300_),
    .Y(_079_));
 sky130_fd_sc_hd__xnor2_1 _596_ (.A(_078_),
    .B(_079_),
    .Y(_080_));
 sky130_fd_sc_hd__xnor2_1 _597_ (.A(_391_),
    .B(_383_),
    .Y(_081_));
 sky130_fd_sc_hd__xnor2_1 _598_ (.A(_080_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__a31o_1 _599_ (.A1(_074_),
    .A2(_076_),
    .A3(_077_),
    .B1(_082_),
    .X(_083_));
 sky130_fd_sc_hd__nand4_1 _600_ (.A(_082_),
    .B(_074_),
    .C(_076_),
    .D(_077_),
    .Y(_084_));
 sky130_fd_sc_hd__nor2_1 _601_ (.A(net24),
    .B(_028_),
    .Y(_085_));
 sky130_fd_sc_hd__a31oi_1 _602_ (.A1(_028_),
    .A2(_083_),
    .A3(_084_),
    .B1(_085_),
    .Y(_008_));
 sky130_fd_sc_hd__nand2_1 _603_ (.A(_311_),
    .B(_028_),
    .Y(_086_));
 sky130_fd_sc_hd__nand2_1 _604_ (.A(net25),
    .B(_020_),
    .Y(_087_));
 sky130_fd_sc_hd__nand2_1 _605_ (.A(_086_),
    .B(_087_),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_1 _606_ (.A(_314_),
    .B(_028_),
    .Y(_088_));
 sky130_fd_sc_hd__nand2_1 _607_ (.A(net26),
    .B(_020_),
    .Y(_089_));
 sky130_fd_sc_hd__nand2_1 _608_ (.A(_088_),
    .B(_089_),
    .Y(_010_));
 sky130_fd_sc_hd__nand2_1 _609_ (.A(_317_),
    .B(_028_),
    .Y(_090_));
 sky130_fd_sc_hd__nand2_1 _610_ (.A(net27),
    .B(_020_),
    .Y(_091_));
 sky130_fd_sc_hd__nand2_1 _611_ (.A(_090_),
    .B(_091_),
    .Y(_011_));
 sky130_fd_sc_hd__nand2_1 _612_ (.A(_327_),
    .B(_028_),
    .Y(_092_));
 sky130_fd_sc_hd__nand2_1 _613_ (.A(net28),
    .B(_020_),
    .Y(_093_));
 sky130_fd_sc_hd__nand2_1 _614_ (.A(_092_),
    .B(_093_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_1 _615_ (.A(_398_),
    .B(_028_),
    .Y(_094_));
 sky130_fd_sc_hd__nand2_1 _616_ (.A(net29),
    .B(_020_),
    .Y(_095_));
 sky130_fd_sc_hd__nand2_1 _617_ (.A(_094_),
    .B(_095_),
    .Y(_013_));
 sky130_fd_sc_hd__nand2_1 _618_ (.A(net30),
    .B(_030_),
    .Y(_096_));
 sky130_fd_sc_hd__o21ai_0 _619_ (.A1(_165_),
    .A2(_020_),
    .B1(_096_),
    .Y(_014_));
 sky130_fd_sc_hd__xor2_1 _620_ (.A(_343_),
    .B(_164_),
    .X(_097_));
 sky130_fd_sc_hd__nand2_1 _621_ (.A(net31),
    .B(_030_),
    .Y(_098_));
 sky130_fd_sc_hd__o21ai_0 _622_ (.A1(_030_),
    .A2(_097_),
    .B1(_098_),
    .Y(_015_));
 sky130_fd_sc_hd__a21o_1 _623_ (.A1(_336_),
    .A2(_339_),
    .B1(_335_),
    .X(_099_));
 sky130_fd_sc_hd__a21oi_1 _624_ (.A1(_343_),
    .A2(_099_),
    .B1(_342_),
    .Y(_100_));
 sky130_fd_sc_hd__xor2_1 _625_ (.A(_353_),
    .B(_100_),
    .X(_101_));
 sky130_fd_sc_hd__nand2_1 _626_ (.A(net32),
    .B(_030_),
    .Y(_102_));
 sky130_fd_sc_hd__o21ai_0 _627_ (.A1(_030_),
    .A2(_101_),
    .B1(_102_),
    .Y(_016_));
 sky130_fd_sc_hd__o21ai_0 _628_ (.A1(_342_),
    .A2(_038_),
    .B1(_353_),
    .Y(_103_));
 sky130_fd_sc_hd__nor2_1 _629_ (.A(_361_),
    .B(_352_),
    .Y(_104_));
 sky130_fd_sc_hd__a211oi_1 _630_ (.A1(_103_),
    .A2(_104_),
    .B1(_040_),
    .C1(_019_),
    .Y(_105_));
 sky130_fd_sc_hd__a21o_1 _631_ (.A1(net33),
    .A2(_019_),
    .B1(_105_),
    .X(_017_));
 sky130_fd_sc_hd__fa_1 _632_ (.A(_106_),
    .B(_107_),
    .CIN(_108_),
    .COUT(_109_),
    .SUM(_110_));
 sky130_fd_sc_hd__fa_1 _633_ (.A(_111_),
    .B(_112_),
    .CIN(_113_),
    .COUT(_114_),
    .SUM(_115_));
 sky130_fd_sc_hd__fa_1 _634_ (.A(_116_),
    .B(_109_),
    .CIN(_115_),
    .COUT(_117_),
    .SUM(_118_));
 sky130_fd_sc_hd__fa_1 _635_ (.A(_119_),
    .B(_120_),
    .CIN(_121_),
    .COUT(_122_),
    .SUM(_123_));
 sky130_fd_sc_hd__fa_1 _636_ (.A(_124_),
    .B(_114_),
    .CIN(_123_),
    .COUT(_125_),
    .SUM(_126_));
 sky130_fd_sc_hd__fa_1 _637_ (.A(_127_),
    .B(_128_),
    .CIN(_129_),
    .COUT(_130_),
    .SUM(_131_));
 sky130_fd_sc_hd__fa_1 _638_ (.A(_132_),
    .B(_133_),
    .CIN(_134_),
    .COUT(_135_),
    .SUM(_136_));
 sky130_fd_sc_hd__fa_1 _639_ (.A(_136_),
    .B(_137_),
    .CIN(_131_),
    .COUT(_138_),
    .SUM(_139_));
 sky130_fd_sc_hd__fa_1 _640_ (.A(_140_),
    .B(_141_),
    .CIN(_142_),
    .COUT(_143_),
    .SUM(_144_));
 sky130_fd_sc_hd__fa_1 _641_ (.A(_145_),
    .B(_146_),
    .CIN(_147_),
    .COUT(_148_),
    .SUM(_149_));
 sky130_fd_sc_hd__fa_1 _642_ (.A(_150_),
    .B(_151_),
    .CIN(_152_),
    .COUT(_153_),
    .SUM(_154_));
 sky130_fd_sc_hd__fa_1 _643_ (.A(_149_),
    .B(_155_),
    .CIN(_156_),
    .COUT(_150_),
    .SUM(_157_));
 sky130_fd_sc_hd__fa_1 _644_ (.A(_158_),
    .B(_125_),
    .CIN(_157_),
    .COUT(_159_),
    .SUM(_160_));
 sky130_fd_sc_hd__fa_1 _645_ (.A(_161_),
    .B(_162_),
    .CIN(_163_),
    .COUT(_164_),
    .SUM(_165_));
 sky130_fd_sc_hd__fa_1 _646_ (.A(_166_),
    .B(_167_),
    .CIN(_168_),
    .COUT(_169_),
    .SUM(_170_));
 sky130_fd_sc_hd__fa_1 _647_ (.A(_171_),
    .B(_172_),
    .CIN(_173_),
    .COUT(_174_),
    .SUM(_175_));
 sky130_fd_sc_hd__fa_1 _648_ (.A(_170_),
    .B(_130_),
    .CIN(_175_),
    .COUT(_176_),
    .SUM(_177_));
 sky130_fd_sc_hd__fa_1 _649_ (.A(_178_),
    .B(_179_),
    .CIN(_180_),
    .COUT(_181_),
    .SUM(_182_));
 sky130_fd_sc_hd__fa_1 _650_ (.A(_138_),
    .B(_177_),
    .CIN(_183_),
    .COUT(_184_),
    .SUM(_185_));
 sky130_fd_sc_hd__fa_1 _651_ (.A(_186_),
    .B(_187_),
    .CIN(_185_),
    .COUT(_188_),
    .SUM(_189_));
 sky130_fd_sc_hd__fa_1 _652_ (.A(_191_),
    .B(_192_),
    .CIN(_193_),
    .COUT(_194_),
    .SUM(_195_));
 sky130_fd_sc_hd__fa_1 _653_ (.A(_195_),
    .B(_196_),
    .CIN(_169_),
    .COUT(_197_),
    .SUM(_198_));
 sky130_fd_sc_hd__fa_1 _654_ (.A(_199_),
    .B(_174_),
    .CIN(_200_),
    .COUT(_201_),
    .SUM(_202_));
 sky130_fd_sc_hd__fa_1 _655_ (.A(_202_),
    .B(_176_),
    .CIN(_198_),
    .COUT(_203_),
    .SUM(_204_));
 sky130_fd_sc_hd__fa_1 _656_ (.A(_205_),
    .B(_206_),
    .CIN(_207_),
    .COUT(_208_),
    .SUM(_209_));
 sky130_fd_sc_hd__fa_1 _657_ (.A(_210_),
    .B(_211_),
    .CIN(_212_),
    .COUT(_213_),
    .SUM(_214_));
 sky130_fd_sc_hd__fa_1 _658_ (.A(_214_),
    .B(_215_),
    .CIN(_216_),
    .COUT(_217_),
    .SUM(_218_));
 sky130_fd_sc_hd__fa_1 _659_ (.A(_219_),
    .B(_220_),
    .CIN(_221_),
    .COUT(_222_),
    .SUM(_223_));
 sky130_fd_sc_hd__fa_1 _660_ (.A(_218_),
    .B(_197_),
    .CIN(_224_),
    .COUT(_225_),
    .SUM(_226_));
 sky130_fd_sc_hd__fa_1 _661_ (.A(_201_),
    .B(_203_),
    .CIN(_226_),
    .COUT(_227_),
    .SUM(_228_));
 sky130_fd_sc_hd__fa_1 _662_ (.A(_229_),
    .B(_230_),
    .CIN(_231_),
    .COUT(_232_),
    .SUM(_233_));
 sky130_fd_sc_hd__fa_1 _663_ (.A(_234_),
    .B(_235_),
    .CIN(_215_),
    .COUT(_236_),
    .SUM(_237_));
 sky130_fd_sc_hd__fa_1 _664_ (.A(_238_),
    .B(_239_),
    .CIN(_240_),
    .COUT(_241_),
    .SUM(_242_));
 sky130_fd_sc_hd__fa_1 _665_ (.A(_237_),
    .B(_217_),
    .CIN(_243_),
    .COUT(_244_),
    .SUM(_245_));
 sky130_fd_sc_hd__fa_1 _666_ (.A(_225_),
    .B(_246_),
    .CIN(_245_),
    .COUT(_247_),
    .SUM(_248_));
 sky130_fd_sc_hd__fa_1 _667_ (.A(_229_),
    .B(_249_),
    .CIN(_250_),
    .COUT(_251_),
    .SUM(_252_));
 sky130_fd_sc_hd__fa_1 _668_ (.A(_234_),
    .B(_215_),
    .CIN(_253_),
    .COUT(_254_),
    .SUM(_255_));
 sky130_fd_sc_hd__fa_1 _669_ (.A(_256_),
    .B(_232_),
    .CIN(_257_),
    .COUT(_258_),
    .SUM(_259_));
 sky130_fd_sc_hd__fa_1 _670_ (.A(_260_),
    .B(_236_),
    .CIN(_255_),
    .COUT(_261_),
    .SUM(_262_));
 sky130_fd_sc_hd__fa_1 _671_ (.A(_262_),
    .B(_244_),
    .CIN(_263_),
    .COUT(_264_),
    .SUM(_265_));
 sky130_fd_sc_hd__fa_2 _672_ (.A(_229_),
    .B(_266_),
    .CIN(_250_),
    .COUT(_267_),
    .SUM(_268_));
 sky130_fd_sc_hd__fa_4 _673_ (.A(_234_),
    .B(_215_),
    .CIN(_269_),
    .COUT(_270_),
    .SUM(_271_));
 sky130_fd_sc_hd__fa_1 _674_ (.A(_251_),
    .B(_272_),
    .CIN(_273_),
    .COUT(_274_),
    .SUM(_275_));
 sky130_fd_sc_hd__fa_1 _675_ (.A(_271_),
    .B(_254_),
    .CIN(_276_),
    .COUT(_277_),
    .SUM(_278_));
 sky130_fd_sc_hd__fa_1 _676_ (.A(_278_),
    .B(_261_),
    .CIN(_279_),
    .COUT(_280_),
    .SUM(_281_));
 sky130_fd_sc_hd__fa_1 _677_ (.A(_267_),
    .B(_282_),
    .CIN(_283_),
    .COUT(_284_),
    .SUM(_285_));
 sky130_fd_sc_hd__fa_1 _678_ (.A(_271_),
    .B(_270_),
    .CIN(_286_),
    .COUT(_287_),
    .SUM(_288_));
 sky130_fd_sc_hd__fa_1 _679_ (.A(_288_),
    .B(_277_),
    .CIN(_289_),
    .COUT(_290_),
    .SUM(_291_));
 sky130_fd_sc_hd__fa_1 _680_ (.A(_267_),
    .B(_292_),
    .CIN(_293_),
    .COUT(_294_),
    .SUM(_295_));
 sky130_fd_sc_hd__fa_1 _681_ (.A(_271_),
    .B(_270_),
    .CIN(_296_),
    .COUT(_297_),
    .SUM(_298_));
 sky130_fd_sc_hd__fa_1 _682_ (.A(_287_),
    .B(_299_),
    .CIN(_298_),
    .COUT(_300_),
    .SUM(_301_));
 sky130_fd_sc_hd__ha_1 _683_ (.A(_302_),
    .B(start_r),
    .COUT(_303_),
    .SUM(_304_));
 sky130_fd_sc_hd__ha_1 _684_ (.A(net16),
    .B(_305_),
    .COUT(_306_),
    .SUM(_307_));
 sky130_fd_sc_hd__ha_1 _685_ (.A(_308_),
    .B(_309_),
    .COUT(_310_),
    .SUM(_311_));
 sky130_fd_sc_hd__ha_1 _686_ (.A(_310_),
    .B(_312_),
    .COUT(_313_),
    .SUM(_314_));
 sky130_fd_sc_hd__ha_1 _687_ (.A(_313_),
    .B(_315_),
    .COUT(_316_),
    .SUM(_317_));
 sky130_fd_sc_hd__ha_1 _688_ (.A(_318_),
    .B(_319_),
    .COUT(_320_),
    .SUM(_321_));
 sky130_fd_sc_hd__ha_1 _689_ (.A(_322_),
    .B(_323_),
    .COUT(_324_),
    .SUM(_325_));
 sky130_fd_sc_hd__ha_1 _690_ (.A(_316_),
    .B(_325_),
    .COUT(_326_),
    .SUM(_327_));
 sky130_fd_sc_hd__ha_1 _691_ (.A(_328_),
    .B(_329_),
    .COUT(_190_),
    .SUM(_151_));
 sky130_fd_sc_hd__ha_1 _692_ (.A(_330_),
    .B(_331_),
    .COUT(_332_),
    .SUM(_333_));
 sky130_fd_sc_hd__ha_1 _693_ (.A(_334_),
    .B(_333_),
    .COUT(_335_),
    .SUM(_336_));
 sky130_fd_sc_hd__ha_1 _694_ (.A(_324_),
    .B(_337_),
    .COUT(_334_),
    .SUM(_338_));
 sky130_fd_sc_hd__ha_1 _695_ (.A(_135_),
    .B(_182_),
    .COUT(_207_),
    .SUM(_340_));
 sky130_fd_sc_hd__ha_1 _696_ (.A(_341_),
    .B(_332_),
    .COUT(_342_),
    .SUM(_343_));
 sky130_fd_sc_hd__ha_1 _697_ (.A(_344_),
    .B(_345_),
    .COUT(_346_),
    .SUM(_347_));
 sky130_fd_sc_hd__ha_1 _698_ (.A(_348_),
    .B(_349_),
    .COUT(_220_),
    .SUM(_350_));
 sky130_fd_sc_hd__ha_1 _699_ (.A(_351_),
    .B(_209_),
    .COUT(_352_),
    .SUM(_353_));
 sky130_fd_sc_hd__ha_1 _700_ (.A(_354_),
    .B(_345_),
    .COUT(_355_),
    .SUM(_356_));
 sky130_fd_sc_hd__ha_1 _701_ (.A(_357_),
    .B(_358_),
    .COUT(_239_),
    .SUM(_221_));
 sky130_fd_sc_hd__ha_1 _702_ (.A(_208_),
    .B(_359_),
    .COUT(_360_),
    .SUM(_361_));
 sky130_fd_sc_hd__ha_1 _703_ (.A(_362_),
    .B(_363_),
    .COUT(_256_),
    .SUM(_238_));
 sky130_fd_sc_hd__ha_2 _704_ (.A(_364_),
    .B(_365_),
    .COUT(_366_),
    .SUM(_367_));
 sky130_fd_sc_hd__ha_1 _705_ (.A(_368_),
    .B(_369_),
    .COUT(_273_),
    .SUM(_257_));
 sky130_fd_sc_hd__ha_1 _706_ (.A(_370_),
    .B(_371_),
    .COUT(_372_),
    .SUM(_373_));
 sky130_fd_sc_hd__ha_1 _707_ (.A(_375_),
    .B(_376_),
    .COUT(_282_),
    .SUM(_272_));
 sky130_fd_sc_hd__ha_1 _708_ (.A(_377_),
    .B(_378_),
    .COUT(_379_),
    .SUM(_380_));
 sky130_fd_sc_hd__ha_1 _709_ (.A(_374_),
    .B(_381_),
    .COUT(_382_),
    .SUM(_383_));
 sky130_fd_sc_hd__ha_1 _710_ (.A(_384_),
    .B(_385_),
    .COUT(_293_),
    .SUM(_283_));
 sky130_fd_sc_hd__ha_1 _711_ (.A(_386_),
    .B(_387_),
    .COUT(_388_),
    .SUM(_389_));
 sky130_fd_sc_hd__ha_1 _712_ (.A(_384_),
    .B(_390_),
    .COUT(_391_),
    .SUM(_292_));
 sky130_fd_sc_hd__ha_1 _713_ (.A(_267_),
    .B(_292_),
    .COUT(_392_),
    .SUM(_393_));
 sky130_fd_sc_hd__ha_1 _714_ (.A(_394_),
    .B(_395_),
    .COUT(_396_),
    .SUM(_397_));
 sky130_fd_sc_hd__ha_1 _715_ (.A(_326_),
    .B(_338_),
    .COUT(_339_),
    .SUM(_398_));
 sky130_fd_sc_hd__dfrtp_1 \done$_DFFE_PP0P_  (.D(_001_),
    .Q(net17),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[0]$_DFFE_PP0P_  (.D(_002_),
    .Q(net18),
    .RESET_B(_000_),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[10]$_DFFE_PP0P_  (.D(_003_),
    .Q(net19),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[11]$_DFFE_PP0P_  (.D(_004_),
    .Q(net20),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[12]$_DFFE_PP0P_  (.D(_005_),
    .Q(net21),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[13]$_DFFE_PP0P_  (.D(_006_),
    .Q(net22),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[14]$_DFFE_PP0P_  (.D(_007_),
    .Q(net23),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[15]$_DFFE_PP0P_  (.D(_008_),
    .Q(net24),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[1]$_DFFE_PP0P_  (.D(_009_),
    .Q(net25),
    .RESET_B(_000_),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[2]$_DFFE_PP0P_  (.D(_010_),
    .Q(net26),
    .RESET_B(_000_),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[3]$_DFFE_PP0P_  (.D(_011_),
    .Q(net27),
    .RESET_B(_000_),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[4]$_DFFE_PP0P_  (.D(_012_),
    .Q(net28),
    .RESET_B(_000_),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[5]$_DFFE_PP0P_  (.D(_013_),
    .Q(net29),
    .RESET_B(_000_),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[6]$_DFFE_PP0P_  (.D(_014_),
    .Q(net30),
    .RESET_B(_000_),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[7]$_DFFE_PP0P_  (.D(_015_),
    .Q(net31),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[8]$_DFFE_PP0P_  (.D(_016_),
    .Q(net32),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[9]$_DFFE_PP0P_  (.D(_017_),
    .Q(net33),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \start_r$_DFF_PP0_  (.D(net16),
    .Q(start_r),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state$_DFF_PP0_  (.D(_399_),
    .Q(state),
    .RESET_B(_000_),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_69 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(multiplicand[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(multiplicand[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(multiplicand[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(multiplicand[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(multiplicand[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(multiplicand[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(multiplicand[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(multiplier[0]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(multiplier[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input10 (.A(multiplier[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(multiplier[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(multiplier[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(multiplier[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(multiplier[7]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(net34),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(start),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(done));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(product[0]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(product[10]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(product[11]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(product[12]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(product[13]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(product[14]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(product[15]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(product[1]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(product[2]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(product[3]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(product[4]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(product[5]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .X(product[6]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .X(product[7]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net32),
    .X(product[8]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .X(product[9]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(rst),
    .X(net34));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_159 ();
endmodule
